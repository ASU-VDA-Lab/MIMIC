module fake_jpeg_13418_n_612 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_612);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_612;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_5),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_66),
.B(n_70),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_19),
.B(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_16),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

INVx2_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_32),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_103),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_101),
.Y(n_173)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_32),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_36),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_114),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_36),
.B(n_1),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

BUFx4f_ASAP7_75t_SL g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_34),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_55),
.A2(n_15),
.B1(n_14),
.B2(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_57),
.B1(n_44),
.B2(n_26),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_27),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_130),
.B(n_155),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_27),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_159),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_49),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_164),
.B(n_167),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_92),
.B(n_49),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_168),
.B(n_201),
.Y(n_226)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx11_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_69),
.A2(n_60),
.B1(n_45),
.B2(n_54),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_171),
.A2(n_102),
.B1(n_105),
.B2(n_91),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_112),
.B(n_44),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_176),
.B(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_62),
.B(n_23),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_193),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_186),
.B1(n_207),
.B2(n_53),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_57),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_89),
.A2(n_26),
.B1(n_23),
.B2(n_59),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_33),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_187),
.B(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_81),
.B(n_33),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_122),
.Y(n_198)
);

INVx5_ASAP7_75t_SL g269 ( 
.A(n_198),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_75),
.Y(n_199)
);

INVx2_ASAP7_75t_R g200 ( 
.A(n_123),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_100),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_72),
.B(n_45),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_71),
.A2(n_45),
.B1(n_35),
.B2(n_59),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_72),
.B(n_29),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_208),
.B(n_121),
.Y(n_243)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_61),
.Y(n_209)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_214),
.B(n_224),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_216),
.Y(n_309)
);

CKINVDCx11_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_217),
.B(n_243),
.Y(n_331)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

BUFx2_ASAP7_75t_SL g321 ( 
.A(n_218),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_219),
.B(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_221),
.A2(n_50),
.B1(n_41),
.B2(n_188),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_158),
.Y(n_224)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_227),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_261),
.Y(n_288)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_229),
.Y(n_343)
);

CKINVDCx9p33_ASAP7_75t_R g230 ( 
.A(n_142),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_230),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_234),
.A2(n_255),
.B1(n_262),
.B2(n_275),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_45),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_235),
.B(n_236),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_121),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_131),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_129),
.Y(n_239)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_239),
.Y(n_342)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_242),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_171),
.A2(n_78),
.B1(n_97),
.B2(n_111),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_244),
.A2(n_252),
.B1(n_286),
.B2(n_230),
.Y(n_326)
);

CKINVDCx9p33_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_246),
.Y(n_293)
);

CKINVDCx12_ASAP7_75t_R g247 ( 
.A(n_142),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_248),
.B(n_182),
.Y(n_311)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_136),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_249),
.Y(n_299)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_138),
.A2(n_96),
.B1(n_107),
.B2(n_99),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_141),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_253),
.Y(n_308)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_175),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_254),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_177),
.A2(n_80),
.B1(n_67),
.B2(n_63),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_165),
.B(n_128),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_260),
.C(n_187),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_160),
.Y(n_259)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_165),
.B(n_200),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_138),
.B(n_31),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_203),
.A2(n_192),
.B1(n_148),
.B2(n_207),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_146),
.B(n_149),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_266),
.Y(n_289)
);

CKINVDCx12_ASAP7_75t_R g265 ( 
.A(n_169),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_265),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_149),
.B(n_31),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_146),
.B(n_29),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_37),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_194),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_208),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_148),
.A2(n_126),
.B1(n_37),
.B2(n_39),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_135),
.Y(n_276)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_157),
.B(n_21),
.Y(n_277)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_160),
.Y(n_278)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_145),
.Y(n_279)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_147),
.Y(n_280)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_172),
.Y(n_281)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_202),
.A2(n_21),
.B1(n_53),
.B2(n_52),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_301)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_172),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_284),
.B(n_285),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_157),
.B(n_52),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_134),
.A2(n_64),
.B1(n_50),
.B2(n_42),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_151),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_294),
.B(n_215),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_153),
.B1(n_205),
.B2(n_184),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_298),
.A2(n_310),
.B1(n_326),
.B2(n_330),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_303),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_245),
.A2(n_163),
.B1(n_134),
.B2(n_152),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_304),
.A2(n_307),
.B1(n_316),
.B2(n_320),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_143),
.B1(n_140),
.B2(n_188),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_311),
.B(n_273),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_262),
.A2(n_143),
.B1(n_140),
.B2(n_152),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_244),
.A2(n_154),
.B1(n_206),
.B2(n_161),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_234),
.A2(n_137),
.B1(n_166),
.B2(n_162),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_260),
.B(n_185),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_286),
.A2(n_159),
.B1(n_156),
.B2(n_133),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_258),
.A2(n_173),
.B1(n_159),
.B2(n_191),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_269),
.B1(n_282),
.B2(n_229),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_255),
.A2(n_145),
.B(n_191),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_337),
.A2(n_275),
.B(n_257),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_260),
.B(n_15),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_257),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_287),
.B(n_258),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_344),
.B(n_346),
.Y(n_394)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_237),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_326),
.A2(n_254),
.B1(n_238),
.B2(n_223),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_347),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_220),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_348),
.B(n_350),
.Y(n_404)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_289),
.B(n_240),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_269),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_355),
.A2(n_344),
.B(n_359),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_356),
.A2(n_382),
.B1(n_305),
.B2(n_299),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_226),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_357),
.B(n_358),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_313),
.B(n_222),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_360),
.B(n_363),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_274),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_361),
.B(n_384),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_362),
.A2(n_370),
.B(n_377),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_233),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_292),
.B(n_263),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_364),
.B(n_368),
.Y(n_419)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_371),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_331),
.B(n_10),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_340),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_324),
.A2(n_242),
.B1(n_250),
.B2(n_279),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_295),
.Y(n_371)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_324),
.A2(n_256),
.B1(n_253),
.B2(n_227),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_380),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_296),
.B(n_232),
.Y(n_380)
);

INVx13_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_381),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_336),
.A2(n_225),
.B1(n_284),
.B2(n_251),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_294),
.B(n_278),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_387),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_301),
.B(n_281),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_302),
.A2(n_256),
.B1(n_253),
.B2(n_218),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_308),
.B(n_299),
.Y(n_422)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_343),
.Y(n_424)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

OAI32xp33_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_301),
.A3(n_317),
.B1(n_328),
.B2(n_304),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_390),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_389),
.B(n_354),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_351),
.A2(n_317),
.B1(n_337),
.B2(n_301),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_393),
.A2(n_407),
.B(n_372),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_372),
.A2(n_311),
.B(n_308),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_355),
.B(n_300),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_418),
.C(n_349),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_351),
.A2(n_317),
.B1(n_302),
.B2(n_314),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_416),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_353),
.A2(n_323),
.B1(n_338),
.B2(n_325),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_413),
.A2(n_414),
.B1(n_376),
.B2(n_378),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_353),
.A2(n_323),
.B1(n_318),
.B2(n_335),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_375),
.A2(n_334),
.B1(n_216),
.B2(n_259),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_335),
.C(n_315),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

AOI32xp33_ASAP7_75t_L g423 ( 
.A1(n_359),
.A2(n_232),
.A3(n_321),
.B1(n_319),
.B2(n_329),
.Y(n_423)
);

A2O1A1O1Ixp25_ASAP7_75t_L g440 ( 
.A1(n_423),
.A2(n_356),
.B(n_373),
.C(n_381),
.D(n_362),
.Y(n_440)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_424),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_425),
.B(n_427),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_426),
.A2(n_440),
.B(n_442),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_421),
.A2(n_375),
.B1(n_361),
.B2(n_372),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_428),
.A2(n_410),
.B1(n_391),
.B2(n_402),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_397),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_452),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_368),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_433),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_404),
.B(n_350),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_L g460 ( 
.A1(n_434),
.A2(n_435),
.B(n_450),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_421),
.B(n_369),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_358),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_449),
.C(n_455),
.Y(n_483)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_438),
.A2(n_456),
.B1(n_416),
.B2(n_408),
.Y(n_465)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_399),
.Y(n_439)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_393),
.A2(n_367),
.B(n_371),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_392),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_446),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_411),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_345),
.Y(n_445)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_415),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_386),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_448),
.B(n_408),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_374),
.C(n_352),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_390),
.A2(n_382),
.B1(n_387),
.B2(n_365),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_412),
.A2(n_293),
.B(n_327),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_378),
.Y(n_458)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_448),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_461),
.B(n_467),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_449),
.C(n_455),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_458),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_395),
.B1(n_413),
.B2(n_412),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_468),
.A2(n_479),
.B1(n_428),
.B2(n_451),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_422),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_469),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_406),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_470),
.B(n_473),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_427),
.B(n_419),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_486),
.Y(n_498)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_432),
.A2(n_414),
.B1(n_391),
.B2(n_401),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_443),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_480),
.B(n_485),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_436),
.B(n_343),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_484),
.B(n_435),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_445),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_429),
.A2(n_398),
.B1(n_405),
.B2(n_402),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_425),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_420),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_442),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_490),
.A2(n_500),
.B1(n_508),
.B2(n_509),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_513),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_495),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_426),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_506),
.Y(n_519)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_499),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_432),
.B1(n_441),
.B2(n_431),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_501),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_SL g502 ( 
.A(n_487),
.B(n_430),
.C(n_431),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_510),
.B(n_511),
.Y(n_538)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_487),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_514),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_444),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_452),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_507),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_468),
.A2(n_441),
.B1(n_456),
.B2(n_437),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_466),
.A2(n_450),
.B1(n_454),
.B2(n_453),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_462),
.B(n_439),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_463),
.B(n_489),
.C(n_478),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_464),
.C(n_469),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_457),
.B(n_405),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_459),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_466),
.A2(n_438),
.B1(n_398),
.B2(n_403),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_475),
.B1(n_461),
.B2(n_481),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_517),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_516),
.Y(n_545)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_496),
.A2(n_469),
.B(n_488),
.Y(n_525)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_529),
.C(n_539),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_498),
.A2(n_460),
.B1(n_482),
.B2(n_485),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_528),
.Y(n_544)
);

INVxp33_ASAP7_75t_SL g528 ( 
.A(n_503),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_482),
.C(n_462),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_480),
.Y(n_531)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_531),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_498),
.A2(n_493),
.B1(n_494),
.B2(n_496),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_536),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_507),
.A2(n_459),
.B1(n_481),
.B2(n_476),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_510),
.B(n_502),
.Y(n_537)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_537),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_497),
.C(n_513),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_507),
.A2(n_476),
.B1(n_472),
.B2(n_471),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_540),
.B(n_509),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_539),
.B(n_491),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_551),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_545),
.B(n_525),
.C(n_518),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_531),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_552),
.Y(n_566)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_549),
.Y(n_565)
);

BUFx12f_ASAP7_75t_SL g550 ( 
.A(n_538),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_550),
.A2(n_522),
.B(n_537),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_535),
.A2(n_490),
.B1(n_508),
.B2(n_500),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_505),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_486),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_554),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_526),
.B(n_472),
.C(n_420),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_519),
.B(n_327),
.C(n_319),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_555),
.B(n_519),
.C(n_536),
.Y(n_560)
);

INVx13_ASAP7_75t_L g556 ( 
.A(n_540),
.Y(n_556)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_556),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_559),
.B(n_560),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_561),
.B(n_564),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_557),
.A2(n_521),
.B1(n_534),
.B2(n_532),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_562),
.A2(n_570),
.B1(n_571),
.B2(n_558),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_533),
.C(n_518),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_535),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_567),
.B(n_572),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_550),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_541),
.A2(n_530),
.B1(n_523),
.B2(n_527),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_542),
.A2(n_379),
.B1(n_366),
.B2(n_334),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_546),
.B(n_366),
.C(n_312),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_312),
.C(n_173),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_574),
.B(n_555),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_576),
.A2(n_574),
.B1(n_549),
.B2(n_556),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_573),
.B(n_542),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_579),
.B(n_580),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_564),
.C(n_560),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_585),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_551),
.C(n_547),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_583),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_563),
.B(n_547),
.C(n_558),
.Y(n_583)
);

INVx11_ASAP7_75t_L g584 ( 
.A(n_569),
.Y(n_584)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_584),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_L g586 ( 
.A(n_572),
.B(n_544),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_586),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_580),
.B(n_566),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_587),
.B(n_589),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_568),
.C(n_565),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_591),
.B(n_593),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_1),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_595),
.B(n_577),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_599),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_575),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_588),
.B(n_584),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_601),
.C(n_577),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_589),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_603),
.B(n_3),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_596),
.A2(n_594),
.B(n_582),
.Y(n_604)
);

AOI322xp5_ASAP7_75t_L g606 ( 
.A1(n_604),
.A2(n_605),
.A3(n_602),
.B1(n_598),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_597),
.A2(n_594),
.B(n_249),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_607),
.C(n_6),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_6),
.C(n_7),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_609),
.B(n_6),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_7),
.B(n_8),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_611),
.A2(n_7),
.B(n_9),
.Y(n_612)
);


endmodule