module fake_jpeg_10158_n_173 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_21),
.Y(n_42)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_50),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_28),
.C(n_16),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_28),
.C(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_52),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_14),
.B1(n_18),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_14),
.B1(n_24),
.B2(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_18),
.C(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_17),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_49),
.B1(n_23),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_14),
.B1(n_37),
.B2(n_36),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_70),
.B1(n_51),
.B2(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_58),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_69),
.CON(n_76),
.SN(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_54),
.B1(n_43),
.B2(n_32),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_15),
.B(n_27),
.C(n_25),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_27),
.B(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_85),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_78),
.B1(n_91),
.B2(n_59),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_52),
.B1(n_40),
.B2(n_41),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_43),
.B(n_27),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_88),
.C(n_90),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_70),
.B(n_60),
.C(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_71),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_70),
.C(n_72),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_43),
.B(n_54),
.C(n_23),
.Y(n_86)
);

OAI31xp33_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_70),
.A3(n_65),
.B(n_61),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_54),
.C(n_20),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_92),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_1),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_12),
.B1(n_10),
.B2(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_1),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_97),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_96),
.B1(n_104),
.B2(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_12),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_2),
.C(n_3),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_90),
.C(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_76),
.B(n_84),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_115),
.B(n_98),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_88),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_124),
.C(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_120),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_75),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_82),
.C(n_5),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_126),
.C(n_128),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_109),
.C(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_132),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_104),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

OA21x2_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_99),
.B(n_94),
.Y(n_135)
);

AOI321xp33_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_113),
.A3(n_117),
.B1(n_119),
.B2(n_124),
.C(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_143),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_131),
.B(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_4),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_104),
.B1(n_118),
.B2(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_146),
.C(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.C(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_129),
.C(n_125),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_138),
.C(n_141),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_134),
.B(n_127),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_139),
.B(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_143),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_161),
.Y(n_165)
);

OAI21x1_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_160),
.B(n_150),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_9),
.C(n_7),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_8),
.B(n_9),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_7),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_162),
.C(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);


endmodule