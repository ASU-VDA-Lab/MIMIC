module fake_jpeg_4644_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_16),
.Y(n_21)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_28),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_10),
.B1(n_11),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_21),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_11),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_27),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_44),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_28),
.B1(n_19),
.B2(n_26),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_24),
.C(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_35),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_11),
.B(n_27),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_35),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_28),
.B1(n_11),
.B2(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_56),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_25),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_34),
.A3(n_29),
.B1(n_35),
.B2(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_37),
.B1(n_33),
.B2(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_68),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_44),
.B1(n_40),
.B2(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_40),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_52),
.B1(n_68),
.B2(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_31),
.C(n_25),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_60),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_52),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_77),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_37),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_62),
.C(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_62),
.B1(n_53),
.B2(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_70),
.B1(n_74),
.B2(n_25),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_24),
.B1(n_27),
.B2(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_91),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_83),
.C(n_86),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_24),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_8),
.B1(n_9),
.B2(n_2),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_92),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.C(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_95),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_96),
.B(n_97),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_9),
.B(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_5),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);


endmodule