module fake_jpeg_2968_n_259 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_69),
.Y(n_82)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_1),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_68),
.B(n_39),
.C(n_27),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_64),
.Y(n_112)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_2),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_13),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_73),
.Y(n_104)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_3),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_35),
.B1(n_17),
.B2(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_76),
.A2(n_96),
.B1(n_111),
.B2(n_12),
.Y(n_136)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_6),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_102),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_34),
.B1(n_31),
.B2(n_17),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_90),
.B1(n_12),
.B2(n_107),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_33),
.B1(n_38),
.B2(n_30),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_38),
.B1(n_30),
.B2(n_33),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_13),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_99),
.C(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_39),
.B1(n_27),
.B2(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_4),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_24),
.B1(n_22),
.B2(n_8),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_72),
.B1(n_74),
.B2(n_50),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_51),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_44),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_56),
.B(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_47),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_119),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2x1_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_74),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_63),
.B1(n_65),
.B2(n_54),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_136),
.B1(n_142),
.B2(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_126),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_9),
.C(n_10),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_113),
.C(n_117),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_10),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_12),
.Y(n_138)
);

BUFx2_ASAP7_75t_SL g139 ( 
.A(n_109),
.Y(n_139)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_108),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_87),
.B1(n_110),
.B2(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_91),
.A2(n_103),
.B1(n_86),
.B2(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_76),
.A2(n_103),
.B1(n_78),
.B2(n_86),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_91),
.B1(n_101),
.B2(n_77),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_108),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_101),
.B(n_97),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_133),
.B(n_130),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_122),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_162),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_169),
.B1(n_142),
.B2(n_137),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_146),
.B1(n_123),
.B2(n_130),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_114),
.B1(n_97),
.B2(n_106),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_147),
.B1(n_137),
.B2(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_106),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_114),
.B1(n_117),
.B2(n_77),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_133),
.C(n_120),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_189),
.B1(n_194),
.B2(n_162),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_127),
.B(n_129),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_166),
.B(n_129),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_180),
.B(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_138),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_124),
.B(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_190),
.B(n_192),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_131),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_173),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_134),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_156),
.B(n_163),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_184),
.B(n_185),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_157),
.B1(n_160),
.B2(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_206),
.B1(n_210),
.B2(n_179),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_169),
.B1(n_154),
.B2(n_160),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_158),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_159),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_180),
.CI(n_183),
.CON(n_211),
.SN(n_211)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_200),
.C(n_203),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_176),
.B1(n_188),
.B2(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_215),
.B1(n_221),
.B2(n_222),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_213),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_223),
.B(n_197),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_186),
.B1(n_193),
.B2(n_194),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_202),
.B(n_197),
.C(n_198),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_209),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_205),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_227),
.C(n_221),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_191),
.C(n_159),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_229),
.B(n_231),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_200),
.C(n_196),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_211),
.B(n_204),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_235),
.B(n_239),
.Y(n_240)
);

OAI322xp33_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_216),
.A3(n_204),
.B1(n_211),
.B2(n_217),
.C1(n_222),
.C2(n_223),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_213),
.B1(n_210),
.B2(n_192),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_225),
.B1(n_232),
.B2(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_228),
.B(n_196),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_172),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_164),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_227),
.C(n_224),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_245),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_244),
.B1(n_236),
.B2(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_172),
.C(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_233),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_248),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_164),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_168),
.B1(n_174),
.B2(n_256),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_174),
.Y(n_259)
);


endmodule