module fake_netlist_5_702_n_137 (n_16, n_0, n_12, n_9, n_25, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_137);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_137;

wire n_91;
wire n_82;
wire n_122;
wire n_124;
wire n_86;
wire n_136;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_123;
wire n_38;
wire n_113;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_120;
wire n_135;
wire n_30;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_29;
wire n_79;
wire n_131;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_26;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_4),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_33),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_10),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_43),
.Y(n_55)
);

AND3x2_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_2),
.C(n_3),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_40),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_59),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_58),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_53),
.Y(n_76)
);

OAI21x1_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_62),
.B(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_46),
.B1(n_62),
.B2(n_48),
.Y(n_80)
);

OR2x6_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

OAI21x1_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_46),
.B(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI21x1_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_46),
.B(n_58),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_46),
.B(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_47),
.B1(n_65),
.B2(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_76),
.Y(n_89)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_74),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_84),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_R g96 ( 
.A(n_81),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_R g100 ( 
.A(n_91),
.B(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_88),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_104),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_83),
.B1(n_85),
.B2(n_93),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_99),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_99),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_105),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_117),
.B(n_119),
.Y(n_129)
);

OAI221xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_119),
.B1(n_120),
.B2(n_113),
.C(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_126),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_127),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_122),
.B1(n_118),
.B2(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_133),
.B1(n_125),
.B2(n_106),
.C(n_118),
.Y(n_137)
);


endmodule