module fake_jpeg_29222_n_94 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_1),
.Y(n_53)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_37),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_35),
.B1(n_17),
.B2(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_16),
.B1(n_4),
.B2(n_6),
.Y(n_69)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_39),
.C(n_15),
.Y(n_63)
);

XNOR2x1_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_67),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_68),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_13),
.B1(n_18),
.B2(n_20),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_3),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_7),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_74),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_80),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_8),
.B(n_12),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_84),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_59),
.B1(n_21),
.B2(n_23),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_76),
.B(n_73),
.C(n_77),
.D(n_24),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_R g88 ( 
.A(n_87),
.B(n_84),
.C(n_85),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_73),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_76),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_92),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_86),
.Y(n_94)
);


endmodule