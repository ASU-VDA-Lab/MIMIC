module fake_jpeg_18246_n_280 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_280);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_27),
.B1(n_26),
.B2(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_32),
.B1(n_27),
.B2(n_13),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_22),
.B1(n_13),
.B2(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_22),
.B1(n_15),
.B2(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_13),
.B1(n_22),
.B2(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_67),
.B1(n_39),
.B2(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_64),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_35),
.B1(n_29),
.B2(n_36),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_76),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_42),
.A3(n_41),
.B1(n_46),
.B2(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_16),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_85),
.B1(n_84),
.B2(n_72),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_53),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_39),
.B1(n_48),
.B2(n_49),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_56),
.B1(n_51),
.B2(n_52),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_21),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_48),
.B1(n_49),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_37),
.B1(n_65),
.B2(n_64),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_27),
.B(n_19),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_66),
.B1(n_47),
.B2(n_58),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_92),
.B1(n_105),
.B2(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_36),
.C(n_35),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_103),
.C(n_21),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_21),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_101),
.B1(n_87),
.B2(n_70),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_21),
.C(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_69),
.B(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_80),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_15),
.B1(n_23),
.B2(n_20),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_122),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_74),
.A3(n_83),
.B1(n_81),
.B2(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_83),
.B1(n_81),
.B2(n_74),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_117),
.B(n_121),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_118),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_77),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_17),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_86),
.B(n_80),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_87),
.B1(n_70),
.B2(n_86),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_23),
.B1(n_24),
.B2(n_20),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_92),
.B1(n_98),
.B2(n_96),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_77),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_21),
.C(n_16),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_99),
.C(n_106),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_133),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_16),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_100),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_138),
.B(n_146),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_97),
.B(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_100),
.B1(n_91),
.B2(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_147),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_119),
.C(n_129),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_93),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_54),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_111),
.B1(n_117),
.B2(n_113),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_20),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_138),
.C(n_146),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_18),
.B(n_17),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_168),
.B1(n_169),
.B2(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_117),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_109),
.B1(n_108),
.B2(n_24),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_109),
.B1(n_108),
.B2(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_18),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_130),
.B(n_20),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_6),
.B(n_10),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_178),
.B1(n_133),
.B2(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_186),
.B1(n_6),
.B2(n_10),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_184),
.C(n_166),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_142),
.C(n_151),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_135),
.B1(n_147),
.B2(n_136),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_137),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_139),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_196),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_191),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_18),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_17),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_16),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_5),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_169),
.B1(n_155),
.B2(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_161),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_216),
.Y(n_221)
);

NOR4xp25_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_166),
.C(n_167),
.D(n_177),
.Y(n_211)
);

NOR2x1_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_5),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_162),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_163),
.C(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_190),
.C(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_217),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_180),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_219),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_192),
.C(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_197),
.C(n_1),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_0),
.C(n_1),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_229),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_5),
.B(n_10),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_230),
.B1(n_232),
.B2(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_240),
.B1(n_220),
.B2(n_5),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_206),
.B1(n_205),
.B2(n_201),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_205),
.B1(n_201),
.B2(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_208),
.Y(n_242)
);

HB1xp67_ASAP7_75t_SL g243 ( 
.A(n_218),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_4),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_208),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_4),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_221),
.C(n_224),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_252),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_7),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_4),
.B(n_8),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_0),
.B(n_1),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_3),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_7),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_3),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_249),
.B1(n_254),
.B2(n_247),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_245),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_261),
.B(n_242),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_3),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_269),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_244),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_260),
.B(n_8),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_3),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_9),
.B(n_1),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_267),
.B(n_268),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_9),
.C(n_1),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_277),
.B(n_275),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_278),
.A2(n_0),
.B(n_2),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_2),
.Y(n_280)
);


endmodule