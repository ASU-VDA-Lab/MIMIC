module fake_jpeg_3482_n_231 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_231);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_14),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_12),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_74),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_74),
.B1(n_59),
.B2(n_58),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_56),
.B1(n_67),
.B2(n_79),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_62),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_89),
.B(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_70),
.B1(n_60),
.B2(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_102),
.B1(n_68),
.B2(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_101),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_107),
.B(n_6),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_110),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_55),
.B1(n_81),
.B2(n_76),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_60),
.B1(n_79),
.B2(n_57),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_115),
.B1(n_118),
.B2(n_2),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_102),
.B1(n_75),
.B2(n_72),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_114),
.Y(n_142)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_73),
.B1(n_64),
.B2(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_61),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_78),
.C(n_5),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_5),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_90),
.Y(n_128)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_133),
.B1(n_138),
.B2(n_143),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_66),
.B1(n_71),
.B2(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_1),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_137),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_24),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_25),
.C(n_53),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_151),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_115),
.B1(n_23),
.B2(n_26),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_171),
.B1(n_10),
.B2(n_13),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_22),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_157),
.B(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_54),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_161),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_21),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_6),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_160),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_14),
.B(n_15),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_165),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_176),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_30),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_181),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_186),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_31),
.B(n_50),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_20),
.B(n_38),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_155),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_52),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_15),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_32),
.C(n_44),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_156),
.B1(n_149),
.B2(n_171),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_169),
.B1(n_170),
.B2(n_166),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_200),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_29),
.B(n_40),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_34),
.B(n_37),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_178),
.B1(n_174),
.B2(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_192),
.B(n_183),
.C(n_175),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_176),
.C(n_187),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_216),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_205),
.A2(n_201),
.B(n_194),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_219),
.A2(n_210),
.B1(n_205),
.B2(n_204),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_216),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_48),
.B1(n_17),
.B2(n_18),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_214),
.B(n_17),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.C(n_223),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_222),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_220),
.B(n_16),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_19),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_19),
.Y(n_231)
);


endmodule