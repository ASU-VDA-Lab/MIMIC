module real_jpeg_1431_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_32),
.B1(n_59),
.B2(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_32),
.B1(n_54),
.B2(n_55),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_3),
.B(n_53),
.C(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_3),
.B(n_52),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_3),
.B(n_37),
.C(n_71),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_3),
.B(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_40),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_26),
.C(n_41),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_96),
.Y(n_193)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_5),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_46),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_94)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_122),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_98),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_16),
.B(n_98),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_75),
.C(n_83),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_17),
.A2(n_18),
.B1(n_75),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_49),
.C(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_21),
.A2(n_33),
.B1(n_34),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_21),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_29),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_22),
.A2(n_27),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_28),
.Y(n_30)
);

AO22x1_ASAP7_75t_SL g40 ( 
.A1(n_23),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_26),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_27),
.B(n_78),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_27),
.A2(n_29),
.B(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_31),
.B(n_113),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_33),
.A2(n_34),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_33),
.B(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_33),
.A2(n_34),
.B1(n_106),
.B2(n_108),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_33),
.B(n_106),
.C(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_35),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_35),
.A2(n_39),
.B(n_44),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

AOI22x1_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_37),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_37),
.B(n_186),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_44),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_67),
.B2(n_68),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_49),
.B(n_106),
.C(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_49),
.A2(n_50),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OA21x2_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_58),
.B(n_63),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_53),
.B(n_59),
.C(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_64),
.B1(n_65),
.B2(n_85),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_59),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_55),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_55),
.B(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_81),
.A2(n_82),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_81),
.A2(n_82),
.B1(n_166),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_82),
.B(n_161),
.C(n_166),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_82),
.B(n_91),
.C(n_193),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.C(n_93),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_93),
.B1(n_109),
.B2(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_86),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_90),
.A2(n_91),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_91),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_181),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_144),
.C(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_93),
.A2(n_128),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_96),
.B(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_108),
.B1(n_136),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_120),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

OAI211xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_147),
.B(n_153),
.C(n_154),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_137),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_137),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_132),
.C(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_143),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_143),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_145),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_155),
.C(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_172),
.B(n_209),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_160),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_203),
.B(n_208),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_197),
.B(n_202),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_189),
.B(n_196),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_183),
.B(n_188),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B(n_182),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_195),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_207),
.Y(n_208)
);


endmodule