module real_aes_9006_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g535 ( .A(n_1), .Y(n_535) );
INVx1_ASAP7_75t_L g201 ( .A(n_2), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_3), .A2(n_39), .B1(n_163), .B2(n_477), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g142 ( .A1(n_4), .A2(n_143), .B(n_150), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_5), .B(n_136), .Y(n_526) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_7), .A2(n_242), .B(n_243), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g160 ( .A(n_9), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_10), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_12), .B(n_173), .Y(n_472) );
INVx1_ASAP7_75t_L g248 ( .A(n_13), .Y(n_248) );
INVx1_ASAP7_75t_L g530 ( .A(n_14), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_15), .B(n_137), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_16), .A2(n_746), .B1(n_747), .B2(n_750), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_16), .Y(n_750) );
AO32x2_ASAP7_75t_L g492 ( .A1(n_17), .A2(n_136), .A3(n_170), .B1(n_493), .B2(n_497), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_18), .B(n_163), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_19), .B(n_189), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_20), .B(n_137), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_21), .A2(n_52), .B1(n_163), .B2(n_477), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_22), .B(n_143), .Y(n_213) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_23), .A2(n_78), .B1(n_163), .B2(n_173), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_24), .B(n_163), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_25), .B(n_134), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_26), .A2(n_246), .B(n_247), .C(n_249), .Y(n_245) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_27), .A2(n_76), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_27), .Y(n_749) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_28), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_29), .B(n_166), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_30), .B(n_158), .Y(n_203) );
INVx1_ASAP7_75t_L g179 ( .A(n_31), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_32), .B(n_166), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_33), .B(n_445), .Y(n_450) );
INVx2_ASAP7_75t_L g146 ( .A(n_34), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_35), .B(n_163), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_36), .B(n_166), .Y(n_478) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_37), .A2(n_64), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_37), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_38), .A2(n_148), .B(n_153), .C(n_215), .Y(n_214) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_40), .A2(n_453), .B1(n_744), .B2(n_745), .C1(n_751), .C2(n_755), .Y(n_452) );
INVx1_ASAP7_75t_L g177 ( .A(n_42), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_43), .B(n_158), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_44), .B(n_163), .Y(n_520) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_45), .A2(n_122), .A3(n_445), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_45), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_46), .A2(n_89), .B1(n_220), .B2(n_477), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_47), .B(n_163), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_48), .B(n_163), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_49), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_50), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_51), .B(n_143), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_53), .A2(n_62), .B1(n_163), .B2(n_173), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_54), .A2(n_153), .B1(n_173), .B2(n_175), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_55), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_56), .B(n_163), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_57), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_58), .B(n_163), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_59), .A2(n_157), .B(n_159), .C(n_162), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_60), .Y(n_266) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
INVx1_ASAP7_75t_L g149 ( .A(n_63), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_64), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_65), .B(n_163), .Y(n_536) );
INVx1_ASAP7_75t_L g140 ( .A(n_66), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
AO32x2_ASAP7_75t_L g502 ( .A1(n_68), .A2(n_136), .A3(n_228), .B1(n_497), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g547 ( .A(n_69), .Y(n_547) );
INVx1_ASAP7_75t_L g485 ( .A(n_70), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_SL g188 ( .A1(n_71), .A2(n_162), .B(n_189), .C(n_190), .Y(n_188) );
INVxp67_ASAP7_75t_L g191 ( .A(n_72), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_73), .B(n_173), .Y(n_486) );
INVx1_ASAP7_75t_L g107 ( .A(n_74), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_75), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_76), .Y(n_748) );
INVx1_ASAP7_75t_L g259 ( .A(n_77), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_79), .A2(n_148), .B(n_153), .C(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_80), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_81), .B(n_173), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_82), .B(n_202), .Y(n_216) );
INVx2_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_84), .B(n_189), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_85), .A2(n_104), .B1(n_115), .B2(n_758), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_86), .B(n_173), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_87), .A2(n_148), .B(n_153), .C(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
OR2x2_ASAP7_75t_L g446 ( .A(n_88), .B(n_111), .Y(n_446) );
OR2x2_ASAP7_75t_L g458 ( .A(n_88), .B(n_112), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_90), .A2(n_102), .B1(n_173), .B2(n_174), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_91), .B(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_92), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_93), .A2(n_148), .B(n_153), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_94), .Y(n_238) );
INVx1_ASAP7_75t_L g187 ( .A(n_95), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_96), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_97), .B(n_202), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_98), .B(n_173), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_99), .B(n_136), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_100), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_101), .A2(n_143), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g759 ( .A(n_105), .Y(n_759) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g756 ( .A(n_109), .Y(n_756) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g460 ( .A(n_110), .B(n_112), .Y(n_460) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AO21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_451), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g757 ( .A(n_119), .Y(n_757) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_122), .B(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_127), .B2(n_444), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_127), .A2(n_462), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_L g444 ( .A(n_128), .Y(n_444) );
AND3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_366), .C(n_411), .Y(n_128) );
NOR4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_289), .C(n_330), .D(n_347), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_193), .B(n_209), .C(n_251), .Y(n_130) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_167), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_132), .B(n_194), .Y(n_193) );
NOR4xp25_ASAP7_75t_L g313 ( .A(n_132), .B(n_307), .C(n_314), .D(n_320), .Y(n_313) );
AND2x2_ASAP7_75t_L g386 ( .A(n_132), .B(n_275), .Y(n_386) );
AND2x2_ASAP7_75t_L g405 ( .A(n_132), .B(n_351), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_132), .B(n_400), .Y(n_414) );
AND2x2_ASAP7_75t_L g427 ( .A(n_132), .B(n_208), .Y(n_427) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_SL g272 ( .A(n_133), .Y(n_272) );
AND2x2_ASAP7_75t_L g279 ( .A(n_133), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g329 ( .A(n_133), .B(n_168), .Y(n_329) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_133), .B(n_275), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_133), .B(n_168), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_133), .B(n_278), .Y(n_353) );
BUFx2_ASAP7_75t_L g376 ( .A(n_133), .Y(n_376) );
AND2x2_ASAP7_75t_L g380 ( .A(n_133), .B(n_184), .Y(n_380) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_142), .B(n_165), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_135), .B(n_223), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_135), .B(n_497), .C(n_513), .Y(n_512) );
AO21x1_ASAP7_75t_L g550 ( .A1(n_135), .A2(n_513), .B(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_136), .A2(n_185), .B(n_192), .Y(n_184) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_136), .A2(n_518), .B(n_526), .Y(n_517) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_138), .B(n_139), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx2_ASAP7_75t_L g242 ( .A(n_143), .Y(n_242) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_144), .B(n_148), .Y(n_181) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g525 ( .A(n_145), .Y(n_525) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx1_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx3_ASAP7_75t_L g161 ( .A(n_147), .Y(n_161) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx1_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
INVx4_ASAP7_75t_SL g164 ( .A(n_148), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_148), .A2(n_470), .B(n_474), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_148), .A2(n_484), .B(n_487), .Y(n_483) );
BUFx3_ASAP7_75t_L g497 ( .A(n_148), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_148), .A2(n_519), .B(n_522), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_148), .A2(n_529), .B(n_533), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_164), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_152), .A2(n_164), .B(n_187), .C(n_188), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_152), .A2(n_164), .B(n_244), .C(n_245), .Y(n_243) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
BUFx3_ASAP7_75t_L g220 ( .A(n_154), .Y(n_220) );
INVx1_ASAP7_75t_L g477 ( .A(n_154), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_157), .A2(n_475), .B(n_476), .Y(n_474) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_157), .A2(n_534), .B(n_547), .C(n_548), .Y(n_546) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g234 ( .A(n_158), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_158), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g503 ( .A1(n_158), .A2(n_161), .B1(n_504), .B2(n_505), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_158), .A2(n_495), .B1(n_514), .B2(n_515), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_161), .B(n_191), .Y(n_190) );
INVx5_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
O2A1O1Ixp5_ASAP7_75t_SL g484 ( .A1(n_162), .A2(n_202), .B(n_485), .C(n_486), .Y(n_484) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_163), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_164), .A2(n_172), .B1(n_180), .B2(n_181), .Y(n_171) );
INVx1_ASAP7_75t_L g207 ( .A(n_166), .Y(n_207) );
INVx2_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_166), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_166), .A2(n_469), .B(n_478), .Y(n_468) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_166), .A2(n_483), .B(n_490), .Y(n_482) );
OR2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
AND2x2_ASAP7_75t_L g208 ( .A(n_168), .B(n_184), .Y(n_208) );
BUFx2_ASAP7_75t_L g282 ( .A(n_168), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_168), .A2(n_315), .B1(n_317), .B2(n_318), .Y(n_314) );
OR2x2_ASAP7_75t_L g336 ( .A(n_168), .B(n_196), .Y(n_336) );
AND2x2_ASAP7_75t_L g400 ( .A(n_168), .B(n_278), .Y(n_400) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g268 ( .A(n_169), .B(n_196), .Y(n_268) );
AND2x2_ASAP7_75t_L g275 ( .A(n_169), .B(n_184), .Y(n_275) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_169), .Y(n_317) );
OR2x2_ASAP7_75t_L g352 ( .A(n_169), .B(n_195), .Y(n_352) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_182), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_170), .B(n_183), .Y(n_182) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_170), .A2(n_197), .B(n_205), .Y(n_196) );
INVx2_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
INVx2_ASAP7_75t_L g204 ( .A(n_173), .Y(n_204) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_175) );
INVx2_ASAP7_75t_L g178 ( .A(n_176), .Y(n_178) );
INVx4_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_181), .A2(n_198), .B(n_199), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_181), .A2(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g271 ( .A(n_184), .Y(n_271) );
INVx3_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
BUFx2_ASAP7_75t_L g304 ( .A(n_184), .Y(n_304) );
AND2x2_ASAP7_75t_L g337 ( .A(n_184), .B(n_272), .Y(n_337) );
INVx1_ASAP7_75t_L g473 ( .A(n_189), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_193), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_208), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_195), .B(n_280), .Y(n_284) );
INVx1_ASAP7_75t_L g312 ( .A(n_195), .Y(n_312) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g278 ( .A(n_196), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .C(n_204), .Y(n_200) );
INVx2_ASAP7_75t_L g495 ( .A(n_202), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_202), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_202), .A2(n_544), .B(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_204), .A2(n_530), .B(n_531), .C(n_532), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_207), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_207), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
NAND2x1_ASAP7_75t_SL g209 ( .A(n_210), .B(n_224), .Y(n_209) );
AND2x2_ASAP7_75t_L g288 ( .A(n_210), .B(n_239), .Y(n_288) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_210), .Y(n_362) );
AND2x2_ASAP7_75t_L g389 ( .A(n_210), .B(n_309), .Y(n_389) );
AND2x2_ASAP7_75t_L g397 ( .A(n_210), .B(n_359), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_210), .B(n_254), .Y(n_424) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g255 ( .A(n_211), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g273 ( .A(n_211), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g294 ( .A(n_211), .Y(n_294) );
INVx1_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_211), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g333 ( .A(n_211), .B(n_257), .Y(n_333) );
OR2x2_ASAP7_75t_L g371 ( .A(n_211), .B(n_326), .Y(n_371) );
AOI32xp33_ASAP7_75t_L g383 ( .A1(n_211), .A2(n_384), .A3(n_387), .B1(n_388), .B2(n_389), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_211), .B(n_359), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_211), .B(n_319), .Y(n_434) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AOI21xp5_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_214), .B(n_221), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_218), .A2(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g249 ( .A(n_220), .Y(n_249) );
INVx1_ASAP7_75t_L g264 ( .A(n_221), .Y(n_264) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_221), .A2(n_528), .B(n_537), .Y(n_527) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_221), .A2(n_542), .B(n_549), .Y(n_541) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g345 ( .A(n_225), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
INVx1_ASAP7_75t_L g307 ( .A(n_226), .Y(n_307) );
AND2x2_ASAP7_75t_L g309 ( .A(n_226), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_226), .B(n_256), .Y(n_326) );
AND2x2_ASAP7_75t_L g359 ( .A(n_226), .B(n_335), .Y(n_359) );
AND2x2_ASAP7_75t_L g396 ( .A(n_226), .B(n_257), .Y(n_396) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_227), .B(n_256), .Y(n_286) );
AND2x2_ASAP7_75t_L g293 ( .A(n_227), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g334 ( .A(n_227), .B(n_335), .Y(n_334) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
INVx2_ASAP7_75t_L g310 ( .A(n_239), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_239), .B(n_256), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_239), .B(n_301), .Y(n_382) );
INVx1_ASAP7_75t_L g404 ( .A(n_239), .Y(n_404) );
INVx1_ASAP7_75t_L g421 ( .A(n_239), .Y(n_421) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g274 ( .A(n_240), .B(n_256), .Y(n_274) );
AND2x2_ASAP7_75t_L g296 ( .A(n_240), .B(n_257), .Y(n_296) );
INVx1_ASAP7_75t_L g335 ( .A(n_240), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_246), .B(n_248), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_246), .A2(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g532 ( .A(n_246), .Y(n_532) );
AOI221x1_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_267), .B1(n_273), .B2(n_275), .C(n_276), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_252), .A2(n_340), .B1(n_407), .B2(n_408), .Y(n_406) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g298 ( .A(n_253), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g393 ( .A(n_253), .B(n_273), .Y(n_393) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g349 ( .A(n_254), .B(n_274), .Y(n_349) );
INVx1_ASAP7_75t_L g361 ( .A(n_255), .Y(n_361) );
AND2x2_ASAP7_75t_L g372 ( .A(n_255), .B(n_359), .Y(n_372) );
AND2x2_ASAP7_75t_L g439 ( .A(n_255), .B(n_334), .Y(n_439) );
INVx2_ASAP7_75t_L g301 ( .A(n_256), .Y(n_301) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_264), .B(n_265), .Y(n_257) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_268), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g391 ( .A(n_268), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_269), .B(n_352), .Y(n_355) );
INVx3_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_270), .A2(n_391), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NOR2xp33_ASAP7_75t_SL g413 ( .A(n_273), .B(n_299), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_274), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g365 ( .A(n_274), .B(n_293), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_274), .B(n_300), .Y(n_442) );
AND2x2_ASAP7_75t_L g311 ( .A(n_275), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g378 ( .A(n_275), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B(n_285), .Y(n_276) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_278), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g327 ( .A(n_278), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g339 ( .A(n_278), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_278), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g363 ( .A(n_279), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_279), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_279), .B(n_282), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_282), .A2(n_321), .B(n_351), .C(n_353), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_282), .A2(n_369), .B1(n_372), .B2(n_373), .C(n_377), .Y(n_368) );
AND2x2_ASAP7_75t_L g364 ( .A(n_283), .B(n_317), .Y(n_364) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g324 ( .A(n_288), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g395 ( .A(n_288), .B(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_297), .C(n_322), .Y(n_289) );
NAND3xp33_ASAP7_75t_SL g408 ( .A(n_290), .B(n_409), .C(n_410), .Y(n_408) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
OR2x2_ASAP7_75t_L g381 ( .A(n_292), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_302), .B1(n_305), .B2(n_311), .C(n_313), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_299), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_299), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g321 ( .A(n_304), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_304), .A2(n_361), .B1(n_362), .B2(n_363), .Y(n_360) );
OR2x2_ASAP7_75t_L g441 ( .A(n_304), .B(n_352), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVxp67_ASAP7_75t_L g415 ( .A(n_307), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_309), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_312), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_312), .B(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_312), .B(n_379), .Y(n_418) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g432 ( .A(n_321), .B(n_352), .Y(n_432) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g410 ( .A(n_327), .Y(n_410) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI322xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_336), .A3(n_337), .B1(n_338), .B2(n_341), .C1(n_343), .C2(n_345), .Y(n_330) );
OAI322xp33_ASAP7_75t_L g412 ( .A1(n_331), .A2(n_413), .A3(n_414), .B1(n_415), .B2(n_416), .C1(n_417), .C2(n_419), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx4_ASAP7_75t_L g346 ( .A(n_333), .Y(n_346) );
AND2x2_ASAP7_75t_L g407 ( .A(n_333), .B(n_359), .Y(n_407) );
AND2x2_ASAP7_75t_L g420 ( .A(n_333), .B(n_421), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_336), .Y(n_431) );
INVx1_ASAP7_75t_L g409 ( .A(n_337), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g343 ( .A(n_339), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g426 ( .A(n_339), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_339), .B(n_380), .Y(n_437) );
OR2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_371), .Y(n_370) );
INVxp33_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
OAI221xp5_ASAP7_75t_SL g347 ( .A1(n_346), .A2(n_348), .B1(n_350), .B2(n_354), .C(n_356), .Y(n_347) );
NOR2xp67_ASAP7_75t_L g403 ( .A(n_346), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g430 ( .A(n_346), .Y(n_430) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx3_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AOI322xp5_ASAP7_75t_L g394 ( .A1(n_353), .A2(n_378), .A3(n_395), .B1(n_397), .B2(n_398), .C1(n_401), .C2(n_405), .Y(n_394) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B1(n_364), .B2(n_365), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_390), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_368), .B(n_383), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_371), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NAND2xp33_ASAP7_75t_SL g388 ( .A(n_374), .B(n_385), .Y(n_388) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OAI322xp33_ASAP7_75t_L g428 ( .A1(n_376), .A2(n_429), .A3(n_431), .B1(n_432), .B2(n_433), .C1(n_435), .C2(n_438), .Y(n_428) );
AOI21xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_379), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_386), .B(n_434), .Y(n_443) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .B(n_394), .C(n_406), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR4xp25_ASAP7_75t_L g411 ( .A(n_412), .B(n_422), .C(n_428), .D(n_440), .Y(n_411) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_442), .B(n_443), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_444), .A2(n_455), .B1(n_459), .B2(n_461), .Y(n_454) );
INVx1_ASAP7_75t_L g449 ( .A(n_445), .Y(n_449) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_450), .A2(n_452), .B(n_757), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g753 ( .A(n_458), .Y(n_753) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx6_ASAP7_75t_L g754 ( .A(n_460), .Y(n_754) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_666), .Y(n_462) );
NAND5xp2_ASAP7_75t_L g463 ( .A(n_464), .B(n_585), .C(n_600), .D(n_626), .E(n_648), .Y(n_463) );
NOR2xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_565), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_506), .B1(n_538), .B2(n_554), .C(n_555), .Y(n_465) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_467), .B(n_498), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_467), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g742 ( .A(n_467), .Y(n_742) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_479), .Y(n_467) );
INVx1_ASAP7_75t_L g582 ( .A(n_468), .Y(n_582) );
AND2x2_ASAP7_75t_L g584 ( .A(n_468), .B(n_492), .Y(n_584) );
AND2x2_ASAP7_75t_L g594 ( .A(n_468), .B(n_491), .Y(n_594) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_468), .Y(n_612) );
INVx1_ASAP7_75t_L g622 ( .A(n_468), .Y(n_622) );
OR2x2_ASAP7_75t_L g660 ( .A(n_468), .B(n_559), .Y(n_660) );
INVx2_ASAP7_75t_L g710 ( .A(n_468), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_468), .B(n_558), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_473), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_480), .B(n_491), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_481), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_481), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_SL g642 ( .A(n_481), .B(n_582), .Y(n_642) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_482), .Y(n_500) );
INVx2_ASAP7_75t_L g559 ( .A(n_482), .Y(n_559) );
OR2x2_ASAP7_75t_L g621 ( .A(n_482), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g560 ( .A(n_491), .B(n_502), .Y(n_560) );
AND2x2_ASAP7_75t_L g577 ( .A(n_491), .B(n_557), .Y(n_577) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g501 ( .A(n_492), .B(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g580 ( .A(n_492), .Y(n_580) );
AND2x2_ASAP7_75t_L g709 ( .A(n_492), .B(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_495), .A2(n_523), .B(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_495), .A2(n_534), .B(n_535), .C(n_536), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_497), .A2(n_543), .B(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g554 ( .A(n_498), .Y(n_554) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x2_ASAP7_75t_L g672 ( .A(n_499), .B(n_560), .Y(n_672) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g673 ( .A(n_500), .B(n_584), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_501), .A2(n_641), .B(n_643), .C(n_645), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_501), .B(n_641), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_501), .A2(n_571), .B1(n_714), .B2(n_715), .C(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g557 ( .A(n_502), .Y(n_557) );
INVx1_ASAP7_75t_L g593 ( .A(n_502), .Y(n_593) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_502), .Y(n_602) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
AND2x2_ASAP7_75t_L g619 ( .A(n_508), .B(n_564), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_508), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_509), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g711 ( .A(n_509), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g743 ( .A(n_509), .Y(n_743) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g573 ( .A(n_510), .Y(n_573) );
AND2x2_ASAP7_75t_L g599 ( .A(n_510), .B(n_553), .Y(n_599) );
NOR2x1_ASAP7_75t_L g608 ( .A(n_510), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g615 ( .A(n_510), .B(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g551 ( .A(n_511), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_516), .B(n_655), .Y(n_690) );
INVx1_ASAP7_75t_SL g694 ( .A(n_516), .Y(n_694) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx3_ASAP7_75t_L g553 ( .A(n_517), .Y(n_553) );
AND2x2_ASAP7_75t_L g564 ( .A(n_517), .B(n_541), .Y(n_564) );
AND2x2_ASAP7_75t_L g586 ( .A(n_517), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g631 ( .A(n_517), .B(n_625), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_517), .B(n_563), .Y(n_712) );
INVx2_ASAP7_75t_L g534 ( .A(n_525), .Y(n_534) );
AND2x2_ASAP7_75t_L g552 ( .A(n_527), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_527), .B(n_541), .Y(n_588) );
AND2x2_ASAP7_75t_L g624 ( .A(n_527), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_552), .Y(n_539) );
INVx1_ASAP7_75t_L g604 ( .A(n_540), .Y(n_604) );
AND2x2_ASAP7_75t_L g646 ( .A(n_540), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_540), .B(n_567), .Y(n_652) );
AOI21xp5_ASAP7_75t_SL g726 ( .A1(n_540), .A2(n_558), .B(n_581), .Y(n_726) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_550), .Y(n_540) );
OR2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_550), .Y(n_569) );
AND2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_553), .Y(n_616) );
INVx2_ASAP7_75t_L g625 ( .A(n_541), .Y(n_625) );
INVx1_ASAP7_75t_L g731 ( .A(n_541), .Y(n_731) );
AND2x2_ASAP7_75t_L g655 ( .A(n_550), .B(n_625), .Y(n_655) );
INVx1_ASAP7_75t_L g680 ( .A(n_550), .Y(n_680) );
AND2x2_ASAP7_75t_L g589 ( .A(n_552), .B(n_573), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_552), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g719 ( .A(n_552), .Y(n_719) );
INVx2_ASAP7_75t_L g609 ( .A(n_553), .Y(n_609) );
AND2x2_ASAP7_75t_L g647 ( .A(n_553), .B(n_563), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_553), .B(n_731), .Y(n_730) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B(n_561), .Y(n_555) );
AND2x2_ASAP7_75t_L g662 ( .A(n_556), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g716 ( .A(n_556), .Y(n_716) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g636 ( .A(n_557), .Y(n_636) );
BUFx2_ASAP7_75t_L g735 ( .A(n_557), .Y(n_735) );
BUFx2_ASAP7_75t_L g606 ( .A(n_558), .Y(n_606) );
AND2x2_ASAP7_75t_L g708 ( .A(n_558), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g691 ( .A(n_559), .Y(n_691) );
AND2x4_ASAP7_75t_L g618 ( .A(n_560), .B(n_581), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_560), .B(n_642), .Y(n_654) );
AOI32xp33_ASAP7_75t_L g578 ( .A1(n_561), .A2(n_579), .A3(n_581), .B1(n_583), .B2(n_584), .Y(n_578) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx3_ASAP7_75t_L g567 ( .A(n_562), .Y(n_567) );
OR2x2_ASAP7_75t_L g703 ( .A(n_562), .B(n_659), .Y(n_703) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_563), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g679 ( .A(n_563), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g571 ( .A(n_564), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g583 ( .A(n_564), .B(n_573), .Y(n_583) );
INVx1_ASAP7_75t_L g704 ( .A(n_564), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_564), .B(n_679), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_570), .B(n_574), .C(n_578), .Y(n_565) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_566), .A2(n_611), .A3(n_675), .B1(n_677), .B2(n_681), .C1(n_682), .C2(n_686), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVxp67_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g693 ( .A(n_569), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_569), .B(n_609), .Y(n_740) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g632 ( .A(n_572), .Y(n_632) );
OR2x2_ASAP7_75t_L g718 ( .A(n_573), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_576), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g627 ( .A(n_577), .B(n_606), .Y(n_627) );
AND2x2_ASAP7_75t_L g698 ( .A(n_577), .B(n_611), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_577), .B(n_685), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_579), .A2(n_586), .B1(n_589), .B2(n_590), .C(n_595), .Y(n_585) );
OR2x2_ASAP7_75t_L g596 ( .A(n_579), .B(n_592), .Y(n_596) );
AND2x2_ASAP7_75t_L g684 ( .A(n_579), .B(n_685), .Y(n_684) );
AOI32xp33_ASAP7_75t_L g723 ( .A1(n_579), .A2(n_609), .A3(n_724), .B1(n_725), .B2(n_728), .Y(n_723) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_580), .B(n_616), .C(n_639), .Y(n_657) );
AND2x2_ASAP7_75t_L g683 ( .A(n_580), .B(n_676), .Y(n_683) );
INVxp67_ASAP7_75t_L g663 ( .A(n_581), .Y(n_663) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_584), .B(n_636), .Y(n_692) );
INVx2_ASAP7_75t_L g702 ( .A(n_584), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_584), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g671 ( .A(n_587), .Y(n_671) );
OR2x2_ASAP7_75t_L g597 ( .A(n_588), .B(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_590), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_593), .Y(n_676) );
AND2x2_ASAP7_75t_L g635 ( .A(n_594), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g681 ( .A(n_594), .Y(n_681) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_594), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI21xp33_ASAP7_75t_SL g620 ( .A1(n_596), .A2(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g714 ( .A(n_599), .B(n_624), .Y(n_714) );
AOI211xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B(n_613), .C(n_620), .Y(n_600) );
AND2x2_ASAP7_75t_L g644 ( .A(n_602), .B(n_612), .Y(n_644) );
INVx2_ASAP7_75t_L g659 ( .A(n_602), .Y(n_659) );
OR2x2_ASAP7_75t_L g697 ( .A(n_602), .B(n_660), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_602), .B(n_740), .Y(n_739) );
AOI211xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_607), .C(n_610), .Y(n_603) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_606), .B(n_644), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_607), .A2(n_702), .B(n_726), .C(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_608), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g665 ( .A(n_609), .B(n_655), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_609), .Y(n_670) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_617), .Y(n_613) );
INVxp33_ASAP7_75t_L g721 ( .A(n_615), .Y(n_721) );
AND2x2_ASAP7_75t_L g700 ( .A(n_616), .B(n_679), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_621), .A2(n_683), .B(n_684), .Y(n_682) );
OAI322xp33_ASAP7_75t_L g701 ( .A1(n_623), .A2(n_702), .A3(n_703), .B1(n_704), .B2(n_705), .C1(n_707), .C2(n_711), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_633), .B2(n_637), .C(n_640), .Y(n_626) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g678 ( .A(n_631), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g722 ( .A(n_635), .Y(n_722) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_638), .B(n_658), .Y(n_724) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g687 ( .A(n_647), .B(n_655), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_655), .C(n_656), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_651), .A2(n_668), .B1(n_672), .B2(n_673), .C(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_655), .B(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_661), .B2(n_664), .Y(n_656) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_SL g685 ( .A(n_660), .Y(n_685) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND5xp2_ASAP7_75t_L g666 ( .A(n_667), .B(n_688), .C(n_713), .D(n_723), .E(n_733), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_671), .Y(n_668) );
NOR4xp25_ASAP7_75t_L g741 ( .A(n_670), .B(n_676), .C(n_742), .D(n_743), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_673), .A2(n_734), .B1(n_736), .B2(n_738), .C(n_741), .Y(n_733) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g732 ( .A(n_679), .Y(n_732) );
OAI322xp33_ASAP7_75t_L g689 ( .A1(n_683), .A2(n_690), .A3(n_691), .B1(n_692), .B2(n_693), .C1(n_695), .C2(n_699), .Y(n_689) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_701), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g734 ( .A(n_709), .B(n_735), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule