module fake_jpeg_2167_n_217 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_217);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_98),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_71),
.B1(n_70),
.B2(n_59),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_69),
.B1(n_73),
.B2(n_56),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_75),
.B1(n_70),
.B2(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_86),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_106),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_58),
.B(n_62),
.C(n_74),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_95),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_110),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_66),
.C(n_71),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_66),
.C(n_55),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_76),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_116),
.A2(n_55),
.B1(n_75),
.B2(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_60),
.B1(n_76),
.B2(n_25),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_119),
.A2(n_39),
.B1(n_52),
.B2(n_30),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_128),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_127),
.B1(n_11),
.B2(n_12),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_31),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_76),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_0),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_23),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_6),
.C(n_8),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_2),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_4),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_8),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_144),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_137),
.B(n_111),
.C(n_5),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_19),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_19),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_151),
.B1(n_158),
.B2(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_155),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_13),
.B(n_14),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_17),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_134),
.B(n_32),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_171),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_134),
.C(n_33),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_175),
.C(n_153),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_177),
.C(n_182),
.Y(n_193)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_34),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_35),
.B(n_36),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_163),
.B1(n_146),
.B2(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_181),
.B(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_153),
.B1(n_44),
.B2(n_45),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_40),
.B(n_46),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_183),
.B(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_53),
.B1(n_47),
.B2(n_50),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_191),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_167),
.C(n_169),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_204),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_187),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_183),
.B(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_206),
.A2(n_180),
.B1(n_196),
.B2(n_197),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_203),
.B1(n_195),
.B2(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_210),
.C(n_209),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_197),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_176),
.B(n_179),
.C(n_170),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_214),
.A2(n_176),
.B(n_193),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_189),
.Y(n_217)
);


endmodule