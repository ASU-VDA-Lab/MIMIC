module real_jpeg_29140_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_343, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_343;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_0),
.A2(n_37),
.B1(n_58),
.B2(n_61),
.Y(n_107)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_118),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_2),
.A2(n_58),
.B1(n_61),
.B2(n_118),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_118),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_3),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_123),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_123),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_3),
.A2(n_58),
.B1(n_61),
.B2(n_123),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_5),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_26),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_31),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_5),
.A2(n_31),
.B(n_163),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_121),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_58),
.B(n_62),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_80),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_5),
.A2(n_100),
.B1(n_213),
.B2(n_214),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_7),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_116),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_116),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_58),
.B1(n_61),
.B2(n_116),
.Y(n_205)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_9),
.A2(n_46),
.B1(n_58),
.B2(n_61),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_9),
.A2(n_27),
.B1(n_31),
.B2(n_46),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_10),
.A2(n_25),
.B1(n_58),
.B2(n_61),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_48),
.B1(n_58),
.B2(n_61),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_12),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_292)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_15),
.Y(n_60)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_341),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_85),
.B(n_339),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_20),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_21),
.A2(n_44),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_22),
.A2(n_33),
.B(n_84),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g120 ( 
.A(n_23),
.B(n_121),
.CON(n_120),
.SN(n_120)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_26),
.A2(n_33),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_31),
.B1(n_69),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_27),
.A2(n_34),
.B1(n_120),
.B2(n_135),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_53),
.A3(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_29),
.B(n_31),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_32),
.A2(n_45),
.B(n_49),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_33),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_36),
.B(n_49),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_39),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_77),
.C(n_82),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_40),
.A2(n_41),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_65),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_42),
.A2(n_43),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_44),
.A2(n_49),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_44),
.A2(n_49),
.B1(n_129),
.B2(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_50),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_50),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_50),
.A2(n_65),
.B1(n_307),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_63),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_63),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_51),
.A2(n_57),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_51),
.A2(n_171),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_51),
.A2(n_57),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_51),
.A2(n_57),
.B1(n_170),
.B2(n_189),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_51),
.A2(n_57),
.B1(n_95),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_51),
.A2(n_111),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_70),
.Y(n_67)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_54),
.B(n_76),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_54),
.A2(n_56),
.B(n_121),
.C(n_191),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_57),
.B(n_121),
.Y(n_211)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_61),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_64),
.B(n_112),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_66),
.A2(n_79),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_74),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_67),
.A2(n_74),
.B1(n_115),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_67),
.A2(n_74),
.B1(n_146),
.B2(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_67),
.B(n_73),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_67),
.A2(n_74),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_72),
.A2(n_80),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_79),
.A2(n_81),
.B(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_79),
.A2(n_256),
.B(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_82),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_332),
.B(n_338),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_302),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_343),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_283),
.B(n_301),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_260),
.B(n_282),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_152),
.B(n_237),
.C(n_259),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_138),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_91),
.B(n_138),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_124),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_93),
.B(n_108),
.C(n_124),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_94),
.B(n_99),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_96),
.B(n_181),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B(n_105),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_100),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_100),
.A2(n_205),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_100),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_106),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_101),
.A2(n_102),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_160),
.Y(n_200)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_102),
.Y(n_277)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_103),
.A2(n_137),
.B(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_119),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_121),
.B(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_133),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_126),
.B(n_131),
.C(n_133),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_136),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_139),
.A2(n_140),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_149),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_200),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_236),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_229),
.B(n_235),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_182),
.B(n_228),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_172),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_156),
.B(n_172),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.C(n_168),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_157),
.A2(n_158),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_161),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_160),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_179),
.C(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_222),
.B(n_227),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_201),
.B(n_221),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_199),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_209),
.B(n_220),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_207),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_215),
.B(n_219),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_239),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_257),
.B2(n_258),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_248),
.C(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_251),
.C(n_255),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_262),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_281),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_274),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_269),
.C(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_270),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_276),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_279),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_276),
.A2(n_295),
.B(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_285),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_299),
.B2(n_300),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_294),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_294),
.C(n_300),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_293),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_292),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_304),
.C(n_314),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_304),
.B1(n_305),
.B2(n_329),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_293),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_313),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_322),
.C(n_323),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_315),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_335),
.Y(n_337)
);


endmodule