module fake_jpeg_5506_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_53),
.B1(n_55),
.B2(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_26),
.B1(n_23),
.B2(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_26),
.B1(n_23),
.B2(n_27),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_64),
.B1(n_67),
.B2(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_17),
.B(n_19),
.C(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_22),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_27),
.B1(n_24),
.B2(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_17),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_24),
.B1(n_33),
.B2(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_68),
.B(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_72),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_24),
.A3(n_25),
.B1(n_30),
.B2(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_67),
.B1(n_53),
.B2(n_54),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_0),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_48),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_66),
.C(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_51),
.B1(n_60),
.B2(n_45),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_92),
.B1(n_51),
.B2(n_77),
.Y(n_95)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_93),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_67),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_106),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_109),
.B1(n_113),
.B2(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_78),
.B1(n_83),
.B2(n_81),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_57),
.B1(n_52),
.B2(n_66),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_45),
.B1(n_56),
.B2(n_64),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_114),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_88),
.B1(n_70),
.B2(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_68),
.B(n_79),
.C(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_0),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_63),
.B(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_86),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_42),
.C(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_126),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_130),
.B1(n_142),
.B2(n_93),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_129),
.B(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_20),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_89),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_92),
.B1(n_89),
.B2(n_90),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_139),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_92),
.B1(n_42),
.B2(n_62),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_129),
.B1(n_119),
.B2(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_20),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_98),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_63),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_62),
.B1(n_19),
.B2(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_34),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_2),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_108),
.B1(n_113),
.B2(n_101),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_98),
.B(n_102),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_163),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_137),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_153),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_114),
.B1(n_118),
.B2(n_115),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_117),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_129),
.B(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_165),
.Y(n_174)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_115),
.B(n_100),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_97),
.B(n_1),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_52),
.C(n_100),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_157),
.C(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_100),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_168),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_107),
.B(n_1),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_107),
.B1(n_1),
.B2(n_0),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_2),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_171),
.B1(n_119),
.B2(n_4),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_124),
.B1(n_132),
.B2(n_125),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_183),
.B1(n_167),
.B2(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_148),
.B(n_149),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_176),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_152),
.C(n_150),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_189),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_131),
.B(n_5),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_190),
.B(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_6),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_195),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_170),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_7),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_204),
.C(n_212),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_159),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_178),
.C(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_160),
.B1(n_146),
.B2(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_150),
.B1(n_159),
.B2(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_190),
.B1(n_176),
.B2(n_182),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_172),
.B(n_166),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_209),
.B(n_186),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_163),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_161),
.C(n_145),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_154),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_161),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_185),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_190),
.B(n_194),
.C(n_187),
.D(n_188),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_229),
.B1(n_201),
.B2(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_209),
.B(n_205),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_192),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_231),
.C(n_232),
.Y(n_234)
);

BUFx12_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_171),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_196),
.C(n_12),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_206),
.C(n_216),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_218),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_217),
.B1(n_203),
.B2(n_200),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_244),
.B1(n_196),
.B2(n_231),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_243),
.B(n_233),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_213),
.B(n_196),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_217),
.B1(n_196),
.B2(n_199),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_215),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_259)
);

OA21x2_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_227),
.B(n_232),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_202),
.C(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_207),
.B1(n_208),
.B2(n_230),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_245),
.B(n_238),
.Y(n_258)
);

NOR2x1_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

OAI321xp33_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_244),
.A3(n_239),
.B1(n_237),
.B2(n_242),
.C(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_267),
.B(n_15),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_250),
.C(n_12),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_10),
.C(n_12),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_260),
.C(n_262),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_10),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.C1(n_260),
.C2(n_265),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_15),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_275),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_274),
.Y(n_277)
);


endmodule