module fake_jpeg_8853_n_73 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_55;
wire n_27;
wire n_64;
wire n_47;
wire n_51;
wire n_22;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_24;
wire n_38;
wire n_28;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_25;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;
wire n_70;
wire n_66;

BUFx12_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_46),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_47),
.B1(n_39),
.B2(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_52),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_23),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_43),
.C(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_37),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_34),
.B(n_44),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_65),
.A2(n_32),
.B(n_24),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_33),
.B1(n_25),
.B2(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_42),
.B(n_22),
.Y(n_72)
);

AOI221xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_55),
.B1(n_53),
.B2(n_26),
.C(n_22),
.Y(n_73)
);


endmodule