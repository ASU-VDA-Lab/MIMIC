module fake_jpeg_29321_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_18),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_52),
.B(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_54),
.B(n_55),
.Y(n_146)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_13),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_82),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_57),
.Y(n_115)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx2_ASAP7_75t_SL g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_13),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_99),
.Y(n_148)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_29),
.B(n_12),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_90),
.Y(n_137)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_25),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_95),
.Y(n_142)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_30),
.B(n_12),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_42),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_30),
.B(n_11),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

CKINVDCx6p67_ASAP7_75t_R g101 ( 
.A(n_25),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_101),
.Y(n_165)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_44),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_116),
.B(n_152),
.Y(n_227)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_57),
.A2(n_50),
.B1(n_45),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_149),
.B1(n_45),
.B2(n_96),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_80),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_54),
.A2(n_32),
.B1(n_42),
.B2(n_35),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_94),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_61),
.B(n_32),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_154),
.B(n_22),
.Y(n_198)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_49),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_21),
.Y(n_195)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_61),
.B(n_20),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_62),
.B(n_20),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_62),
.B(n_39),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_68),
.B(n_49),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_68),
.B(n_39),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_101),
.C(n_65),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_167),
.B(n_112),
.C(n_156),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_74),
.B1(n_64),
.B2(n_73),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_168),
.A2(n_170),
.B1(n_197),
.B2(n_112),
.Y(n_235)
);

INVx6_ASAP7_75t_SL g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_169),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_115),
.A2(n_97),
.B1(n_70),
.B2(n_102),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_171),
.A2(n_194),
.B1(n_200),
.B2(n_212),
.Y(n_237)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_175),
.B(n_205),
.Y(n_230)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_179),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_181),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_182),
.Y(n_275)
);

OR2x2_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_27),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_184),
.Y(n_274)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_104),
.A2(n_22),
.B1(n_37),
.B2(n_47),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_191),
.B(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_115),
.A2(n_37),
.B(n_47),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_214),
.B(n_195),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_113),
.A2(n_93),
.B1(n_84),
.B2(n_79),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_210),
.Y(n_234)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_66),
.B1(n_78),
.B2(n_76),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_206),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_123),
.A2(n_45),
.B1(n_83),
.B2(n_35),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_113),
.B(n_11),
.Y(n_205)
);

CKINVDCx12_ASAP7_75t_R g206 ( 
.A(n_122),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_208),
.Y(n_262)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

OR2x2_ASAP7_75t_SL g210 ( 
.A(n_157),
.B(n_35),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_143),
.A2(n_45),
.B1(n_83),
.B2(n_27),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_213),
.B(n_215),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_165),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_216),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_217),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_142),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_218),
.B(n_220),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_114),
.A2(n_11),
.B(n_1),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_219),
.A2(n_2),
.B(n_4),
.Y(n_261)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_143),
.A2(n_75),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_133),
.B1(n_145),
.B2(n_124),
.Y(n_252)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_114),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_118),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_140),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_232),
.B(n_187),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_233),
.A2(n_188),
.B(n_217),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_235),
.A2(n_38),
.B1(n_21),
.B2(n_23),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_138),
.B1(n_156),
.B2(n_153),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_239),
.A2(n_248),
.B1(n_268),
.B2(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_153),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_243),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_140),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_197),
.A2(n_126),
.B1(n_138),
.B2(n_139),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_128),
.B1(n_139),
.B2(n_126),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_252),
.B1(n_263),
.B2(n_271),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_173),
.B(n_145),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_256),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_122),
.B(n_107),
.C(n_159),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_253),
.B(n_259),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_180),
.B(n_0),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_122),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_261),
.B(n_5),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_223),
.B1(n_171),
.B2(n_200),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_193),
.A2(n_124),
.B1(n_107),
.B2(n_38),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_202),
.A2(n_23),
.B1(n_21),
.B2(n_38),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_183),
.B(n_2),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_6),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_209),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_279),
.Y(n_344)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_214),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_295),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_282),
.B(n_284),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_199),
.C(n_172),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_312),
.C(n_231),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_201),
.Y(n_284)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_209),
.B1(n_226),
.B2(n_179),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_287),
.A2(n_290),
.B1(n_270),
.B2(n_242),
.Y(n_339)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_189),
.B1(n_207),
.B2(n_190),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_291),
.Y(n_342)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_296),
.Y(n_349)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_297),
.B(n_306),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_298),
.B(n_310),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_299),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_236),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_307),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_303),
.Y(n_346)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_313),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_246),
.B(n_6),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_309),
.B(n_311),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_251),
.B(n_177),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_234),
.B(n_182),
.C(n_181),
.Y(n_312)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_235),
.A2(n_21),
.B1(n_23),
.B2(n_38),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_317),
.B1(n_320),
.B2(n_249),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_256),
.B(n_240),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_316),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_243),
.A2(n_233),
.B1(n_237),
.B2(n_253),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_258),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_321),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_232),
.B(n_21),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_322),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_7),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_234),
.B(n_7),
.Y(n_322)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_323),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_324),
.B(n_361),
.Y(n_396)
);

AOI32xp33_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_230),
.A3(n_261),
.B1(n_267),
.B2(n_262),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_283),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_305),
.A2(n_248),
.B1(n_244),
.B2(n_241),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_329),
.A2(n_338),
.B1(n_348),
.B2(n_350),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_340),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_244),
.B1(n_241),
.B2(n_260),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_343),
.B1(n_345),
.B2(n_354),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_254),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_254),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_359),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_294),
.A2(n_276),
.B1(n_275),
.B2(n_247),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_294),
.A2(n_285),
.B1(n_314),
.B2(n_302),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_315),
.A2(n_247),
.B1(n_271),
.B2(n_275),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_285),
.A2(n_242),
.B1(n_265),
.B2(n_277),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_281),
.A2(n_265),
.B1(n_273),
.B2(n_266),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_351),
.A2(n_287),
.B1(n_304),
.B2(n_296),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_290),
.A2(n_273),
.B1(n_266),
.B2(n_9),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_23),
.C(n_38),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_302),
.B(n_23),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_286),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_366),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_326),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_353),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_368),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_312),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_371),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_333),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_335),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_375),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_347),
.A2(n_281),
.B(n_322),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_373),
.A2(n_398),
.B(n_351),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_374),
.A2(n_390),
.B1(n_356),
.B2(n_332),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_321),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_378),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_288),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_380),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_342),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_383),
.Y(n_401)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_387),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_328),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_386),
.B(n_391),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_291),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_332),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_389),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_352),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_L g390 ( 
.A1(n_339),
.A2(n_304),
.B1(n_306),
.B2(n_297),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_328),
.B(n_298),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_394),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_278),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_393),
.Y(n_428)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_363),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_336),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_340),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_303),
.B(n_279),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_368),
.B(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_402),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_369),
.A2(n_324),
.B1(n_329),
.B2(n_338),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_404),
.A2(n_418),
.B1(n_427),
.B2(n_398),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_417),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_374),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_365),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_362),
.Y(n_416)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_369),
.A2(n_392),
.B1(n_394),
.B2(n_396),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_419),
.B(n_395),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_363),
.C(n_359),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_419),
.C(n_367),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_348),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_365),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_378),
.B(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_396),
.A2(n_362),
.B1(n_358),
.B2(n_361),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_429),
.A2(n_387),
.B1(n_382),
.B2(n_356),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_432),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_446),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_380),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_435),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_397),
.C(n_385),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_440),
.C(n_451),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_421),
.B(n_408),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_388),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_438),
.B(n_441),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_385),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_410),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_403),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_442),
.B(n_455),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_444),
.A2(n_445),
.B1(n_417),
.B2(n_413),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_427),
.A2(n_393),
.B1(n_373),
.B2(n_383),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_448),
.A2(n_452),
.B1(n_454),
.B2(n_422),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_391),
.C(n_376),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_428),
.A2(n_408),
.B1(n_429),
.B2(n_414),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_400),
.B(n_384),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_405),
.C(n_422),
.Y(n_466)
);

AOI211xp5_ASAP7_75t_L g454 ( 
.A1(n_428),
.A2(n_389),
.B(n_346),
.C(n_301),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_400),
.B(n_313),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_457),
.A2(n_406),
.B1(n_423),
.B2(n_407),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_421),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_458),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_443),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_463),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_445),
.A2(n_426),
.B(n_404),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_469),
.B(n_448),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_454),
.Y(n_463)
);

XOR2x2_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_416),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_466),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_467),
.A2(n_433),
.B1(n_452),
.B2(n_449),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_444),
.A2(n_409),
.B(n_401),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_474),
.Y(n_488)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_434),
.C(n_440),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_476),
.C(n_477),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_401),
.C(n_409),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_405),
.C(n_406),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_485),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_481),
.A2(n_457),
.B1(n_474),
.B2(n_472),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_453),
.C(n_446),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_465),
.C(n_456),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_468),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_490),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_469),
.A2(n_423),
.B1(n_407),
.B2(n_330),
.Y(n_489)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_489),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_470),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_463),
.A2(n_330),
.B1(n_307),
.B2(n_293),
.Y(n_491)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_462),
.A2(n_458),
.B(n_467),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_459),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_471),
.B(n_280),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_494),
.B(n_458),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_497),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_478),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_456),
.C(n_477),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_508),
.C(n_487),
.Y(n_509)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_466),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_501),
.A2(n_507),
.B(n_488),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_484),
.A2(n_476),
.B(n_473),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_505),
.A2(n_500),
.B(n_493),
.Y(n_513)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_484),
.Y(n_506)
);

CKINVDCx11_ASAP7_75t_R g511 ( 
.A(n_506),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_473),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_465),
.C(n_464),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_512),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_515),
.C(n_519),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_513),
.A2(n_503),
.B(n_508),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_502),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_514),
.A2(n_498),
.B1(n_492),
.B2(n_461),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_485),
.C(n_479),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_479),
.B1(n_486),
.B2(n_489),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_496),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_492),
.C(n_486),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_525),
.C(n_526),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_516),
.C(n_515),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_523),
.B(n_524),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_496),
.C(n_460),
.Y(n_525)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_511),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_530),
.B(n_517),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_521),
.C(n_513),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_532),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_512),
.B1(n_292),
.B2(n_323),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_531),
.B(n_528),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_8),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_533),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_537),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_538),
.B(n_10),
.Y(n_539)
);


endmodule