module real_aes_17125_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_0), .Y(n_556) );
AND2x4_ASAP7_75t_L g865 ( .A(n_1), .B(n_866), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_2), .A2(n_4), .B1(n_258), .B2(n_259), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_3), .A2(n_23), .B1(n_158), .B2(n_239), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_5), .A2(n_53), .B1(n_166), .B2(n_195), .Y(n_194) );
BUFx3_ASAP7_75t_L g590 ( .A(n_6), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_7), .A2(n_13), .B1(n_129), .B2(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g866 ( .A(n_8), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_9), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_10), .B(n_164), .Y(n_604) );
OR2x2_ASAP7_75t_L g110 ( .A(n_11), .B(n_33), .Y(n_110) );
BUFx2_ASAP7_75t_L g862 ( .A(n_11), .Y(n_862) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_12), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_14), .B(n_200), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_15), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_16), .B(n_173), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_17), .A2(n_86), .B1(n_200), .B2(n_239), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_18), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_19), .A2(n_59), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_19), .Y(n_114) );
INVx1_ASAP7_75t_L g847 ( .A(n_20), .Y(n_847) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_21), .A2(n_49), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_22), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_24), .B(n_158), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_25), .B(n_134), .Y(n_214) );
INVx4_ASAP7_75t_R g182 ( .A(n_26), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_27), .Y(n_848) );
AO32x2_ASAP7_75t_L g515 ( .A1(n_28), .A2(n_152), .A3(n_153), .B1(n_516), .B2(n_519), .Y(n_515) );
AO32x1_ASAP7_75t_L g620 ( .A1(n_28), .A2(n_152), .A3(n_153), .B1(n_516), .B2(n_519), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_29), .B(n_158), .Y(n_221) );
INVx1_ASAP7_75t_L g263 ( .A(n_30), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_SL g236 ( .A1(n_31), .A2(n_129), .B(n_133), .C(n_237), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_32), .A2(n_46), .B1(n_129), .B2(n_136), .Y(n_245) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_33), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_34), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_35), .A2(n_52), .B1(n_158), .B2(n_183), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_36), .A2(n_91), .B1(n_136), .B2(n_239), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_37), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_38), .B(n_528), .Y(n_532) );
INVx1_ASAP7_75t_L g218 ( .A(n_39), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_40), .B(n_129), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_41), .A2(n_68), .B1(n_136), .B2(n_541), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_42), .Y(n_156) );
INVx2_ASAP7_75t_L g105 ( .A(n_43), .Y(n_105) );
BUFx3_ASAP7_75t_L g109 ( .A(n_44), .Y(n_109) );
INVx1_ASAP7_75t_L g842 ( .A(n_44), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_45), .B(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_47), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_48), .A2(n_85), .B1(n_129), .B2(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_50), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_51), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_54), .A2(n_78), .B1(n_202), .B2(n_528), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_55), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_56), .A2(n_82), .B1(n_200), .B2(n_239), .Y(n_586) );
INVx1_ASAP7_75t_L g142 ( .A(n_57), .Y(n_142) );
AND2x4_ASAP7_75t_L g144 ( .A(n_58), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g115 ( .A(n_59), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_60), .A2(n_90), .B1(n_136), .B2(n_256), .Y(n_255) );
AO22x1_ASAP7_75t_L g198 ( .A1(n_61), .A2(n_73), .B1(n_199), .B2(n_201), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_62), .B(n_239), .Y(n_603) );
INVx1_ASAP7_75t_L g145 ( .A(n_63), .Y(n_145) );
AND2x2_ASAP7_75t_L g240 ( .A(n_64), .B(n_152), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_65), .B(n_152), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_66), .A2(n_166), .B(n_193), .C(n_555), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_67), .B(n_239), .C(n_607), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_69), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_70), .Y(n_231) );
AND2x2_ASAP7_75t_L g557 ( .A(n_71), .B(n_187), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_72), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_74), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_75), .A2(n_96), .B1(n_200), .B2(n_202), .Y(n_579) );
INVx2_ASAP7_75t_L g134 ( .A(n_76), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_77), .B(n_159), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_79), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_80), .B(n_152), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_81), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_83), .A2(n_102), .B1(n_856), .B2(n_867), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_84), .B(n_140), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_87), .B(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_88), .A2(n_100), .B1(n_136), .B2(n_183), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_89), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_92), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g506 ( .A(n_93), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_93), .B(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_94), .B(n_173), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_95), .A2(n_138), .B(n_166), .C(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g186 ( .A(n_97), .B(n_187), .Y(n_186) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_98), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_99), .Y(n_566) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_106), .B(n_834), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g837 ( .A(n_104), .Y(n_837) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_111), .B1(n_831), .B2(n_832), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g833 ( .A(n_108), .B(n_505), .Y(n_833) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
NOR3x1_ASAP7_75t_L g863 ( .A(n_109), .B(n_843), .C(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g844 ( .A(n_110), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_113), .B1(n_116), .B2(n_830), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g830 ( .A(n_116), .Y(n_830) );
AOI22x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_503), .B1(n_507), .B2(n_827), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
XNOR2x1_ASAP7_75t_L g845 ( .A(n_118), .B(n_846), .Y(n_845) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_412), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_328), .C(n_359), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_294), .Y(n_120) );
AOI211x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_206), .B(n_249), .C(n_280), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_170), .Y(n_123) );
AND2x2_ASAP7_75t_L g435 ( .A(n_124), .B(n_310), .Y(n_435) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_149), .Y(n_124) );
INVx1_ASAP7_75t_L g320 ( .A(n_125), .Y(n_320) );
OR2x2_ASAP7_75t_L g441 ( .A(n_125), .B(n_292), .Y(n_441) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g277 ( .A(n_126), .B(n_150), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_126), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g309 ( .A(n_126), .Y(n_309) );
OR2x2_ASAP7_75t_L g340 ( .A(n_126), .B(n_171), .Y(n_340) );
AND2x2_ASAP7_75t_L g354 ( .A(n_126), .B(n_171), .Y(n_354) );
AND2x2_ASAP7_75t_L g391 ( .A(n_126), .B(n_347), .Y(n_391) );
AO31x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_139), .A3(n_143), .B(n_146), .Y(n_126) );
OAI22x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B1(n_135), .B2(n_137), .Y(n_127) );
INVx4_ASAP7_75t_L g131 ( .A(n_129), .Y(n_131) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_130), .Y(n_164) );
INVx1_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
INVx1_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_130), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_130), .Y(n_202) );
INVx1_ASAP7_75t_L g233 ( .A(n_130), .Y(n_233) );
INVx2_ASAP7_75t_L g239 ( .A(n_130), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_131), .A2(n_156), .B(n_157), .C(n_159), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_132), .A2(n_192), .B1(n_244), .B2(n_245), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_132), .A2(n_137), .B1(n_255), .B2(n_257), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_132), .A2(n_532), .B(n_533), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_132), .A2(n_192), .B1(n_540), .B2(n_542), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_132), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_132), .A2(n_133), .B1(n_586), .B2(n_587), .Y(n_585) );
INVx6_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_163), .B(n_165), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_133), .B(n_198), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_133), .A2(n_191), .B(n_198), .C(n_204), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_133), .A2(n_235), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_133), .A2(n_603), .B(n_604), .Y(n_602) );
BUFx8_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g138 ( .A(n_134), .Y(n_138) );
INVx2_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
INVx1_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_136), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g258 ( .A(n_136), .Y(n_258) );
INVx2_ASAP7_75t_L g530 ( .A(n_136), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_137), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g553 ( .A(n_138), .Y(n_553) );
INVx1_ASAP7_75t_SL g578 ( .A(n_138), .Y(n_578) );
INVx2_ASAP7_75t_L g600 ( .A(n_139), .Y(n_600) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
OAI21xp33_ASAP7_75t_L g204 ( .A1(n_140), .A2(n_196), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
INVx2_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
BUFx10_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx10_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
INVx1_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx1_ASAP7_75t_L g261 ( .A(n_144), .Y(n_261) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_144), .A2(n_538), .A3(n_539), .B(n_543), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx2_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
BUFx2_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_148), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_148), .B(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_148), .B(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g271 ( .A(n_149), .Y(n_271) );
AND2x2_ASAP7_75t_L g322 ( .A(n_149), .B(n_188), .Y(n_322) );
AND2x2_ASAP7_75t_L g465 ( .A(n_149), .B(n_171), .Y(n_465) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g289 ( .A(n_150), .Y(n_289) );
AND2x2_ASAP7_75t_L g308 ( .A(n_150), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g345 ( .A(n_150), .Y(n_345) );
AND2x2_ASAP7_75t_L g369 ( .A(n_150), .B(n_171), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_154), .Y(n_150) );
NOR2x1_ASAP7_75t_L g167 ( .A(n_152), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g246 ( .A(n_152), .Y(n_246) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g222 ( .A(n_153), .B(n_169), .Y(n_222) );
INVx2_ASAP7_75t_SL g524 ( .A(n_153), .Y(n_524) );
BUFx3_ASAP7_75t_L g538 ( .A(n_153), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_153), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g563 ( .A(n_153), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_153), .B(n_589), .Y(n_588) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_162), .B(n_167), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_158), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g541 ( .A(n_158), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_158), .A2(n_183), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx2_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_160), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_164), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
INVx2_ASAP7_75t_L g256 ( .A(n_164), .Y(n_256) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_169), .A2(n_243), .A3(n_246), .B(n_247), .Y(n_242) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_169), .A2(n_565), .B(n_568), .Y(n_564) );
AOI31xp67_ASAP7_75t_L g584 ( .A1(n_169), .A2(n_246), .A3(n_585), .B(n_588), .Y(n_584) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_169), .A2(n_602), .B(n_605), .Y(n_601) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_170), .Y(n_269) );
AND2x2_ASAP7_75t_L g330 ( .A(n_170), .B(n_319), .Y(n_330) );
INVx2_ASAP7_75t_L g462 ( .A(n_170), .Y(n_462) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_188), .Y(n_170) );
INVx1_ASAP7_75t_L g267 ( .A(n_171), .Y(n_267) );
AND2x4_ASAP7_75t_L g279 ( .A(n_171), .B(n_189), .Y(n_279) );
INVx2_ASAP7_75t_L g347 ( .A(n_171), .Y(n_347) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_186), .Y(n_171) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_172), .A2(n_548), .B(n_557), .Y(n_547) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_180), .B(n_185), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx2_ASAP7_75t_L g195 ( .A(n_178), .Y(n_195) );
INVx1_ASAP7_75t_L g570 ( .A(n_183), .Y(n_570) );
AND2x2_ASAP7_75t_L g346 ( .A(n_188), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g353 ( .A(n_188), .Y(n_353) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g431 ( .A(n_189), .B(n_347), .Y(n_431) );
AOI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_197), .B(n_203), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_196), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_192), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_192), .A2(n_527), .B(n_529), .Y(n_526) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g534 ( .A(n_200), .Y(n_534) );
OAI21xp33_ASAP7_75t_SL g213 ( .A1(n_201), .A2(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_202), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_205), .A2(n_229), .B(n_236), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_205), .A2(n_549), .B(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_223), .Y(n_207) );
OR2x2_ASAP7_75t_L g336 ( .A(n_208), .B(n_224), .Y(n_336) );
AND2x2_ASAP7_75t_L g474 ( .A(n_208), .B(n_418), .Y(n_474) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x4_ASAP7_75t_L g251 ( .A(n_209), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g356 ( .A(n_209), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_209), .B(n_298), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_209), .B(n_274), .Y(n_411) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g268 ( .A(n_210), .Y(n_268) );
AND2x2_ASAP7_75t_L g284 ( .A(n_210), .B(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_SL g297 ( .A(n_210), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g305 ( .A(n_210), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_210), .B(n_274), .Y(n_376) );
AND2x2_ASAP7_75t_L g424 ( .A(n_210), .B(n_253), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_210), .B(n_252), .Y(n_467) );
BUFx2_ASAP7_75t_L g486 ( .A(n_210), .Y(n_486) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_222), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
INVx1_ASAP7_75t_L g607 ( .A(n_217), .Y(n_607) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g383 ( .A(n_224), .Y(n_383) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_241), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_225), .B(n_253), .Y(n_286) );
INVx2_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
AND2x2_ASAP7_75t_L g334 ( .A(n_225), .B(n_242), .Y(n_334) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
AOI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_240), .Y(n_226) );
AO31x2_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_254), .A3(n_260), .B(n_262), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_232), .B(n_235), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
O2A1O1Ixp5_ASAP7_75t_L g565 ( .A1(n_235), .A2(n_259), .B(n_566), .C(n_567), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_SL g528 ( .A(n_239), .Y(n_528) );
INVx1_ASAP7_75t_L g358 ( .A(n_241), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_241), .B(n_253), .Y(n_375) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g285 ( .A(n_242), .Y(n_285) );
OR2x2_ASAP7_75t_L g317 ( .A(n_242), .B(n_253), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_242), .B(n_253), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B1(n_272), .B2(n_276), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_264), .B1(n_268), .B2(n_269), .Y(n_250) );
INVx2_ASAP7_75t_L g275 ( .A(n_251), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_251), .B(n_334), .Y(n_348) );
AND2x2_ASAP7_75t_L g382 ( .A(n_251), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g300 ( .A(n_253), .Y(n_300) );
INVx1_ASAP7_75t_L g306 ( .A(n_253), .Y(n_306) );
AO31x2_ASAP7_75t_L g575 ( .A1(n_260), .A2(n_538), .A3(n_576), .B(n_580), .Y(n_575) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_SL g519 ( .A(n_261), .Y(n_519) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g440 ( .A(n_266), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g321 ( .A(n_267), .Y(n_321) );
AND3x1_ASAP7_75t_L g425 ( .A(n_267), .B(n_288), .C(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g381 ( .A(n_268), .Y(n_381) );
AND2x4_ASAP7_75t_L g417 ( .A(n_268), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g455 ( .A(n_271), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_272), .Y(n_459) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
OR2x2_ASAP7_75t_L g432 ( .A(n_273), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_273), .Y(n_480) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g380 ( .A(n_274), .B(n_358), .Y(n_380) );
AND2x2_ASAP7_75t_L g422 ( .A(n_274), .B(n_289), .Y(n_422) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_274), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_277), .B(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_277), .A2(n_278), .B(n_342), .C(n_348), .Y(n_341) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_277), .B(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_277), .B(n_435), .Y(n_481) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_279), .B(n_308), .Y(n_327) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_287), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_286), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_287), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
AND2x2_ASAP7_75t_L g337 ( .A(n_288), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_288), .B(n_354), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_288), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_288), .B(n_346), .Y(n_502) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g485 ( .A(n_289), .Y(n_485) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_307), .B(n_312), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_301), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OAI33xp33_ASAP7_75t_L g361 ( .A1(n_297), .A2(n_302), .A3(n_362), .B1(n_363), .B2(n_365), .B3(n_366), .Y(n_361) );
OR2x2_ASAP7_75t_L g493 ( .A(n_297), .B(n_317), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_297), .Y(n_495) );
INVx1_ASAP7_75t_L g316 ( .A(n_298), .Y(n_316) );
OR2x2_ASAP7_75t_L g357 ( .A(n_298), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_302), .B(n_484), .C(n_486), .Y(n_483) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_303), .B(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_303), .B(n_467), .Y(n_471) );
AND2x4_ASAP7_75t_L g500 ( .A(n_303), .B(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
OR2x2_ASAP7_75t_L g332 ( .A(n_305), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g445 ( .A(n_305), .B(n_380), .Y(n_445) );
INVx1_ASAP7_75t_L g501 ( .A(n_305), .Y(n_501) );
AND2x4_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_308), .Y(n_324) );
INVx1_ASAP7_75t_L g367 ( .A(n_309), .Y(n_367) );
AND2x2_ASAP7_75t_L g408 ( .A(n_309), .B(n_311), .Y(n_408) );
INVx1_ASAP7_75t_L g448 ( .A(n_310), .Y(n_448) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g339 ( .A(n_311), .B(n_340), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_318), .B1(n_325), .B2(n_327), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g404 ( .A(n_317), .Y(n_404) );
INVx2_ASAP7_75t_L g418 ( .A(n_317), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_322), .C(n_323), .Y(n_318) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_320), .B(n_345), .Y(n_447) );
OR2x2_ASAP7_75t_L g463 ( .A(n_320), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g476 ( .A(n_320), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_322), .B(n_390), .Y(n_451) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_349), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_335), .B2(n_337), .C(n_341), .Y(n_329) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI32xp33_ASAP7_75t_L g498 ( .A1(n_332), .A2(n_429), .A3(n_447), .B1(n_499), .B2(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g468 ( .A(n_334), .Y(n_468) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_337), .A2(n_350), .B(n_355), .Y(n_349) );
NAND2x1_ASAP7_75t_L g497 ( .A(n_338), .B(n_485), .Y(n_497) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AND2x2_ASAP7_75t_L g491 ( .A(n_344), .B(n_372), .Y(n_491) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g439 ( .A(n_345), .Y(n_439) );
INVx2_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
AND2x2_ASAP7_75t_L g368 ( .A(n_352), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_377), .C(n_388), .D(n_399), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_368), .B1(n_370), .B2(n_373), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_362), .A2(n_490), .B1(n_492), .B2(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g472 ( .A(n_367), .B(n_431), .Y(n_472) );
AND2x2_ASAP7_75t_L g475 ( .A(n_369), .B(n_476), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_389), .B1(n_393), .B2(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OR2x2_ASAP7_75t_L g410 ( .A(n_375), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g394 ( .A(n_376), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B(n_384), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_378), .A2(n_483), .B(n_487), .C(n_489), .Y(n_482) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g457 ( .A(n_380), .Y(n_457) );
AND2x4_ASAP7_75t_L g450 ( .A(n_383), .B(n_424), .Y(n_450) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_390), .A2(n_416), .B(n_419), .Y(n_415) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g421 ( .A(n_391), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_391), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g397 ( .A(n_395), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_428), .B1(n_432), .B2(n_434), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B1(n_406), .B2(n_409), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_404), .Y(n_420) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_477), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_436), .C(n_452), .D(n_469), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_427), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g479 ( .A(n_417), .B(n_480), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_423), .B2(n_425), .Y(n_419) );
INVxp67_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
BUFx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g433 ( .A(n_424), .Y(n_433) );
AND2x2_ASAP7_75t_L g456 ( .A(n_424), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_442), .B(n_444), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x6_ASAP7_75t_L g461 ( .A(n_439), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g458 ( .A(n_440), .Y(n_458) );
OAI32xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .A3(n_448), .B1(n_449), .B2(n_451), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .B1(n_458), .B2(n_459), .C(n_460), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B(n_466), .Y(n_460) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
INVx1_ASAP7_75t_L g488 ( .A(n_472), .Y(n_488) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
OAI211xp5_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_481), .B(n_482), .C(n_494), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_498), .Y(n_494) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
BUFx8_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_505), .Y(n_829) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g843 ( .A(n_506), .Y(n_843) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR2x1p5_ASAP7_75t_L g508 ( .A(n_509), .B(n_735), .Y(n_508) );
NAND4xp75_ASAP7_75t_L g509 ( .A(n_510), .B(n_632), .C(n_666), .D(n_715), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_558), .B(n_591), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g711 ( .A(n_514), .Y(n_711) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g596 ( .A(n_515), .B(n_522), .Y(n_596) );
AND2x4_ASAP7_75t_L g627 ( .A(n_515), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g648 ( .A(n_515), .Y(n_648) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_519), .A2(n_526), .B(n_531), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_520), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_536), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_521), .B(n_662), .Y(n_739) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_521), .Y(n_766) );
OR2x2_ASAP7_75t_L g815 ( .A(n_521), .B(n_619), .Y(n_815) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g631 ( .A(n_522), .Y(n_631) );
INVx3_ASAP7_75t_L g639 ( .A(n_522), .Y(n_639) );
OR2x2_ASAP7_75t_L g647 ( .A(n_522), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g675 ( .A(n_522), .B(n_645), .Y(n_675) );
INVx1_ASAP7_75t_L g686 ( .A(n_522), .Y(n_686) );
AND2x2_ASAP7_75t_L g707 ( .A(n_522), .B(n_648), .Y(n_707) );
INVxp67_ASAP7_75t_L g731 ( .A(n_522), .Y(n_731) );
BUFx2_ASAP7_75t_L g775 ( .A(n_522), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_522), .B(n_537), .Y(n_784) );
AND2x2_ASAP7_75t_L g791 ( .A(n_522), .B(n_792), .Y(n_791) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI21x1_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_535), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_530), .A2(n_606), .B(n_608), .Y(n_605) );
AND2x2_ASAP7_75t_L g649 ( .A(n_536), .B(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_536), .A2(n_561), .B1(n_765), .B2(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
OR2x2_ASAP7_75t_L g619 ( .A(n_537), .B(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g628 ( .A(n_537), .Y(n_628) );
AND2x2_ASAP7_75t_L g640 ( .A(n_537), .B(n_620), .Y(n_640) );
AND2x2_ASAP7_75t_L g698 ( .A(n_537), .B(n_546), .Y(n_698) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g595 ( .A(n_546), .Y(n_595) );
INVx1_ASAP7_75t_L g689 ( .A(n_546), .Y(n_689) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_546), .Y(n_792) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g645 ( .A(n_547), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_573), .Y(n_559) );
AND2x2_ASAP7_75t_L g746 ( .A(n_560), .B(n_692), .Y(n_746) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI32xp33_ASAP7_75t_L g776 ( .A1(n_561), .A2(n_669), .A3(n_743), .B1(n_777), .B2(n_779), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_561), .B(n_806), .Y(n_805) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g598 ( .A(n_562), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g615 ( .A(n_562), .B(n_575), .Y(n_615) );
BUFx2_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
INVx1_ASAP7_75t_L g681 ( .A(n_562), .Y(n_681) );
AND2x2_ASAP7_75t_L g714 ( .A(n_562), .B(n_693), .Y(n_714) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_572), .Y(n_562) );
OA21x2_ASAP7_75t_L g660 ( .A1(n_563), .A2(n_564), .B(n_572), .Y(n_660) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g597 ( .A(n_574), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g802 ( .A(n_574), .B(n_686), .Y(n_802) );
INVx1_ASAP7_75t_L g806 ( .A(n_574), .Y(n_806) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_582), .Y(n_574) );
INVx2_ASAP7_75t_L g630 ( .A(n_575), .Y(n_630) );
AND2x2_ASAP7_75t_L g654 ( .A(n_575), .B(n_613), .Y(n_654) );
AND2x2_ASAP7_75t_L g665 ( .A(n_575), .B(n_660), .Y(n_665) );
INVx1_ASAP7_75t_L g672 ( .A(n_575), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_575), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g693 ( .A(n_575), .Y(n_693) );
AND2x2_ASAP7_75t_L g759 ( .A(n_575), .B(n_582), .Y(n_759) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g623 ( .A(n_583), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g613 ( .A(n_584), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_597), .B1(n_610), .B2(n_616), .C(n_621), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_593), .A2(n_743), .B(n_746), .Y(n_742) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
AND2x4_ASAP7_75t_L g818 ( .A(n_594), .B(n_618), .Y(n_818) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g662 ( .A(n_595), .B(n_628), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_596), .B(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g727 ( .A(n_596), .Y(n_727) );
OR2x2_ASAP7_75t_L g671 ( .A(n_598), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g733 ( .A(n_598), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g804 ( .A(n_598), .Y(n_804) );
AND2x2_ASAP7_75t_L g612 ( .A(n_599), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g761 ( .A(n_599), .B(n_660), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_609), .Y(n_599) );
OAI21x1_ASAP7_75t_L g624 ( .A1(n_600), .A2(n_601), .B(n_609), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_610), .A2(n_642), .B1(n_643), .B2(n_652), .C(n_661), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_610), .A2(n_725), .B1(n_738), .B2(n_740), .C(n_742), .Y(n_737) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
AND2x2_ASAP7_75t_L g664 ( .A(n_612), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g677 ( .A(n_613), .B(n_660), .Y(n_677) );
INVx2_ASAP7_75t_L g683 ( .A(n_613), .Y(n_683) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g747 ( .A1(n_616), .A2(n_748), .B1(n_753), .B2(n_757), .C(n_762), .Y(n_747) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g799 ( .A(n_619), .B(n_769), .Y(n_799) );
INVx1_ASAP7_75t_L g651 ( .A(n_620), .Y(n_651) );
INVx1_ASAP7_75t_L g688 ( .A(n_620), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g637 ( .A(n_623), .Y(n_637) );
OR2x2_ASAP7_75t_L g700 ( .A(n_623), .B(n_636), .Y(n_700) );
INVx2_ASAP7_75t_L g713 ( .A(n_623), .Y(n_713) );
INVx2_ASAP7_75t_L g658 ( .A(n_624), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g663 ( .A(n_627), .Y(n_663) );
AND2x4_ASAP7_75t_L g669 ( .A(n_627), .B(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_627), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g743 ( .A(n_627), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g820 ( .A(n_627), .B(n_775), .Y(n_820) );
AND2x2_ASAP7_75t_L g644 ( .A(n_628), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g706 ( .A(n_628), .Y(n_706) );
INVx1_ASAP7_75t_L g765 ( .A(n_628), .Y(n_765) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx2_ASAP7_75t_SL g636 ( .A(n_630), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_630), .B(n_657), .Y(n_678) );
AND2x2_ASAP7_75t_L g752 ( .A(n_631), .B(n_706), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_638), .B(n_641), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g718 ( .A(n_634), .Y(n_718) );
AND2x2_ASAP7_75t_L g785 ( .A(n_634), .B(n_713), .Y(n_785) );
AND2x2_ASAP7_75t_L g800 ( .A(n_634), .B(n_759), .Y(n_800) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx2_ASAP7_75t_L g754 ( .A(n_636), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_636), .B(n_761), .Y(n_771) );
OAI33xp33_ASAP7_75t_L g808 ( .A1(n_636), .A2(n_710), .A3(n_778), .B1(n_809), .B2(n_810), .B3(n_811), .Y(n_808) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_639), .B(n_645), .Y(n_769) );
AND2x2_ASAP7_75t_L g797 ( .A(n_640), .B(n_745), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g670 ( .A(n_645), .Y(n_670) );
INVx1_ASAP7_75t_L g745 ( .A(n_645), .Y(n_745) );
OAI32xp33_ASAP7_75t_L g690 ( .A1(n_646), .A2(n_671), .A3(n_691), .B1(n_694), .B2(n_696), .Y(n_690) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g725 ( .A(n_647), .B(n_670), .Y(n_725) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g703 ( .A(n_651), .Y(n_703) );
INVx2_ASAP7_75t_L g751 ( .A(n_651), .Y(n_751) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g734 ( .A(n_654), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_655), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g794 ( .A(n_655), .B(n_741), .Y(n_794) );
INVx2_ASAP7_75t_L g825 ( .A(n_655), .Y(n_825) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g740 ( .A(n_656), .B(n_741), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
AND2x2_ASAP7_75t_L g682 ( .A(n_657), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g724 ( .A(n_658), .Y(n_724) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B(n_664), .Y(n_661) );
INVx2_ASAP7_75t_L g732 ( .A(n_662), .Y(n_732) );
AND2x2_ASAP7_75t_L g716 ( .A(n_663), .B(n_717), .Y(n_716) );
NOR3x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_690), .C(n_699), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_671), .B(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_670), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_672), .B(n_723), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B1(n_679), .B2(n_684), .Y(n_673) );
INVx3_ASAP7_75t_L g708 ( .A(n_675), .Y(n_708) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVxp67_ASAP7_75t_L g721 ( .A(n_677), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_677), .B(n_756), .Y(n_755) );
AND2x4_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
AND2x2_ASAP7_75t_L g822 ( .A(n_680), .B(n_713), .Y(n_822) );
AND2x2_ASAP7_75t_L g692 ( .A(n_683), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g741 ( .A(n_683), .Y(n_741) );
INVx1_ASAP7_75t_L g778 ( .A(n_683), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_683), .B(n_724), .Y(n_812) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g809 ( .A(n_687), .Y(n_809) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g695 ( .A(n_689), .Y(n_695) );
AND2x2_ASAP7_75t_L g821 ( .A(n_692), .B(n_761), .Y(n_821) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
BUFx2_ASAP7_75t_L g729 ( .A(n_698), .Y(n_729) );
AND2x2_ASAP7_75t_L g826 ( .A(n_698), .B(n_707), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_709), .B2(n_712), .Y(n_699) );
AOI211xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_704), .B(n_707), .C(n_708), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g783 ( .A(n_703), .B(n_784), .Y(n_783) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp33_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
AND2x2_ASAP7_75t_L g717 ( .A(n_713), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g795 ( .A(n_714), .B(n_756), .Y(n_795) );
INVx1_ASAP7_75t_L g810 ( .A(n_714), .Y(n_810) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .C(n_726), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_725), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g756 ( .A(n_724), .Y(n_756) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B(n_730), .C(n_733), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_727), .A2(n_820), .B1(n_821), .B2(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_787), .Y(n_735) );
NOR3xp33_ASAP7_75t_SL g736 ( .A(n_737), .B(n_747), .C(n_772), .Y(n_736) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_743), .A2(n_782), .B1(n_785), .B2(n_786), .Y(n_781) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
AND2x2_ASAP7_75t_L g767 ( .A(n_750), .B(n_768), .Y(n_767) );
AND2x4_ASAP7_75t_L g790 ( .A(n_750), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g786 ( .A(n_755), .Y(n_786) );
OR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_761), .B(n_778), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_767), .B(n_770), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_767), .A2(n_822), .B1(n_824), .B2(n_826), .Y(n_823) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI21xp33_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_776), .B(n_781), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_774), .B(n_818), .Y(n_817) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g813 ( .A(n_784), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_786), .A2(n_808), .B1(n_813), .B2(n_814), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_816), .Y(n_787) );
OAI211xp5_ASAP7_75t_SL g788 ( .A1(n_789), .A2(n_793), .B(n_796), .C(n_807), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
O2A1O1Ixp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B(n_800), .C(n_801), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_799), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_801) );
OAI211xp5_ASAP7_75t_L g816 ( .A1(n_810), .A2(n_817), .B(n_819), .C(n_823), .Y(n_816) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx8_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
BUFx12f_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
OAI21xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_838), .B(n_849), .Y(n_834) );
INVxp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_845), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AND3x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .C(n_844), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g854 ( .A(n_842), .Y(n_854) );
AND2x6_ASAP7_75t_SL g852 ( .A(n_844), .B(n_853), .Y(n_852) );
XOR2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_855), .Y(n_850) );
INVx5_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
INVx4_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
CKINVDCx14_ASAP7_75t_R g867 ( .A(n_858), .Y(n_867) );
AND2x6_ASAP7_75t_L g858 ( .A(n_859), .B(n_863), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
INVx2_ASAP7_75t_SL g864 ( .A(n_865), .Y(n_864) );
endmodule