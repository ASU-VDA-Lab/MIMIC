module fake_jpeg_15325_n_152 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_53),
.B1(n_64),
.B2(n_49),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_81),
.B1(n_84),
.B2(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_53),
.B1(n_64),
.B2(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_61),
.B1(n_58),
.B2(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_98),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_97),
.B1(n_103),
.B2(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_95),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_76),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_96),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_58),
.B1(n_47),
.B2(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_106),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_56),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_54),
.B(n_63),
.C(n_62),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_51),
.B1(n_22),
.B2(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_1),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_21),
.B1(n_44),
.B2(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_3),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_101),
.B1(n_102),
.B2(n_10),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_89),
.C(n_90),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_115),
.B1(n_97),
.B2(n_106),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_121),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_117),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_121),
.A2(n_123),
.B(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_28),
.B1(n_42),
.B2(n_41),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_110),
.B1(n_108),
.B2(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_8),
.B(n_9),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_120),
.C(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_108),
.B1(n_111),
.B2(n_10),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_29),
.CI(n_39),
.CON(n_138),
.SN(n_138)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_132),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_133),
.B1(n_9),
.B2(n_12),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_25),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_136),
.B(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.C(n_19),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_138),
.B(n_137),
.Y(n_142)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_30),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_35),
.B1(n_45),
.B2(n_14),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_144),
.C(n_18),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_38),
.B(n_15),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_16),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_36),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_37),
.B(n_12),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_13),
.Y(n_152)
);


endmodule