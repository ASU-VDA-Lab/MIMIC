module real_jpeg_15384_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_0),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_0),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_0),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_0),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_0),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_0),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_1),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_1),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_1),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_1),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_1),
.B(n_367),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_2),
.Y(n_120)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_3),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_4),
.B(n_111),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_4),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_54),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_5),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_7),
.B1(n_39),
.B2(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_7),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_7),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_7),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_7),
.B(n_354),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_8),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_8),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_8),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_8),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_8),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_8),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_8),
.B(n_313),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_11),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_11),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_11),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_13),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_13),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_13),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_13),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_13),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_13),
.B(n_258),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_13),
.B(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g204 ( 
.A(n_14),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_14),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_14),
.Y(n_352)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_15),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_220),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_218),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_169),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_19),
.B(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.C(n_143),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_21),
.A2(n_22),
.B1(n_100),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_23),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.C(n_49),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_24),
.B(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_29),
.C(n_33),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_30),
.Y(n_264)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_33),
.B(n_201),
.Y(n_253)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_35),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_36),
.B(n_201),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_37),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_389)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_38),
.A2(n_277),
.B(n_283),
.Y(n_276)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_43),
.Y(n_151)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_46),
.Y(n_190)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_59),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_51),
.B(n_59),
.Y(n_146)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_56),
.B(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_58),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_75),
.B1(n_97),
.B2(n_98),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_74),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_67),
.B(n_74),
.C(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_69),
.Y(n_260)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_71),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B(n_83),
.C(n_94),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_76),
.A2(n_80),
.B1(n_95),
.B2(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_79),
.Y(n_338)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_83),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_92),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_84),
.A2(n_92),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_84),
.Y(n_288)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_88),
.B(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_92),
.B(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_92),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_97),
.B(n_171),
.C(n_172),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_100),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_114),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_101),
.B(n_115),
.C(n_141),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_102),
.B(n_107),
.C(n_110),
.Y(n_191)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_109),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_130),
.B1(n_141),
.B2(n_142),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_126),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_117),
.B1(n_126),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_122),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_125),
.Y(n_309)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_136),
.C(n_140),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_132),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_132),
.B(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_136),
.A2(n_137),
.B1(n_149),
.B2(n_150),
.Y(n_232)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_138),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_140),
.B1(n_201),
.B2(n_205),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_138),
.B(n_262),
.Y(n_320)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_139),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_139),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_140),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_143),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_161),
.C(n_166),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_144),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_152),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_145),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_147),
.A2(n_148),
.B1(n_152),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_152),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_159),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_153),
.A2(n_159),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_153),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_155),
.B(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_157),
.Y(n_336)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_162),
.B(n_167),
.Y(n_386)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_194),
.B1(n_216),
.B2(n_217),
.Y(n_173)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_193),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_192),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_206),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_382),
.B(n_397),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_290),
.B(n_381),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_265),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_224),
.B(n_265),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_242),
.C(n_254),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_225),
.A2(n_226),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_232),
.C(n_233),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_240),
.Y(n_325)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_237),
.B(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_242),
.B(n_254),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_248),
.B1(n_249),
.B2(n_252),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_252),
.C(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.C(n_261),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_261),
.B(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_267),
.B(n_272),
.C(n_273),
.Y(n_391)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_274),
.B(n_276),
.C(n_286),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_375),
.B(n_380),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_329),
.B(n_374),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_321),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_293),
.B(n_321),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_310),
.C(n_319),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_294),
.A2(n_295),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_305),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_303),
.C(n_305),
.Y(n_323)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_319),
.B1(n_320),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_324),
.C(n_326),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_343),
.B(n_373),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_339),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_331),
.B(n_339),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.C(n_337),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_333),
.A2(n_334),
.B1(n_337),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_337),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_340),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_358),
.B(n_372),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_355),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_345),
.B(n_355),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_353),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_353),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_362),
.B(n_371),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_360),
.B(n_361),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_376),
.B(n_377),
.Y(n_380)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_391),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_391),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_388),
.C(n_390),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

OAI21x1_ASAP7_75t_SL g397 ( 
.A1(n_392),
.A2(n_398),
.B(n_399),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_394),
.Y(n_399)
);


endmodule