module fake_netlist_6_3446_n_187 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_187);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_187;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_186;
wire n_87;
wire n_32;
wire n_85;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_66;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_155;
wire n_29;
wire n_62;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_171;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVxp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVxp33_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_16),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2x1p5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_33),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_52),
.B1(n_55),
.B2(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

OAI221xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_50),
.B1(n_47),
.B2(n_38),
.C(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

OR2x6_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_36),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_34),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_36),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_80),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_68),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_69),
.B1(n_65),
.B2(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_86),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_88),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_88),
.B(n_86),
.C(n_64),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_80),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_75),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_95),
.B(n_96),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_84),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_97),
.Y(n_113)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_101),
.B(n_99),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_101),
.B(n_99),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_84),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

NOR2x1p5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_106),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

AOI31xp33_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_112),
.A3(n_116),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_117),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AOI21x1_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_114),
.B(n_115),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_104),
.B(n_116),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_116),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_123),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_127),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_87),
.B1(n_89),
.B2(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_127),
.B1(n_107),
.B2(n_33),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_127),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_34),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_57),
.C(n_85),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_130),
.C(n_125),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_89),
.B(n_87),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_111),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND3x1_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_5),
.C(n_7),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_111),
.B(n_130),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.C(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_67),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_115),
.B(n_111),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_8),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_8),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_142),
.B(n_63),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_67),
.Y(n_168)
);

NAND3x1_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_10),
.C(n_11),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_168),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_63),
.B(n_62),
.C(n_56),
.Y(n_172)
);

NOR3x1_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_114),
.C(n_83),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_114),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_125),
.B1(n_126),
.B2(n_66),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_68),
.C(n_66),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_64),
.Y(n_177)
);

OAI211xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_164),
.B(n_53),
.C(n_56),
.Y(n_178)
);

AOI211xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_176),
.B(n_172),
.C(n_170),
.Y(n_179)
);

NOR2x1p5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_169),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_63),
.B(n_53),
.C(n_62),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_53),
.C(n_62),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_175),
.B1(n_113),
.B2(n_71),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_178),
.B1(n_181),
.B2(n_71),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_113),
.B1(n_70),
.B2(n_93),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_185),
.B1(n_70),
.B2(n_113),
.C(n_93),
.Y(n_187)
);


endmodule