module fake_jpeg_22686_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_47),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_53),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_34),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_67),
.B(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_55),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_62),
.B1(n_74),
.B2(n_27),
.Y(n_93)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_57),
.B(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_41),
.B(n_47),
.C(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_17),
.B1(n_22),
.B2(n_31),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_30),
.B1(n_27),
.B2(n_32),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_31),
.C(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_34),
.B1(n_25),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_72),
.B1(n_33),
.B2(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_27),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_34),
.B1(n_25),
.B2(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_0),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_88),
.Y(n_120)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_93),
.B1(n_110),
.B2(n_50),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_13),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_61),
.C(n_67),
.Y(n_115)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_58),
.B1(n_65),
.B2(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_12),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_12),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_58),
.Y(n_127)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_52),
.B(n_13),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_113),
.B(n_14),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_13),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_49),
.B(n_11),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_14),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_45),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_63),
.A2(n_10),
.B1(n_8),
.B2(n_15),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_50),
.B(n_10),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_126),
.B1(n_132),
.B2(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_51),
.B1(n_81),
.B2(n_106),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_63),
.B(n_55),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_124),
.B1(n_111),
.B2(n_103),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_95),
.B1(n_102),
.B2(n_94),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_58),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_139),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_79),
.A2(n_65),
.B1(n_51),
.B2(n_57),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_65),
.B1(n_75),
.B2(n_51),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_79),
.B(n_87),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_10),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_138),
.B(n_0),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_36),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_135),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_158),
.B(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_119),
.B1(n_118),
.B2(n_115),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_152),
.B1(n_175),
.B2(n_124),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_82),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_96),
.B1(n_91),
.B2(n_89),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_87),
.C(n_83),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_8),
.C(n_36),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_92),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_90),
.CI(n_83),
.CON(n_155),
.SN(n_155)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_160),
.B(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_90),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_157),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_111),
.Y(n_157)
);

XOR2x2_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_133),
.B1(n_45),
.B2(n_18),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_1),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_88),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_16),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_14),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_85),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_142),
.B(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_78),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_138),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_120),
.A2(n_111),
.B1(n_18),
.B2(n_24),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_122),
.B(n_117),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_179),
.B(n_180),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_122),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_145),
.B(n_173),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_172),
.B(n_153),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_185),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_122),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_197),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_166),
.A2(n_142),
.B1(n_128),
.B2(n_121),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_203),
.B1(n_204),
.B2(n_163),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_84),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_164),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_45),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_146),
.A2(n_128),
.B1(n_133),
.B2(n_54),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_161),
.B(n_156),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_152),
.B1(n_159),
.B2(n_150),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_214),
.B1(n_216),
.B2(n_229),
.Y(n_233)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_190),
.A2(n_159),
.B1(n_148),
.B2(n_155),
.Y(n_214)
);

AOI32xp33_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_183),
.A3(n_189),
.B1(n_206),
.B2(n_186),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_155),
.B1(n_151),
.B2(n_157),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_179),
.A2(n_162),
.B1(n_165),
.B2(n_18),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_197),
.C(n_185),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_234),
.C(n_241),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_196),
.C(n_202),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_207),
.B(n_176),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_248),
.B(n_249),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_176),
.B1(n_178),
.B2(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_213),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_191),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_198),
.C(n_182),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_195),
.B1(n_181),
.B2(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_1),
.B(n_3),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_225),
.B(n_229),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_224),
.B1(n_223),
.B2(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_210),
.B(n_209),
.C(n_217),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_260),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_1),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_36),
.B1(n_32),
.B2(n_24),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_237),
.Y(n_269)
);

NAND2x1_ASAP7_75t_SL g260 ( 
.A(n_243),
.B(n_3),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_24),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_246),
.C(n_241),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_239),
.C(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_238),
.C(n_235),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_235),
.C(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_251),
.C(n_249),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_251),
.B(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_274),
.C(n_278),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_253),
.B1(n_256),
.B2(n_233),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_230),
.C(n_259),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.C(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_260),
.C(n_5),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_4),
.B(n_6),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_282),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_266),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_4),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_272),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_279),
.A3(n_281),
.B1(n_283),
.B2(n_273),
.C1(n_4),
.C2(n_6),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_287),
.B(n_7),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_285),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_291),
.Y(n_292)
);


endmodule