module fake_ibex_1915_n_4733 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_848, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4733);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4733;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_4688;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4687;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4364;
wire n_4204;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_4632;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_3838;
wire n_957;
wire n_4514;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_4668;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_4731;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_4142;
wire n_2322;
wire n_1233;
wire n_3025;
wire n_2335;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_4239;
wire n_3175;
wire n_3729;
wire n_4169;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4708;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_4673;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_4690;
wire n_1668;
wire n_3982;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_4672;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_3711;
wire n_1595;
wire n_2164;
wire n_4267;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_4723;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_4312;
wire n_4567;
wire n_917;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4430;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4223;
wire n_2260;
wire n_3977;
wire n_4724;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_4721;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_3822;
wire n_1276;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_4667;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_4711;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_4671;
wire n_1326;
wire n_971;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_4676;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_4714;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_3199;
wire n_1616;
wire n_2723;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4732;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_4692;
wire n_4713;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2646;
wire n_2387;
wire n_3375;
wire n_3241;
wire n_1121;
wire n_2397;
wire n_2746;
wire n_4615;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_4710;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_4680;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_4693;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4549;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_4700;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4523;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_4712;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_3626;
wire n_1831;
wire n_3733;
wire n_864;
wire n_1987;
wire n_4571;
wire n_959;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_4725;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4681;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3529;
wire n_1711;
wire n_3222;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_4033;
wire n_3855;
wire n_4485;
wire n_4608;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_3364;
wire n_1236;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_2999;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2910;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_4706;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_2699;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4674;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4679;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_1395;
wire n_998;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4660;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_4664;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_4709;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3646;
wire n_3477;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_4683;
wire n_3557;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_3398;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_4694;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_4717;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_4719;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_4685;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_4716;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_3284;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_4185;
wire n_2422;
wire n_3927;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_3314;
wire n_2997;
wire n_961;
wire n_1349;
wire n_1331;
wire n_991;
wire n_1223;
wire n_2127;
wire n_3891;
wire n_1323;
wire n_1739;
wire n_4704;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1601;
wire n_1294;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_4707;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_4695;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_4638;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_3356;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_4149;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_3930;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_4637;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_3773;
wire n_2528;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_3506;
wire n_2845;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_2732;
wire n_3162;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_4697;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_4730;
wire n_1415;
wire n_1238;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_4720;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_4715;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_4698;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_3604;
wire n_1740;
wire n_1989;
wire n_3649;
wire n_1838;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2576;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4200;
wire n_4111;
wire n_4162;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_4666;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_4663;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_4611;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2816;
wire n_2433;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_4670;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1542;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_4696;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_3368;
wire n_3561;
wire n_956;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_4729;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3173;
wire n_2872;
wire n_3102;
wire n_4345;
wire n_4281;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_4675;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_3163;
wire n_2701;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1912;
wire n_1297;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3791;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_4686;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4682;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_4705;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_4684;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_3296;
wire n_1911;
wire n_2293;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_1193;
wire n_3067;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_1074;
wire n_3380;
wire n_3225;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4718;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_4412;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_3286;
wire n_999;
wire n_2634;
wire n_2982;
wire n_4038;
wire n_1092;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1027;
wire n_1516;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_4448;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_4727;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_4701;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_4726;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_4544;
wire n_4728;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_4275;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_4689;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_4702;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2619;
wire n_3873;
wire n_3738;
wire n_4506;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1947;
wire n_1675;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_856;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_4703;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_4691;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_4662;
wire n_2658;

INVx1_ASAP7_75t_L g853 ( 
.A(n_557),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_606),
.Y(n_854)
);

CKINVDCx16_ASAP7_75t_R g855 ( 
.A(n_146),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_705),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_475),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_520),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_144),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_344),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_526),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_113),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_215),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_807),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_243),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_173),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_332),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_507),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_14),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_131),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_788),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_827),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_304),
.Y(n_873)
);

CKINVDCx16_ASAP7_75t_R g874 ( 
.A(n_264),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_42),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_523),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_210),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_341),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_16),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_819),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_570),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_201),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_500),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_503),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_747),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_583),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_782),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_830),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_727),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_673),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_509),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_726),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_614),
.Y(n_893)
);

BUFx10_ASAP7_75t_L g894 ( 
.A(n_340),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_485),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_238),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_118),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_468),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_711),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_482),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_39),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_507),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_167),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_787),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_561),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_543),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_606),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_390),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_688),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_786),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_812),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_499),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_460),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_808),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_587),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_844),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_303),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_408),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_270),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_790),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_845),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_794),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_109),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_710),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_738),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_113),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_126),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_776),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_753),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_657),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_469),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_175),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_452),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_775),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_778),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_842),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_804),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_652),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_48),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_284),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_825),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_750),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_260),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_824),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_822),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_457),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_116),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_568),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_221),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_277),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_223),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_803),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_82),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_383),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_793),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_640),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_612),
.Y(n_957)
);

BUFx10_ASAP7_75t_L g958 ( 
.A(n_634),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_228),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_628),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_445),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_653),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_485),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_100),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_372),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_668),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_605),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_558),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_798),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_842),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_411),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_471),
.Y(n_972)
);

CKINVDCx14_ASAP7_75t_R g973 ( 
.A(n_24),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_564),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_453),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_536),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_818),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_532),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_291),
.Y(n_979)
);

CKINVDCx14_ASAP7_75t_R g980 ( 
.A(n_174),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_516),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_624),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_700),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_772),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_478),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_728),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_437),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_142),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_720),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_702),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_832),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_635),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_740),
.Y(n_993)
);

HB1xp67_ASAP7_75t_SL g994 ( 
.A(n_355),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_427),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_458),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_425),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_489),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_246),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_275),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_851),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_267),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_640),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_455),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_719),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_64),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_791),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_329),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_30),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_799),
.Y(n_1010)
);

CKINVDCx14_ASAP7_75t_R g1011 ( 
.A(n_69),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_80),
.Y(n_1012)
);

BUFx8_ASAP7_75t_SL g1013 ( 
.A(n_577),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_267),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_311),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_416),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_419),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_61),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_482),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_355),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_565),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_42),
.Y(n_1022)
);

CKINVDCx16_ASAP7_75t_R g1023 ( 
.A(n_454),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_443),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_731),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_623),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_351),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_168),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_716),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_667),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_340),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_537),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_611),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_538),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_747),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_736),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_411),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_62),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_585),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_119),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_472),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_510),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_36),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_809),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_563),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_409),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_116),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_818),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_279),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_264),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_761),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_477),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_139),
.Y(n_1053)
);

CKINVDCx16_ASAP7_75t_R g1054 ( 
.A(n_629),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_774),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_715),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_102),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_801),
.Y(n_1058)
);

BUFx5_ASAP7_75t_L g1059 ( 
.A(n_526),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_734),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_220),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_851),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_723),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_221),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_830),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_758),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_658),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_533),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_153),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_240),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_800),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_387),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_820),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_795),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_28),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_784),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_554),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_364),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_627),
.Y(n_1079)
);

CKINVDCx16_ASAP7_75t_R g1080 ( 
.A(n_326),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_440),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_199),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_551),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_588),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_600),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_217),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_813),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_468),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_228),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_669),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_736),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_803),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_128),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_564),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_558),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_476),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_635),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_541),
.Y(n_1098)
);

BUFx2_ASAP7_75t_SL g1099 ( 
.A(n_583),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_790),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_843),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_708),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_431),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_729),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_143),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_273),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_143),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_317),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_791),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_327),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_428),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_787),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_773),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_587),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_838),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_658),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_814),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_281),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_493),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_777),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_802),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_287),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_712),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_529),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_33),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_29),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_778),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_797),
.Y(n_1128)
);

CKINVDCx14_ASAP7_75t_R g1129 ( 
.A(n_178),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_106),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_197),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_764),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_5),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_243),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_475),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_380),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_819),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_721),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_302),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_427),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_609),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_415),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_614),
.Y(n_1143)
);

CKINVDCx14_ASAP7_75t_R g1144 ( 
.A(n_179),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_62),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_275),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_65),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_786),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_142),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_810),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_160),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_383),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_795),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_202),
.Y(n_1154)
);

BUFx5_ASAP7_75t_L g1155 ( 
.A(n_809),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_432),
.Y(n_1156)
);

BUFx10_ASAP7_75t_L g1157 ( 
.A(n_91),
.Y(n_1157)
);

BUFx5_ASAP7_75t_L g1158 ( 
.A(n_429),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_254),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_442),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_767),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_530),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_780),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_682),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_56),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_829),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_574),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_495),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_234),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_222),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_607),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_40),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_687),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_582),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_484),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_821),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_377),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_435),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_586),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_378),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_554),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_685),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_63),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_282),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_561),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_196),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_282),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_204),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_815),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_205),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_833),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_665),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_805),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_653),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_647),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_792),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_806),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_241),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_664),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_121),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_705),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_607),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_651),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_428),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_356),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_114),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_111),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_811),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_612),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_367),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_556),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_823),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_779),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_401),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_813),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_42),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_299),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_47),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_518),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_668),
.Y(n_1220)
);

BUFx2_ASAP7_75t_SL g1221 ( 
.A(n_308),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_416),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_194),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_670),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_104),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_796),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_715),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_512),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_513),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_817),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_710),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_499),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_534),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_577),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_762),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_222),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_281),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_829),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_104),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_364),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_148),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_783),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_531),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_164),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_288),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_388),
.Y(n_1246)
);

INVxp33_ASAP7_75t_SL g1247 ( 
.A(n_158),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_93),
.Y(n_1248)
);

CKINVDCx16_ASAP7_75t_R g1249 ( 
.A(n_127),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_207),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_845),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_525),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_248),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_597),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_832),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_458),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_70),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_555),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_828),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_263),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_167),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_514),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_530),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_58),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_313),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_604),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_337),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_75),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_190),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_374),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_65),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_681),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_744),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_55),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_588),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_804),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_477),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_666),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_444),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_816),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_602),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_570),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_538),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_618),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_382),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_352),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_11),
.Y(n_1287)
);

BUFx10_ASAP7_75t_L g1288 ( 
.A(n_553),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_469),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_160),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_186),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_50),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_78),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_651),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_504),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_50),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_831),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_626),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_509),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_402),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_112),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_168),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_233),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_628),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_445),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_841),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_474),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_785),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_180),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_781),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_123),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_178),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_305),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_517),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_191),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_463),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_146),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_339),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_220),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_806),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_757),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_522),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_50),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_30),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_158),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_38),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_90),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_695),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_609),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_278),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_714),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_45),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_835),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_215),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_208),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_193),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_254),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_333),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_70),
.Y(n_1339)
);

BUFx2_ASAP7_75t_SL g1340 ( 
.A(n_122),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_180),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_699),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_734),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_48),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_274),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_10),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_449),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_592),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_139),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_81),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_374),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_181),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_756),
.Y(n_1353)
);

BUFx10_ASAP7_75t_L g1354 ( 
.A(n_339),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_13),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_43),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_500),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_789),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_601),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1018),
.B(n_0),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_894),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_902),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_888),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1247),
.B(n_0),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_888),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_872),
.B(n_0),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1247),
.B(n_1),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_894),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_967),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_967),
.Y(n_1370)
);

INVx5_ASAP7_75t_L g1371 ( 
.A(n_967),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1018),
.B(n_1),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1059),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_901),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1059),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1059),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_902),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_904),
.B(n_1),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_894),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1142),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1059),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_973),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1142),
.B(n_2),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_973),
.B(n_2),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_924),
.B(n_997),
.Y(n_1385)
);

INVxp33_ASAP7_75t_SL g1386 ( 
.A(n_961),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1228),
.B(n_2),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1059),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_901),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1289),
.B(n_3),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_902),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1170),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_958),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_902),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_980),
.B(n_3),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_958),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_980),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_977),
.Y(n_1398)
);

AND2x6_ASAP7_75t_L g1399 ( 
.A(n_977),
.B(n_3),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_984),
.B(n_4),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1059),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1011),
.B(n_4),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_925),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_925),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1132),
.B(n_4),
.Y(n_1405)
);

INVx5_ASAP7_75t_L g1406 ( 
.A(n_901),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_901),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1324),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_925),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_958),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1157),
.Y(n_1411)
);

BUFx12f_ASAP7_75t_L g1412 ( 
.A(n_1157),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1157),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1253),
.B(n_5),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1303),
.B(n_5),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1315),
.B(n_7),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_925),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_887),
.B(n_6),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1011),
.B(n_1129),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1182),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1059),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1155),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_928),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1182),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1170),
.B(n_6),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_899),
.B(n_6),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1201),
.B(n_7),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1129),
.B(n_7),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_928),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_928),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1217),
.B(n_8),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_928),
.Y(n_1432)
);

INVx5_ASAP7_75t_L g1433 ( 
.A(n_1324),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1251),
.B(n_8),
.Y(n_1434)
);

AND2x6_ASAP7_75t_L g1435 ( 
.A(n_1141),
.B(n_8),
.Y(n_1435)
);

BUFx8_ASAP7_75t_SL g1436 ( 
.A(n_875),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1284),
.B(n_9),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1182),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_960),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1185),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1144),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1347),
.B(n_9),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1155),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1144),
.B(n_9),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1185),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1284),
.B(n_10),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1185),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1237),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_960),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1155),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1155),
.Y(n_1451)
);

INVx5_ASAP7_75t_L g1452 ( 
.A(n_1324),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1141),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1181),
.B(n_10),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1181),
.B(n_11),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_960),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_960),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1155),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1074),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1186),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_855),
.B(n_11),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_869),
.B(n_12),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1074),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1074),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1324),
.Y(n_1465)
);

AND2x6_ASAP7_75t_L g1466 ( 
.A(n_1186),
.B(n_12),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_939),
.B(n_12),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1383),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1368),
.B(n_1099),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1416),
.A2(n_889),
.B1(n_917),
.B2(n_874),
.Y(n_1470)
);

BUFx10_ASAP7_75t_L g1471 ( 
.A(n_1383),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1386),
.A2(n_879),
.B1(n_1133),
.B2(n_875),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1425),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1366),
.A2(n_994),
.B1(n_1054),
.B2(n_1023),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1382),
.B(n_1397),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1441),
.B(n_1080),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1419),
.B(n_1123),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_R g1478 ( 
.A1(n_1436),
.A2(n_975),
.B1(n_987),
.B2(n_945),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1411),
.B(n_1221),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1385),
.A2(n_1249),
.B1(n_1301),
.B2(n_1138),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1363),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1378),
.A2(n_1038),
.B1(n_1043),
.B2(n_1009),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1387),
.A2(n_1133),
.B1(n_879),
.B2(n_1126),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1379),
.Y(n_1484)
);

AO22x2_ASAP7_75t_L g1485 ( 
.A1(n_1461),
.A2(n_1384),
.B1(n_1402),
.B2(n_1395),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1365),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1379),
.B(n_1393),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1393),
.B(n_1396),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1428),
.A2(n_1145),
.B1(n_1172),
.B2(n_1165),
.Y(n_1489)
);

AO22x2_ASAP7_75t_L g1490 ( 
.A1(n_1444),
.A2(n_1340),
.B1(n_1072),
.B2(n_1124),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1390),
.A2(n_1274),
.B1(n_1296),
.B2(n_1218),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1412),
.B(n_1013),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1415),
.A2(n_1356),
.B1(n_854),
.B2(n_858),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1462),
.A2(n_1353),
.B1(n_866),
.B2(n_907),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1396),
.B(n_1413),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_R g1496 ( 
.A1(n_1400),
.A2(n_1405),
.B1(n_1414),
.B2(n_1410),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1467),
.A2(n_1446),
.B1(n_1424),
.B2(n_1440),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1425),
.Y(n_1498)
);

OA22x2_ASAP7_75t_L g1499 ( 
.A1(n_1361),
.A2(n_1346),
.B1(n_1125),
.B2(n_856),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1360),
.A2(n_1022),
.B1(n_1183),
.B2(n_1075),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1413),
.B(n_1357),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1364),
.A2(n_863),
.B1(n_864),
.B2(n_861),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1420),
.B(n_1237),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1398),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1437),
.Y(n_1505)
);

OAI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1367),
.A2(n_873),
.B1(n_876),
.B2(n_870),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1453),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1420),
.B(n_1237),
.Y(n_1508)
);

AND2x2_ASAP7_75t_SL g1509 ( 
.A(n_1360),
.B(n_867),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1418),
.A2(n_880),
.B1(n_881),
.B2(n_878),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1372),
.A2(n_1216),
.B1(n_1287),
.B2(n_1264),
.Y(n_1511)
);

OA22x2_ASAP7_75t_L g1512 ( 
.A1(n_1447),
.A2(n_912),
.B1(n_921),
.B2(n_903),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1438),
.A2(n_1353),
.B1(n_866),
.B2(n_907),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1448),
.B(n_1255),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1448),
.B(n_1358),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1445),
.Y(n_1516)
);

XOR2xp5_ASAP7_75t_L g1517 ( 
.A(n_1372),
.B(n_862),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1434),
.A2(n_913),
.B1(n_952),
.B2(n_862),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1399),
.A2(n_1323),
.B1(n_1326),
.B2(n_1292),
.Y(n_1519)
);

AO22x2_ASAP7_75t_L g1520 ( 
.A1(n_1454),
.A2(n_1260),
.B1(n_1349),
.B2(n_1108),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1437),
.Y(n_1521)
);

NAND2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1454),
.B(n_913),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1455),
.A2(n_1332),
.B1(n_1355),
.B2(n_1005),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1455),
.A2(n_885),
.B1(n_892),
.B2(n_884),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1380),
.B(n_1351),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1442),
.A2(n_1000),
.B1(n_1001),
.B2(n_952),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1460),
.Y(n_1527)
);

AND2x2_ASAP7_75t_SL g1528 ( 
.A(n_1426),
.B(n_867),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1369),
.B(n_1255),
.Y(n_1529)
);

AO22x2_ASAP7_75t_L g1530 ( 
.A1(n_1392),
.A2(n_1359),
.B1(n_857),
.B2(n_859),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1362),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1466),
.A2(n_898),
.B1(n_900),
.B2(n_895),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1427),
.A2(n_906),
.B1(n_909),
.B2(n_905),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1369),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1431),
.A2(n_911),
.B1(n_914),
.B2(n_910),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1399),
.A2(n_916),
.B1(n_918),
.B2(n_915),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1371),
.B(n_1255),
.Y(n_1537)
);

OAI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1370),
.A2(n_926),
.B1(n_927),
.B2(n_923),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1371),
.B(n_1288),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1371),
.B(n_1288),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1370),
.B(n_1013),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1399),
.A2(n_930),
.B1(n_931),
.B2(n_929),
.Y(n_1542)
);

OAI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1373),
.A2(n_933),
.B1(n_934),
.B2(n_932),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1373),
.B(n_1288),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1466),
.A2(n_936),
.B1(n_937),
.B2(n_935),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1381),
.B(n_947),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1466),
.A2(n_941),
.B1(n_942),
.B2(n_938),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1381),
.B(n_1331),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1443),
.A2(n_1001),
.B1(n_1034),
.B2(n_1000),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1465),
.B(n_1334),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1465),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1443),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1375),
.Y(n_1553)
);

AO22x2_ASAP7_75t_L g1554 ( 
.A1(n_1450),
.A2(n_860),
.B1(n_865),
.B2(n_853),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1450),
.B(n_1331),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1376),
.B(n_868),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1466),
.A2(n_944),
.B1(n_946),
.B2(n_943),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1388),
.A2(n_949),
.B1(n_950),
.B2(n_948),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1401),
.B(n_1350),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1421),
.A2(n_953),
.B1(n_955),
.B2(n_951),
.Y(n_1560)
);

AND2x2_ASAP7_75t_SL g1561 ( 
.A(n_1399),
.B(n_947),
.Y(n_1561)
);

AO22x2_ASAP7_75t_L g1562 ( 
.A1(n_1422),
.A2(n_1341),
.B1(n_1343),
.B2(n_1338),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1435),
.A2(n_959),
.B1(n_962),
.B2(n_956),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1451),
.A2(n_969),
.B1(n_970),
.B2(n_966),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1458),
.A2(n_1111),
.B1(n_1118),
.B2(n_1034),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1435),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1435),
.B(n_1331),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1435),
.A2(n_978),
.B1(n_979),
.B2(n_974),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1374),
.Y(n_1569)
);

AO22x2_ASAP7_75t_L g1570 ( 
.A1(n_1374),
.A2(n_877),
.B1(n_882),
.B2(n_871),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1374),
.B(n_1348),
.Y(n_1571)
);

CKINVDCx6p67_ASAP7_75t_R g1572 ( 
.A(n_1389),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1389),
.Y(n_1573)
);

AO22x2_ASAP7_75t_L g1574 ( 
.A1(n_1389),
.A2(n_1345),
.B1(n_1352),
.B2(n_1328),
.Y(n_1574)
);

BUFx10_ASAP7_75t_L g1575 ( 
.A(n_1362),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1362),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1406),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1406),
.A2(n_985),
.B1(n_986),
.B2(n_982),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1377),
.B(n_883),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1377),
.B(n_972),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1406),
.Y(n_1581)
);

OAI22xp33_ASAP7_75t_R g1582 ( 
.A1(n_1407),
.A2(n_890),
.B1(n_891),
.B2(n_886),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1407),
.A2(n_992),
.B1(n_993),
.B2(n_990),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1407),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1408),
.A2(n_998),
.B1(n_999),
.B2(n_996),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1408),
.B(n_1348),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1408),
.A2(n_1004),
.B1(n_1006),
.B2(n_1003),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1433),
.B(n_1348),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1377),
.B(n_893),
.Y(n_1589)
);

AND2x2_ASAP7_75t_SL g1590 ( 
.A(n_1391),
.B(n_972),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1433),
.Y(n_1591)
);

AO22x2_ASAP7_75t_L g1592 ( 
.A1(n_1433),
.A2(n_897),
.B1(n_908),
.B2(n_896),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1452),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1452),
.Y(n_1594)
);

OR2x6_ASAP7_75t_L g1595 ( 
.A(n_1391),
.B(n_1046),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1452),
.B(n_1354),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1391),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1394),
.A2(n_1008),
.B1(n_1010),
.B2(n_1007),
.Y(n_1598)
);

OAI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1394),
.A2(n_1118),
.B1(n_1121),
.B2(n_1111),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1394),
.B(n_1290),
.Y(n_1600)
);

INVx8_ASAP7_75t_L g1601 ( 
.A(n_1403),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1403),
.A2(n_1019),
.B1(n_1020),
.B2(n_1012),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1403),
.A2(n_1025),
.B1(n_1026),
.B2(n_1021),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1404),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_R g1605 ( 
.A1(n_1404),
.A2(n_920),
.B1(n_922),
.B2(n_919),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1404),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1409),
.B(n_1354),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1409),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1409),
.A2(n_1147),
.B1(n_1152),
.B2(n_1121),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1417),
.A2(n_1030),
.B1(n_1031),
.B2(n_1029),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1417),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1417),
.A2(n_1033),
.B1(n_1035),
.B2(n_1032),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1423),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1423),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1423),
.B(n_1354),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1429),
.B(n_1199),
.Y(n_1616)
);

OR2x6_ASAP7_75t_L g1617 ( 
.A(n_1429),
.B(n_1290),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1429),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1430),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1430),
.A2(n_1039),
.B1(n_1041),
.B2(n_1036),
.Y(n_1620)
);

AO22x2_ASAP7_75t_L g1621 ( 
.A1(n_1430),
.A2(n_954),
.B1(n_957),
.B2(n_940),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1432),
.B(n_1199),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1432),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1432),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1439),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1439),
.A2(n_1044),
.B1(n_1045),
.B2(n_1042),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1439),
.B(n_1236),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1449),
.B(n_1236),
.Y(n_1628)
);

AO22x2_ASAP7_75t_L g1629 ( 
.A1(n_1449),
.A2(n_964),
.B1(n_965),
.B2(n_963),
.Y(n_1629)
);

AO22x2_ASAP7_75t_L g1630 ( 
.A1(n_1449),
.A2(n_971),
.B1(n_981),
.B2(n_968),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1456),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1456),
.A2(n_1050),
.B1(n_1051),
.B2(n_1048),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1456),
.B(n_1258),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1457),
.Y(n_1634)
);

AOI22x1_ASAP7_75t_SL g1635 ( 
.A1(n_1457),
.A2(n_1152),
.B1(n_1161),
.B2(n_1147),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1457),
.B(n_983),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1459),
.A2(n_1189),
.B1(n_1205),
.B2(n_1161),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1459),
.B(n_1258),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1459),
.B(n_1155),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1463),
.A2(n_1056),
.B1(n_1057),
.B2(n_1055),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1463),
.B(n_1300),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1463),
.A2(n_1064),
.B1(n_1067),
.B2(n_1061),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1464),
.A2(n_1319),
.B1(n_1205),
.B2(n_1208),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1464),
.A2(n_1208),
.B1(n_1215),
.B2(n_1189),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1464),
.A2(n_1231),
.B1(n_1241),
.B2(n_1215),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1416),
.A2(n_1241),
.B1(n_1259),
.B2(n_1231),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1383),
.Y(n_1647)
);

AO22x2_ASAP7_75t_L g1648 ( 
.A1(n_1461),
.A2(n_988),
.B1(n_991),
.B2(n_989),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1382),
.B(n_1300),
.Y(n_1649)
);

AND2x2_ASAP7_75t_SL g1650 ( 
.A(n_1397),
.B(n_976),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1416),
.A2(n_1279),
.B1(n_1318),
.B2(n_1259),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_SL g1652 ( 
.A(n_1399),
.B(n_1069),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1416),
.A2(n_1073),
.B1(n_1076),
.B2(n_1071),
.Y(n_1653)
);

NAND3x1_ASAP7_75t_L g1654 ( 
.A(n_1461),
.B(n_1318),
.C(n_1279),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1363),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1385),
.B(n_995),
.Y(n_1656)
);

OAI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1416),
.A2(n_1319),
.B1(n_1002),
.B2(n_1016),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1382),
.B(n_1316),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1382),
.B(n_1316),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1416),
.A2(n_1017),
.B1(n_1024),
.B2(n_1015),
.Y(n_1660)
);

AO22x2_ASAP7_75t_L g1661 ( 
.A1(n_1461),
.A2(n_1028),
.B1(n_1037),
.B2(n_1027),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1363),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1386),
.A2(n_1082),
.B1(n_1083),
.B2(n_1077),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1382),
.B(n_1155),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1382),
.B(n_1322),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1386),
.A2(n_1085),
.B1(n_1086),
.B2(n_1084),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1382),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1386),
.A2(n_1089),
.B1(n_1090),
.B2(n_1087),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1363),
.Y(n_1669)
);

OAI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1416),
.A2(n_1094),
.B1(n_1097),
.B2(n_1092),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1473),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1484),
.B(n_1098),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1552),
.A2(n_1014),
.B(n_976),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1498),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1665),
.B(n_1100),
.Y(n_1675)
);

XNOR2xp5_ASAP7_75t_L g1676 ( 
.A(n_1517),
.B(n_1101),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_SL g1677 ( 
.A(n_1566),
.B(n_1104),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1522),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1468),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1505),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1544),
.B(n_1040),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1476),
.B(n_1106),
.Y(n_1682)
);

INVxp67_ASAP7_75t_SL g1683 ( 
.A(n_1652),
.Y(n_1683)
);

XOR2xp5_ASAP7_75t_L g1684 ( 
.A(n_1472),
.B(n_1325),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1475),
.B(n_1114),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_R g1686 ( 
.A(n_1492),
.B(n_1115),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1561),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1616),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1622),
.Y(n_1689)
);

INVx4_ASAP7_75t_SL g1690 ( 
.A(n_1469),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1580),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1521),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1647),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1621),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1562),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1562),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_SL g1697 ( 
.A(n_1492),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1667),
.B(n_1477),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1487),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1628),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1488),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1548),
.B(n_1049),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1555),
.A2(n_1046),
.B(n_1014),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1495),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_1516),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1579),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1567),
.B(n_1047),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1541),
.B(n_1047),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1589),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1471),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1483),
.B(n_1333),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1501),
.B(n_1116),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1636),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1621),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1503),
.B(n_1052),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1633),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1534),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1637),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1607),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1515),
.B(n_1120),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1615),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1529),
.Y(n_1722)
);

INVxp33_ASAP7_75t_L g1723 ( 
.A(n_1565),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1520),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1664),
.B(n_1158),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1469),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1629),
.Y(n_1727)
);

XOR2xp5_ASAP7_75t_L g1728 ( 
.A(n_1635),
.B(n_1339),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1530),
.Y(n_1729)
);

XOR2xp5_ASAP7_75t_L g1730 ( 
.A(n_1646),
.B(n_1342),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1530),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1554),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1554),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1650),
.B(n_1485),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1629),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1630),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1479),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1630),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1556),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1485),
.B(n_1122),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1481),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1486),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1656),
.B(n_1127),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1504),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1507),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1638),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1527),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1655),
.Y(n_1748)
);

NAND2xp33_ASAP7_75t_R g1749 ( 
.A(n_1541),
.B(n_1128),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1662),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1519),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1489),
.B(n_1130),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1669),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1508),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1649),
.B(n_1136),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1479),
.B(n_1648),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1514),
.B(n_1137),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1571),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1658),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1586),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1509),
.B(n_1158),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1659),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1588),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1553),
.A2(n_1149),
.B(n_1062),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1596),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1537),
.Y(n_1766)
);

AND2x6_ASAP7_75t_L g1767 ( 
.A(n_1532),
.B(n_1344),
.Y(n_1767)
);

INVx3_ASAP7_75t_R g1768 ( 
.A(n_1525),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1539),
.Y(n_1769)
);

XNOR2x2_ASAP7_75t_L g1770 ( 
.A(n_1520),
.B(n_1053),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1559),
.A2(n_1149),
.B(n_1062),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1540),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1546),
.Y(n_1773)
);

OR2x6_ASAP7_75t_L g1774 ( 
.A(n_1648),
.B(n_1177),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1546),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1500),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_1663),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1590),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1511),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1523),
.B(n_1058),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1666),
.B(n_1139),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1661),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1661),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1528),
.B(n_1140),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1627),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1494),
.B(n_1148),
.C(n_1143),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1641),
.Y(n_1787)
);

INVxp33_ASAP7_75t_L g1788 ( 
.A(n_1668),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1512),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1572),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1580),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1595),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1536),
.B(n_1158),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1595),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1600),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1600),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1524),
.B(n_1150),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1499),
.B(n_1151),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1617),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1617),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1497),
.B(n_1153),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1542),
.B(n_1344),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1570),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1545),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1570),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1578),
.B(n_1154),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1574),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1547),
.B(n_1158),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1490),
.B(n_1156),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1657),
.B(n_1480),
.Y(n_1810)
);

CKINVDCx14_ASAP7_75t_R g1811 ( 
.A(n_1583),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1569),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_1557),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1574),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1592),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1592),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1550),
.Y(n_1817)
);

NOR2xp67_ASAP7_75t_L g1818 ( 
.A(n_1602),
.B(n_13),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1605),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1490),
.B(n_1159),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1598),
.Y(n_1821)
);

XNOR2xp5_ASAP7_75t_L g1822 ( 
.A(n_1654),
.B(n_1160),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1585),
.B(n_1162),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1612),
.Y(n_1824)
);

AND2x6_ASAP7_75t_L g1825 ( 
.A(n_1563),
.B(n_1344),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1551),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1603),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1518),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1610),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1620),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1626),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1632),
.Y(n_1832)
);

NAND2xp33_ASAP7_75t_R g1833 ( 
.A(n_1496),
.B(n_1164),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1640),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1642),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1587),
.B(n_1168),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1584),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1591),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1470),
.B(n_1171),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1526),
.B(n_1174),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1573),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1533),
.B(n_1175),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1593),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1568),
.Y(n_1844)
);

OR2x6_ASAP7_75t_L g1845 ( 
.A(n_1478),
.B(n_1177),
.Y(n_1845)
);

BUFx2_ASAP7_75t_SL g1846 ( 
.A(n_1581),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_1651),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1535),
.B(n_1558),
.Y(n_1848)
);

OR2x6_ASAP7_75t_L g1849 ( 
.A(n_1582),
.B(n_1198),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1482),
.Y(n_1850)
);

XOR2xp5_ASAP7_75t_L g1851 ( 
.A(n_1513),
.B(n_1330),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1560),
.B(n_1176),
.Y(n_1852)
);

XNOR2x2_ASAP7_75t_L g1853 ( 
.A(n_1599),
.B(n_1060),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1491),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1549),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1564),
.Y(n_1856)
);

XOR2x2_ASAP7_75t_L g1857 ( 
.A(n_1474),
.B(n_13),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1543),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1594),
.Y(n_1859)
);

XOR2xp5_ASAP7_75t_L g1860 ( 
.A(n_1609),
.B(n_1179),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1538),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1577),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1601),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1493),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1502),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1660),
.B(n_1158),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1643),
.B(n_1180),
.Y(n_1867)
);

AND2x2_ASAP7_75t_SL g1868 ( 
.A(n_1644),
.B(n_1198),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1575),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1506),
.B(n_1158),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1510),
.B(n_1187),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1639),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1653),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1645),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1670),
.B(n_1188),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1623),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1601),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1625),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1606),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1608),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1531),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1613),
.B(n_1314),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1619),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1631),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_1531),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1597),
.B(n_1190),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1576),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1634),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1576),
.Y(n_1889)
);

XOR2xp5_ASAP7_75t_L g1890 ( 
.A(n_1604),
.B(n_1327),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1611),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1614),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1618),
.B(n_1191),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1624),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1473),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_SL g1896 ( 
.A(n_1566),
.B(n_1192),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1473),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1468),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1484),
.B(n_1195),
.Y(n_1899)
);

XOR2x2_ASAP7_75t_L g1900 ( 
.A(n_1654),
.B(n_14),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1473),
.Y(n_1901)
);

XOR2xp5_ASAP7_75t_L g1902 ( 
.A(n_1517),
.B(n_1329),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1476),
.B(n_1196),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1544),
.B(n_1158),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1473),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_SL g1906 ( 
.A(n_1566),
.B(n_1197),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1616),
.Y(n_1907)
);

XNOR2x2_ASAP7_75t_L g1908 ( 
.A(n_1520),
.B(n_1063),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1476),
.B(n_1200),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1552),
.A2(n_1267),
.B(n_1263),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1484),
.B(n_1202),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1476),
.B(n_1203),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1476),
.B(n_1206),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1484),
.B(n_1207),
.Y(n_1914)
);

XOR2x2_ASAP7_75t_L g1915 ( 
.A(n_1654),
.B(n_14),
.Y(n_1915)
);

XOR2xp5_ASAP7_75t_L g1916 ( 
.A(n_1517),
.B(n_1310),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1473),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1473),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1476),
.B(n_1209),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1473),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1616),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1473),
.A2(n_1267),
.B(n_1263),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1473),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1616),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1616),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1473),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1473),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1566),
.B(n_1335),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_SL g1929 ( 
.A(n_1492),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1473),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1476),
.B(n_1210),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1516),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1484),
.B(n_1211),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1473),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1473),
.Y(n_1935)
);

XNOR2xp5_ASAP7_75t_L g1936 ( 
.A(n_1517),
.B(n_1220),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1476),
.B(n_1224),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1473),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1468),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1473),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1476),
.B(n_1225),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1517),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1484),
.B(n_1227),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1473),
.Y(n_1944)
);

BUFx8_ASAP7_75t_L g1945 ( 
.A(n_1476),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1473),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1473),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1476),
.B(n_1229),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1473),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1566),
.Y(n_1950)
);

XOR2xp5_ASAP7_75t_L g1951 ( 
.A(n_1517),
.B(n_1304),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1468),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1484),
.B(n_1233),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1484),
.B(n_1235),
.Y(n_1954)
);

XOR2xp5_ASAP7_75t_L g1955 ( 
.A(n_1517),
.B(n_1307),
.Y(n_1955)
);

XOR2xp5_ASAP7_75t_L g1956 ( 
.A(n_1517),
.B(n_1308),
.Y(n_1956)
);

INVx4_ASAP7_75t_L g1957 ( 
.A(n_1566),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1473),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1743),
.B(n_1238),
.Y(n_1959)
);

INVx1_ASAP7_75t_SL g1960 ( 
.A(n_1932),
.Y(n_1960)
);

AND2x6_ASAP7_75t_L g1961 ( 
.A(n_1735),
.B(n_1736),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1671),
.B(n_1240),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1694),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1671),
.B(n_1674),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1674),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1870),
.A2(n_1066),
.B(n_1065),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1680),
.B(n_1245),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1680),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1685),
.B(n_1252),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1840),
.B(n_1254),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1837),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1705),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1938),
.B(n_1256),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1838),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1828),
.B(n_1698),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1697),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1690),
.B(n_1773),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1774),
.B(n_1257),
.Y(n_1978)
);

BUFx2_ASAP7_75t_L g1979 ( 
.A(n_1774),
.Y(n_1979)
);

INVx3_ASAP7_75t_SL g1980 ( 
.A(n_1690),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1863),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1950),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1881),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1756),
.B(n_1265),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1950),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1756),
.B(n_1266),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1775),
.B(n_1068),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1681),
.B(n_1070),
.Y(n_1988)
);

NAND2x1p5_ASAP7_75t_L g1989 ( 
.A(n_1691),
.B(n_1270),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1843),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1691),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1885),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1938),
.B(n_1268),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1810),
.B(n_1269),
.Y(n_1994)
);

AND2x2_ASAP7_75t_SL g1995 ( 
.A(n_1724),
.B(n_1344),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1940),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1940),
.B(n_1271),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1682),
.B(n_1272),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1944),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1903),
.B(n_1273),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1944),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1946),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1812),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1863),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1714),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1681),
.B(n_1078),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1909),
.B(n_1276),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1946),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1793),
.A2(n_1088),
.B(n_1081),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1841),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1727),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1947),
.B(n_1277),
.Y(n_2012)
);

AND2x2_ASAP7_75t_SL g2013 ( 
.A(n_1738),
.B(n_1270),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1912),
.B(n_1278),
.Y(n_2014)
);

NAND2x1p5_ASAP7_75t_L g2015 ( 
.A(n_1691),
.B(n_1309),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1695),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1863),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1947),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1949),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1913),
.B(n_1282),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1896),
.B(n_1283),
.Y(n_2021)
);

AND2x2_ASAP7_75t_SL g2022 ( 
.A(n_1868),
.B(n_1309),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1919),
.B(n_1285),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1859),
.Y(n_2024)
);

NOR2xp67_ASAP7_75t_L g2025 ( 
.A(n_1726),
.B(n_15),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1949),
.B(n_1291),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1808),
.A2(n_1093),
.B(n_1091),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1679),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1957),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1816),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1958),
.B(n_1294),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1697),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1958),
.B(n_1295),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1717),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1692),
.B(n_1297),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1679),
.Y(n_2036)
);

AND2x2_ASAP7_75t_SL g2037 ( 
.A(n_1707),
.B(n_1074),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1741),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1931),
.B(n_1298),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1742),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1957),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1950),
.Y(n_2042)
);

NAND2x1p5_ASAP7_75t_L g2043 ( 
.A(n_1729),
.B(n_1095),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1768),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1722),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1906),
.B(n_1299),
.Y(n_2046)
);

INVxp67_ASAP7_75t_SL g2047 ( 
.A(n_1696),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1739),
.Y(n_2048)
);

INVx3_ASAP7_75t_L g2049 ( 
.A(n_1687),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1937),
.B(n_1941),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1693),
.B(n_1306),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_1687),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1687),
.B(n_1311),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1948),
.B(n_1336),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_1702),
.B(n_1096),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1699),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1895),
.B(n_1897),
.Y(n_2057)
);

AND2x2_ASAP7_75t_SL g2058 ( 
.A(n_1732),
.B(n_1079),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1702),
.B(n_1337),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1701),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1740),
.B(n_1102),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1744),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1901),
.B(n_1103),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1704),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1867),
.B(n_1105),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1745),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1905),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1711),
.B(n_1107),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1754),
.B(n_1109),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1790),
.Y(n_2070)
);

AND2x4_ASAP7_75t_L g2071 ( 
.A(n_1710),
.B(n_1110),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1855),
.B(n_1112),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1755),
.B(n_1113),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1752),
.B(n_1819),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1734),
.B(n_1117),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1839),
.B(n_1119),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1688),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1747),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1781),
.B(n_1131),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1898),
.B(n_1134),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1730),
.B(n_1135),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1759),
.B(n_1146),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1917),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1703),
.A2(n_1166),
.B(n_1163),
.Y(n_2084)
);

INVx4_ASAP7_75t_L g2085 ( 
.A(n_1708),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1748),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1939),
.B(n_1167),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_1860),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_1952),
.B(n_1169),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1689),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1700),
.Y(n_2091)
);

AND2x2_ASAP7_75t_SL g2092 ( 
.A(n_1786),
.B(n_1173),
.Y(n_2092)
);

INVxp67_ASAP7_75t_SL g2093 ( 
.A(n_1733),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1762),
.B(n_1178),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1809),
.B(n_1184),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1918),
.Y(n_2096)
);

AND2x2_ASAP7_75t_SL g2097 ( 
.A(n_1874),
.B(n_1193),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1820),
.B(n_1194),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1920),
.B(n_1212),
.Y(n_2099)
);

INVx3_ASAP7_75t_L g2100 ( 
.A(n_1716),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1923),
.B(n_1213),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1926),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1776),
.B(n_1214),
.Y(n_2103)
);

INVx2_ASAP7_75t_SL g2104 ( 
.A(n_1945),
.Y(n_2104)
);

CKINVDCx12_ASAP7_75t_R g2105 ( 
.A(n_1708),
.Y(n_2105)
);

AND2x4_ASAP7_75t_SL g2106 ( 
.A(n_1942),
.B(n_1219),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1715),
.B(n_1719),
.Y(n_2107)
);

AND2x2_ASAP7_75t_SL g2108 ( 
.A(n_1731),
.B(n_1079),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1683),
.B(n_1079),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1927),
.B(n_1222),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_1945),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1930),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1887),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1934),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1746),
.Y(n_2115)
);

BUFx3_ASAP7_75t_L g2116 ( 
.A(n_1737),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1803),
.B(n_1079),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1935),
.Y(n_2118)
);

AND2x2_ASAP7_75t_SL g2119 ( 
.A(n_1782),
.B(n_1783),
.Y(n_2119)
);

INVx1_ASAP7_75t_SL g2120 ( 
.A(n_1846),
.Y(n_2120)
);

INVx4_ASAP7_75t_L g2121 ( 
.A(n_1929),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1817),
.B(n_1779),
.Y(n_2122)
);

INVxp67_ASAP7_75t_SL g2123 ( 
.A(n_1751),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1750),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1780),
.B(n_1223),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1721),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1827),
.B(n_1230),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1780),
.B(n_1232),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1753),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1907),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1706),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1715),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1829),
.B(n_1234),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1826),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1921),
.Y(n_2135)
);

AND2x2_ASAP7_75t_SL g2136 ( 
.A(n_1678),
.B(n_1239),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_1924),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_1805),
.Y(n_2138)
);

INVx4_ASAP7_75t_L g2139 ( 
.A(n_1929),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1830),
.B(n_1242),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1833),
.A2(n_1244),
.B1(n_1246),
.B2(n_1243),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_1869),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1784),
.B(n_1248),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1925),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1836),
.B(n_1250),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1758),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1760),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_1882),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1763),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1877),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1718),
.B(n_1261),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_1684),
.B(n_1262),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_1831),
.B(n_1275),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1832),
.B(n_1280),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1709),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1807),
.Y(n_2156)
);

BUFx3_ASAP7_75t_L g2157 ( 
.A(n_1785),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1788),
.B(n_1281),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_1791),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_1814),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1765),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_SL g2162 ( 
.A(n_1815),
.B(n_1286),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1713),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1849),
.B(n_1302),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1766),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1769),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1849),
.B(n_1305),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1845),
.B(n_1312),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1845),
.B(n_1313),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_1902),
.B(n_1317),
.Y(n_2170)
);

AND2x4_ASAP7_75t_SL g2171 ( 
.A(n_1847),
.B(n_1321),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1834),
.B(n_15),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1835),
.B(n_15),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1771),
.B(n_16),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1922),
.B(n_1844),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1851),
.B(n_16),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1866),
.B(n_17),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1677),
.B(n_1204),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1856),
.B(n_1204),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1767),
.Y(n_2180)
);

BUFx3_ASAP7_75t_L g2181 ( 
.A(n_1787),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1801),
.B(n_17),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1797),
.B(n_17),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1904),
.B(n_18),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1798),
.B(n_18),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_1862),
.Y(n_2186)
);

INVx2_ASAP7_75t_SL g2187 ( 
.A(n_1792),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1757),
.B(n_18),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1673),
.B(n_19),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1767),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1772),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1910),
.B(n_19),
.Y(n_2192)
);

NAND2x1p5_ASAP7_75t_L g2193 ( 
.A(n_1794),
.B(n_1204),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1850),
.B(n_19),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1886),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_1795),
.Y(n_2196)
);

BUFx3_ASAP7_75t_L g2197 ( 
.A(n_1821),
.Y(n_2197)
);

OAI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_1725),
.A2(n_1226),
.B(n_1204),
.Y(n_2198)
);

INVx4_ASAP7_75t_L g2199 ( 
.A(n_1767),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1854),
.B(n_20),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1858),
.B(n_20),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1864),
.B(n_20),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1878),
.Y(n_2203)
);

INVx3_ASAP7_75t_SL g2204 ( 
.A(n_1900),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_1818),
.Y(n_2205)
);

BUFx3_ASAP7_75t_L g2206 ( 
.A(n_1824),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1893),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_1796),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1761),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_1789),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1767),
.Y(n_2211)
);

INVx4_ASAP7_75t_L g2212 ( 
.A(n_1825),
.Y(n_2212)
);

BUFx3_ASAP7_75t_L g2213 ( 
.A(n_1861),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_1799),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1723),
.B(n_21),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1800),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1764),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1872),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_1770),
.Y(n_2219)
);

BUFx6f_ASAP7_75t_L g2220 ( 
.A(n_1825),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_1675),
.B(n_21),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1873),
.Y(n_2222)
);

AND2x2_ASAP7_75t_SL g2223 ( 
.A(n_1848),
.B(n_1908),
.Y(n_2223)
);

INVx4_ASAP7_75t_L g2224 ( 
.A(n_1825),
.Y(n_2224)
);

INVxp67_ASAP7_75t_L g2225 ( 
.A(n_1890),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1875),
.B(n_21),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1802),
.B(n_1825),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1712),
.B(n_1720),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1956),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1822),
.B(n_1806),
.Y(n_2230)
);

AND2x2_ASAP7_75t_SL g2231 ( 
.A(n_1916),
.B(n_1226),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1880),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1876),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_1823),
.B(n_22),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1853),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1842),
.B(n_22),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1852),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_1676),
.B(n_22),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1928),
.B(n_1226),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_1951),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1871),
.B(n_23),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_R g2242 ( 
.A(n_1749),
.B(n_23),
.Y(n_2242)
);

INVx4_ASAP7_75t_L g2243 ( 
.A(n_1865),
.Y(n_2243)
);

INVx4_ASAP7_75t_L g2244 ( 
.A(n_1889),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1778),
.B(n_1672),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1915),
.Y(n_2246)
);

AND2x2_ASAP7_75t_SL g2247 ( 
.A(n_1955),
.B(n_1226),
.Y(n_2247)
);

AND2x6_ASAP7_75t_L g2248 ( 
.A(n_1899),
.B(n_1293),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1936),
.B(n_23),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_1911),
.B(n_1293),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1811),
.B(n_24),
.Y(n_2251)
);

INVx1_ASAP7_75t_SL g2252 ( 
.A(n_1728),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_1889),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1914),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_1686),
.Y(n_2255)
);

AND2x2_ASAP7_75t_SL g2256 ( 
.A(n_1777),
.B(n_1933),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1883),
.Y(n_2257)
);

AND2x2_ASAP7_75t_SL g2258 ( 
.A(n_1943),
.B(n_1293),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_1953),
.B(n_1293),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1954),
.Y(n_2260)
);

AND2x6_ASAP7_75t_L g2261 ( 
.A(n_1884),
.B(n_1320),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1804),
.B(n_24),
.Y(n_2262)
);

BUFx3_ASAP7_75t_L g2263 ( 
.A(n_1813),
.Y(n_2263)
);

OAI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_1888),
.A2(n_1320),
.B(n_25),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1879),
.B(n_1320),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1857),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1891),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_1892),
.B(n_25),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1894),
.B(n_1320),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1671),
.B(n_25),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_1690),
.B(n_26),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_1743),
.B(n_26),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1837),
.Y(n_2273)
);

HB1xp67_ASAP7_75t_L g2274 ( 
.A(n_1694),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1671),
.B(n_26),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1837),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1671),
.Y(n_2277)
);

NOR2xp67_ASAP7_75t_SL g2278 ( 
.A(n_1950),
.B(n_28),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_1743),
.B(n_27),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1837),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1743),
.B(n_27),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1671),
.B(n_27),
.Y(n_2282)
);

AND2x2_ASAP7_75t_SL g2283 ( 
.A(n_1868),
.B(n_28),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1743),
.B(n_29),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1837),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1694),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_1681),
.B(n_29),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1671),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_1694),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1743),
.B(n_30),
.Y(n_2290)
);

INVx4_ASAP7_75t_L g2291 ( 
.A(n_1863),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1671),
.B(n_31),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1671),
.B(n_31),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1837),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1837),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1743),
.B(n_31),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1950),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1950),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1837),
.Y(n_2299)
);

OR2x2_ASAP7_75t_SL g2300 ( 
.A(n_1810),
.B(n_32),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_1743),
.B(n_32),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_1690),
.B(n_32),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1837),
.Y(n_2303)
);

NAND2x1p5_ASAP7_75t_L g2304 ( 
.A(n_1691),
.B(n_33),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1837),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_1681),
.B(n_33),
.Y(n_2306)
);

INVx2_ASAP7_75t_SL g2307 ( 
.A(n_1960),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_1982),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_1994),
.B(n_34),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1964),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2291),
.Y(n_2311)
);

INVx4_ASAP7_75t_L g2312 ( 
.A(n_1980),
.Y(n_2312)
);

AND2x2_ASAP7_75t_SL g2313 ( 
.A(n_1995),
.B(n_34),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1964),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1965),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2048),
.B(n_34),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1968),
.Y(n_2317)
);

OR2x6_ASAP7_75t_L g2318 ( 
.A(n_2104),
.B(n_35),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_SL g2319 ( 
.A(n_1995),
.B(n_35),
.Y(n_2319)
);

OR2x6_ASAP7_75t_L g2320 ( 
.A(n_2121),
.B(n_35),
.Y(n_2320)
);

BUFx4f_ASAP7_75t_L g2321 ( 
.A(n_1980),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2122),
.B(n_36),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2048),
.B(n_36),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1960),
.B(n_38),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_2120),
.Y(n_2325)
);

BUFx4f_ASAP7_75t_L g2326 ( 
.A(n_2271),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2122),
.B(n_37),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_1982),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2120),
.B(n_37),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1975),
.B(n_37),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2068),
.B(n_38),
.Y(n_2331)
);

BUFx2_ASAP7_75t_L g2332 ( 
.A(n_1972),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1996),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_1982),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2131),
.B(n_39),
.Y(n_2335)
);

BUFx3_ASAP7_75t_L g2336 ( 
.A(n_1983),
.Y(n_2336)
);

BUFx4f_ASAP7_75t_L g2337 ( 
.A(n_2271),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2155),
.B(n_39),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_1985),
.Y(n_2339)
);

OR2x6_ASAP7_75t_L g2340 ( 
.A(n_2121),
.B(n_2139),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_1992),
.Y(n_2341)
);

OR2x2_ASAP7_75t_L g2342 ( 
.A(n_2088),
.B(n_2240),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2163),
.B(n_40),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2075),
.B(n_40),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2213),
.B(n_41),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_2139),
.B(n_41),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2061),
.B(n_41),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1999),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2097),
.B(n_43),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_2088),
.B(n_43),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2001),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2002),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2148),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2008),
.Y(n_2354)
);

AO21x2_ASAP7_75t_L g2355 ( 
.A1(n_2198),
.A2(n_44),
.B(n_45),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2198),
.A2(n_66),
.B(n_64),
.Y(n_2356)
);

INVx2_ASAP7_75t_SL g2357 ( 
.A(n_2113),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2291),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2074),
.B(n_44),
.Y(n_2359)
);

INVx2_ASAP7_75t_SL g2360 ( 
.A(n_2111),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_1985),
.Y(n_2361)
);

AND2x6_ASAP7_75t_L g2362 ( 
.A(n_2180),
.B(n_44),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2148),
.B(n_45),
.Y(n_2363)
);

BUFx4f_ASAP7_75t_L g2364 ( 
.A(n_2302),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2029),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_SL g2366 ( 
.A(n_2058),
.B(n_46),
.Y(n_2366)
);

AND2x6_ASAP7_75t_L g2367 ( 
.A(n_2180),
.B(n_46),
.Y(n_2367)
);

AND2x2_ASAP7_75t_SL g2368 ( 
.A(n_2037),
.B(n_2283),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2050),
.B(n_46),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2065),
.B(n_47),
.Y(n_2370)
);

NAND2x1p5_ASAP7_75t_L g2371 ( 
.A(n_1991),
.B(n_47),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_1979),
.B(n_48),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2222),
.B(n_2076),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2057),
.B(n_49),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2018),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2019),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2057),
.B(n_49),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2277),
.Y(n_2378)
);

NAND2xp33_ASAP7_75t_L g2379 ( 
.A(n_2180),
.B(n_2190),
.Y(n_2379)
);

NAND2x1p5_ASAP7_75t_L g2380 ( 
.A(n_1991),
.B(n_49),
.Y(n_2380)
);

INVxp67_ASAP7_75t_L g2381 ( 
.A(n_2287),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2045),
.B(n_51),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_1970),
.B(n_51),
.Y(n_2383)
);

BUFx12f_ASAP7_75t_L g2384 ( 
.A(n_1976),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2067),
.B(n_51),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2083),
.B(n_52),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2197),
.B(n_52),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_1959),
.B(n_1969),
.Y(n_2388)
);

BUFx3_ASAP7_75t_L g2389 ( 
.A(n_2017),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2096),
.B(n_52),
.Y(n_2390)
);

INVxp67_ASAP7_75t_SL g2391 ( 
.A(n_2005),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_1985),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2032),
.Y(n_2393)
);

INVx2_ASAP7_75t_SL g2394 ( 
.A(n_2111),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2116),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2029),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2237),
.B(n_2132),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2206),
.B(n_53),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2288),
.Y(n_2399)
);

OR2x6_ASAP7_75t_L g2400 ( 
.A(n_2085),
.B(n_53),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2041),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2102),
.B(n_53),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2112),
.B(n_54),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2042),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2085),
.B(n_54),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_1998),
.B(n_54),
.Y(n_2406)
);

BUFx4f_ASAP7_75t_L g2407 ( 
.A(n_2302),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2114),
.B(n_55),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2256),
.B(n_55),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2228),
.B(n_56),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2118),
.B(n_56),
.Y(n_2411)
);

AND2x4_ASAP7_75t_L g2412 ( 
.A(n_2186),
.B(n_57),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2134),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_2042),
.Y(n_2414)
);

OR2x6_ASAP7_75t_L g2415 ( 
.A(n_2304),
.B(n_57),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2138),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2142),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_1977),
.B(n_57),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_SL g2419 ( 
.A(n_2231),
.B(n_58),
.Y(n_2419)
);

OR2x2_ASAP7_75t_L g2420 ( 
.A(n_2240),
.B(n_58),
.Y(n_2420)
);

INVxp67_ASAP7_75t_L g2421 ( 
.A(n_2287),
.Y(n_2421)
);

INVxp67_ASAP7_75t_L g2422 ( 
.A(n_2306),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2105),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_1971),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1974),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2138),
.Y(n_2426)
);

BUFx10_ASAP7_75t_L g2427 ( 
.A(n_1977),
.Y(n_2427)
);

BUFx6f_ASAP7_75t_L g2428 ( 
.A(n_2042),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_1990),
.Y(n_2429)
);

INVx2_ASAP7_75t_SL g2430 ( 
.A(n_2070),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2000),
.B(n_59),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2228),
.B(n_59),
.Y(n_2432)
);

NAND2x1p5_ASAP7_75t_L g2433 ( 
.A(n_2037),
.B(n_59),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_SL g2434 ( 
.A(n_2247),
.B(n_60),
.Y(n_2434)
);

BUFx12f_ASAP7_75t_L g2435 ( 
.A(n_2243),
.Y(n_2435)
);

OR2x2_ASAP7_75t_L g2436 ( 
.A(n_2081),
.B(n_60),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2072),
.B(n_60),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2056),
.B(n_61),
.Y(n_2438)
);

CKINVDCx20_ASAP7_75t_R g2439 ( 
.A(n_2242),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2095),
.B(n_61),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2007),
.B(n_62),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2160),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_2242),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2297),
.Y(n_2444)
);

NAND2x1p5_ASAP7_75t_L g2445 ( 
.A(n_1981),
.B(n_2004),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2098),
.B(n_63),
.Y(n_2446)
);

AND2x2_ASAP7_75t_SL g2447 ( 
.A(n_2058),
.B(n_63),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2044),
.Y(n_2448)
);

OR2x6_ASAP7_75t_L g2449 ( 
.A(n_2304),
.B(n_66),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2230),
.B(n_848),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_2041),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2153),
.B(n_67),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2160),
.Y(n_2453)
);

INVxp67_ASAP7_75t_L g2454 ( 
.A(n_2306),
.Y(n_2454)
);

NAND2x1p5_ASAP7_75t_L g2455 ( 
.A(n_1981),
.B(n_68),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2273),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2153),
.B(n_2158),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2016),
.Y(n_2458)
);

BUFx2_ASAP7_75t_SL g2459 ( 
.A(n_2044),
.Y(n_2459)
);

INVxp67_ASAP7_75t_L g2460 ( 
.A(n_2059),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_SL g2461 ( 
.A(n_2108),
.B(n_67),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2276),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2152),
.B(n_68),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2016),
.Y(n_2464)
);

INVx6_ASAP7_75t_L g2465 ( 
.A(n_2090),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2014),
.B(n_69),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2079),
.B(n_71),
.Y(n_2467)
);

AND2x2_ASAP7_75t_SL g2468 ( 
.A(n_2108),
.B(n_71),
.Y(n_2468)
);

INVx3_ASAP7_75t_L g2469 ( 
.A(n_2297),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2047),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2297),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_SL g2472 ( 
.A(n_2199),
.B(n_72),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2280),
.Y(n_2473)
);

AND2x4_ASAP7_75t_L g2474 ( 
.A(n_2060),
.B(n_72),
.Y(n_2474)
);

INVx5_ASAP7_75t_L g2475 ( 
.A(n_2298),
.Y(n_2475)
);

BUFx4f_ASAP7_75t_L g2476 ( 
.A(n_2194),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2020),
.B(n_2023),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2285),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2272),
.B(n_73),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2047),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2064),
.B(n_73),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2093),
.Y(n_2482)
);

BUFx2_ASAP7_75t_L g2483 ( 
.A(n_1989),
.Y(n_2483)
);

INVx3_ASAP7_75t_L g2484 ( 
.A(n_2298),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2262),
.B(n_74),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2279),
.B(n_74),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2294),
.Y(n_2487)
);

INVx3_ASAP7_75t_L g2488 ( 
.A(n_2298),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2233),
.B(n_75),
.Y(n_2489)
);

INVx2_ASAP7_75t_SL g2490 ( 
.A(n_2107),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2295),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_2052),
.Y(n_2492)
);

INVx6_ASAP7_75t_L g2493 ( 
.A(n_2090),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2093),
.Y(n_2494)
);

BUFx4f_ASAP7_75t_L g2495 ( 
.A(n_2194),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2004),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2299),
.Y(n_2497)
);

INVx5_ASAP7_75t_L g2498 ( 
.A(n_2052),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2270),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2039),
.B(n_76),
.Y(n_2500)
);

OR2x6_ASAP7_75t_L g2501 ( 
.A(n_2255),
.B(n_76),
.Y(n_2501)
);

INVx5_ASAP7_75t_L g2502 ( 
.A(n_2052),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2281),
.B(n_2284),
.Y(n_2503)
);

BUFx3_ASAP7_75t_L g2504 ( 
.A(n_2107),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2270),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2290),
.B(n_77),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2195),
.B(n_77),
.Y(n_2507)
);

OR2x6_ASAP7_75t_L g2508 ( 
.A(n_2255),
.B(n_78),
.Y(n_2508)
);

NAND2x1p5_ASAP7_75t_L g2509 ( 
.A(n_2028),
.B(n_80),
.Y(n_2509)
);

AND2x2_ASAP7_75t_SL g2510 ( 
.A(n_2022),
.B(n_79),
.Y(n_2510)
);

INVx4_ASAP7_75t_L g2511 ( 
.A(n_1989),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2275),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_2049),
.Y(n_2513)
);

INVx4_ASAP7_75t_L g2514 ( 
.A(n_2015),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2275),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2282),
.Y(n_2516)
);

BUFx12f_ASAP7_75t_L g2517 ( 
.A(n_2243),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2282),
.Y(n_2518)
);

NAND2x1_ASAP7_75t_SL g2519 ( 
.A(n_2204),
.B(n_1984),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2162),
.B(n_79),
.Y(n_2520)
);

OR2x2_ASAP7_75t_L g2521 ( 
.A(n_2262),
.B(n_81),
.Y(n_2521)
);

AND2x4_ASAP7_75t_L g2522 ( 
.A(n_2207),
.B(n_82),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2015),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2296),
.B(n_83),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2303),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2054),
.B(n_83),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2301),
.B(n_84),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2292),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2292),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2176),
.B(n_84),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2145),
.B(n_85),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_1978),
.B(n_2171),
.Y(n_2532)
);

INVxp67_ASAP7_75t_L g2533 ( 
.A(n_2059),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2136),
.B(n_849),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2049),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2183),
.B(n_85),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_SL g2537 ( 
.A(n_2199),
.B(n_86),
.Y(n_2537)
);

OR2x6_ASAP7_75t_L g2538 ( 
.A(n_2229),
.B(n_86),
.Y(n_2538)
);

OR2x2_ASAP7_75t_L g2539 ( 
.A(n_2170),
.B(n_87),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_2190),
.Y(n_2540)
);

BUFx2_ASAP7_75t_L g2541 ( 
.A(n_2005),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2234),
.B(n_87),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2106),
.Y(n_2543)
);

AOI21x1_ASAP7_75t_L g2544 ( 
.A1(n_2109),
.A2(n_88),
.B(n_89),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2146),
.B(n_88),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2143),
.B(n_89),
.Y(n_2546)
);

BUFx2_ASAP7_75t_L g2547 ( 
.A(n_2011),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2165),
.B(n_90),
.Y(n_2548)
);

OR2x6_ASAP7_75t_L g2549 ( 
.A(n_2229),
.B(n_91),
.Y(n_2549)
);

BUFx6f_ASAP7_75t_L g2550 ( 
.A(n_2190),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2147),
.B(n_92),
.Y(n_2551)
);

INVx3_ASAP7_75t_L g2552 ( 
.A(n_2090),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_L g2553 ( 
.A(n_2254),
.B(n_838),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2191),
.B(n_92),
.Y(n_2554)
);

CKINVDCx8_ASAP7_75t_R g2555 ( 
.A(n_1988),
.Y(n_2555)
);

AND2x4_ASAP7_75t_L g2556 ( 
.A(n_2149),
.B(n_93),
.Y(n_2556)
);

NOR2xp33_ASAP7_75t_L g2557 ( 
.A(n_2260),
.B(n_841),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2293),
.Y(n_2558)
);

BUFx6f_ASAP7_75t_L g2559 ( 
.A(n_2211),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2161),
.B(n_94),
.Y(n_2560)
);

INVx6_ASAP7_75t_L g2561 ( 
.A(n_2115),
.Y(n_2561)
);

INVx4_ASAP7_75t_L g2562 ( 
.A(n_2212),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2125),
.B(n_94),
.Y(n_2563)
);

BUFx2_ASAP7_75t_L g2564 ( 
.A(n_2011),
.Y(n_2564)
);

BUFx4f_ASAP7_75t_L g2565 ( 
.A(n_2119),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2128),
.B(n_95),
.Y(n_2566)
);

OR2x6_ASAP7_75t_L g2567 ( 
.A(n_2225),
.B(n_95),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2103),
.B(n_2126),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_L g2569 ( 
.A(n_2211),
.Y(n_2569)
);

HB1xp67_ASAP7_75t_L g2570 ( 
.A(n_2274),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2293),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2245),
.B(n_846),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2182),
.B(n_96),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2266),
.B(n_96),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2305),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_1988),
.B(n_2006),
.Y(n_2576)
);

CKINVDCx8_ASAP7_75t_R g2577 ( 
.A(n_2006),
.Y(n_2577)
);

OR2x6_ASAP7_75t_L g2578 ( 
.A(n_2225),
.B(n_97),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_2245),
.B(n_847),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2166),
.B(n_97),
.Y(n_2580)
);

NAND2x1p5_ASAP7_75t_L g2581 ( 
.A(n_2036),
.B(n_2150),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2175),
.Y(n_2582)
);

AND2x4_ASAP7_75t_L g2583 ( 
.A(n_2214),
.B(n_98),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2226),
.B(n_98),
.Y(n_2584)
);

AND2x6_ASAP7_75t_L g2585 ( 
.A(n_2211),
.B(n_99),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2172),
.B(n_99),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2172),
.B(n_100),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2175),
.Y(n_2588)
);

NOR2x1_ASAP7_75t_L g2589 ( 
.A(n_2212),
.B(n_101),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2173),
.B(n_101),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2156),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2115),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_L g2593 ( 
.A(n_2220),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2156),
.Y(n_2594)
);

BUFx6f_ASAP7_75t_SL g2595 ( 
.A(n_2263),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2156),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2214),
.B(n_102),
.Y(n_2597)
);

BUFx12f_ASAP7_75t_L g2598 ( 
.A(n_2300),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2203),
.Y(n_2599)
);

OR2x6_ASAP7_75t_L g2600 ( 
.A(n_2043),
.B(n_103),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2274),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2205),
.B(n_833),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2135),
.B(n_103),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2055),
.B(n_105),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2232),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2205),
.B(n_835),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2055),
.B(n_105),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_2035),
.B(n_837),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2038),
.Y(n_2609)
);

CKINVDCx20_ASAP7_75t_R g2610 ( 
.A(n_2204),
.Y(n_2610)
);

INVx6_ASAP7_75t_L g2611 ( 
.A(n_2115),
.Y(n_2611)
);

AND2x2_ASAP7_75t_SL g2612 ( 
.A(n_2022),
.B(n_106),
.Y(n_2612)
);

NOR2x1_ASAP7_75t_L g2613 ( 
.A(n_2224),
.B(n_107),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2286),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2173),
.B(n_107),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2257),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2040),
.Y(n_2617)
);

INVxp67_ASAP7_75t_SL g2618 ( 
.A(n_2286),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_1962),
.B(n_108),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2062),
.Y(n_2620)
);

OR2x6_ASAP7_75t_L g2621 ( 
.A(n_2043),
.B(n_108),
.Y(n_2621)
);

INVx4_ASAP7_75t_L g2622 ( 
.A(n_2224),
.Y(n_2622)
);

INVx3_ASAP7_75t_L g2623 ( 
.A(n_2244),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2030),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2030),
.Y(n_2625)
);

BUFx2_ASAP7_75t_L g2626 ( 
.A(n_2289),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2289),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_SL g2628 ( 
.A(n_2252),
.B(n_109),
.Y(n_2628)
);

AND2x4_ASAP7_75t_L g2629 ( 
.A(n_2144),
.B(n_110),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2066),
.Y(n_2630)
);

AND2x4_ASAP7_75t_L g2631 ( 
.A(n_2077),
.B(n_110),
.Y(n_2631)
);

BUFx2_ASAP7_75t_L g2632 ( 
.A(n_2071),
.Y(n_2632)
);

CKINVDCx8_ASAP7_75t_R g2633 ( 
.A(n_2071),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2034),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2220),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2078),
.Y(n_2636)
);

OR2x6_ASAP7_75t_L g2637 ( 
.A(n_2025),
.B(n_111),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2035),
.B(n_847),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2267),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_1962),
.B(n_112),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2051),
.B(n_849),
.Y(n_2641)
);

INVxp67_ASAP7_75t_L g2642 ( 
.A(n_2080),
.Y(n_2642)
);

BUFx4f_ASAP7_75t_L g2643 ( 
.A(n_2119),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2051),
.B(n_850),
.Y(n_2644)
);

NAND2x1p5_ASAP7_75t_L g2645 ( 
.A(n_2150),
.B(n_115),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2086),
.Y(n_2646)
);

BUFx3_ASAP7_75t_L g2647 ( 
.A(n_2077),
.Y(n_2647)
);

BUFx12f_ASAP7_75t_L g2648 ( 
.A(n_1987),
.Y(n_2648)
);

BUFx6f_ASAP7_75t_L g2649 ( 
.A(n_2220),
.Y(n_2649)
);

NAND2x1p5_ASAP7_75t_L g2650 ( 
.A(n_2244),
.B(n_115),
.Y(n_2650)
);

BUFx2_ASAP7_75t_SL g2651 ( 
.A(n_2261),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_SL g2652 ( 
.A(n_2162),
.B(n_114),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_L g2653 ( 
.A(n_2141),
.B(n_117),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_1967),
.B(n_117),
.Y(n_2654)
);

BUFx3_ASAP7_75t_L g2655 ( 
.A(n_2091),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_1967),
.B(n_1973),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2124),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_1973),
.B(n_118),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2218),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2217),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2003),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2129),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2193),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2010),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2024),
.Y(n_2665)
);

OR2x2_ASAP7_75t_L g2666 ( 
.A(n_2246),
.B(n_2238),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2249),
.B(n_2080),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_1993),
.B(n_119),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2193),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2268),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2151),
.B(n_120),
.Y(n_2671)
);

BUFx3_ASAP7_75t_L g2672 ( 
.A(n_2091),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2189),
.Y(n_2673)
);

AND2x4_ASAP7_75t_L g2674 ( 
.A(n_2100),
.B(n_120),
.Y(n_2674)
);

AND2x6_ASAP7_75t_L g2675 ( 
.A(n_2209),
.B(n_121),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_1993),
.B(n_122),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2189),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2192),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2100),
.B(n_123),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2087),
.B(n_124),
.Y(n_2680)
);

HB1xp67_ASAP7_75t_L g2681 ( 
.A(n_2087),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2258),
.B(n_124),
.Y(n_2682)
);

BUFx8_ASAP7_75t_SL g2683 ( 
.A(n_2164),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_1997),
.B(n_125),
.Y(n_2684)
);

BUFx4f_ASAP7_75t_L g2685 ( 
.A(n_2013),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_1997),
.B(n_125),
.Y(n_2686)
);

BUFx3_ASAP7_75t_L g2687 ( 
.A(n_2130),
.Y(n_2687)
);

OR2x6_ASAP7_75t_L g2688 ( 
.A(n_2210),
.B(n_126),
.Y(n_2688)
);

NAND2x1p5_ASAP7_75t_L g2689 ( 
.A(n_1986),
.B(n_128),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2192),
.Y(n_2690)
);

AND2x4_ASAP7_75t_L g2691 ( 
.A(n_2130),
.B(n_127),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2012),
.B(n_129),
.Y(n_2692)
);

BUFx8_ASAP7_75t_L g2693 ( 
.A(n_2251),
.Y(n_2693)
);

INVx6_ASAP7_75t_L g2694 ( 
.A(n_2089),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2137),
.Y(n_2695)
);

NOR2xp33_ASAP7_75t_L g2696 ( 
.A(n_2012),
.B(n_846),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_L g2697 ( 
.A(n_2026),
.B(n_848),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2089),
.B(n_129),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2137),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2216),
.Y(n_2700)
);

BUFx6f_ASAP7_75t_L g2701 ( 
.A(n_2261),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2184),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2159),
.B(n_130),
.Y(n_2703)
);

AND2x4_ASAP7_75t_L g2704 ( 
.A(n_2187),
.B(n_130),
.Y(n_2704)
);

INVx4_ASAP7_75t_L g2705 ( 
.A(n_2261),
.Y(n_2705)
);

CKINVDCx8_ASAP7_75t_R g2706 ( 
.A(n_2069),
.Y(n_2706)
);

BUFx12f_ASAP7_75t_L g2707 ( 
.A(n_1987),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2174),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2026),
.B(n_2031),
.Y(n_2709)
);

OR2x6_ASAP7_75t_L g2710 ( 
.A(n_2196),
.B(n_131),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2252),
.B(n_132),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2031),
.B(n_132),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2184),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2221),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2157),
.Y(n_2715)
);

AND2x6_ASAP7_75t_L g2716 ( 
.A(n_2235),
.B(n_2227),
.Y(n_2716)
);

INVx5_ASAP7_75t_L g2717 ( 
.A(n_2261),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2073),
.B(n_133),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_2261),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2174),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2033),
.B(n_133),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2181),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2188),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_1961),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_1961),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_1961),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2033),
.B(n_134),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2177),
.Y(n_2728)
);

INVxp67_ASAP7_75t_L g2729 ( 
.A(n_2208),
.Y(n_2729)
);

BUFx8_ASAP7_75t_SL g2730 ( 
.A(n_2167),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2127),
.B(n_134),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2127),
.B(n_135),
.Y(n_2732)
);

AND2x4_ASAP7_75t_L g2733 ( 
.A(n_2208),
.B(n_2069),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_1961),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2200),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2215),
.B(n_135),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2133),
.B(n_136),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2200),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2133),
.B(n_136),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2185),
.B(n_137),
.Y(n_2740)
);

INVx4_ASAP7_75t_L g2741 ( 
.A(n_1961),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2168),
.B(n_137),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2177),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2202),
.Y(n_2744)
);

NOR2xp33_ASAP7_75t_L g2745 ( 
.A(n_2092),
.B(n_834),
.Y(n_2745)
);

INVx8_ASAP7_75t_L g2746 ( 
.A(n_2248),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2169),
.Y(n_2747)
);

BUFx3_ASAP7_75t_L g2748 ( 
.A(n_2082),
.Y(n_2748)
);

INVx3_ASAP7_75t_L g2749 ( 
.A(n_2253),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2094),
.B(n_138),
.Y(n_2750)
);

INVx6_ASAP7_75t_L g2751 ( 
.A(n_2223),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2053),
.B(n_138),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2253),
.Y(n_2753)
);

AND2x4_ASAP7_75t_L g2754 ( 
.A(n_1963),
.B(n_140),
.Y(n_2754)
);

AO21x2_ASAP7_75t_L g2755 ( 
.A1(n_2264),
.A2(n_140),
.B(n_141),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2013),
.B(n_141),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2223),
.B(n_144),
.Y(n_2757)
);

OR2x6_ASAP7_75t_L g2758 ( 
.A(n_2219),
.B(n_145),
.Y(n_2758)
);

INVx1_ASAP7_75t_SL g2759 ( 
.A(n_2236),
.Y(n_2759)
);

BUFx6f_ASAP7_75t_L g2760 ( 
.A(n_2248),
.Y(n_2760)
);

NOR2x1_ASAP7_75t_R g2761 ( 
.A(n_1963),
.B(n_145),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2140),
.B(n_147),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2140),
.B(n_147),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2154),
.B(n_844),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2154),
.B(n_148),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2202),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2236),
.B(n_149),
.Y(n_2767)
);

NOR2x1_ASAP7_75t_L g2768 ( 
.A(n_2264),
.B(n_149),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2063),
.B(n_150),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2201),
.Y(n_2770)
);

OR2x6_ASAP7_75t_L g2771 ( 
.A(n_2219),
.B(n_150),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2248),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2063),
.B(n_825),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2241),
.B(n_151),
.Y(n_2774)
);

BUFx8_ASAP7_75t_L g2775 ( 
.A(n_2248),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2241),
.Y(n_2776)
);

NAND2x1p5_ASAP7_75t_L g2777 ( 
.A(n_2278),
.B(n_152),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2201),
.B(n_151),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2099),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2099),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2101),
.Y(n_2781)
);

BUFx12f_ASAP7_75t_L g2782 ( 
.A(n_2248),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2258),
.B(n_152),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2101),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2084),
.B(n_153),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2227),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2110),
.B(n_154),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2110),
.Y(n_2788)
);

OR2x2_ASAP7_75t_L g2789 ( 
.A(n_2084),
.B(n_154),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_1966),
.B(n_155),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_1966),
.B(n_155),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2123),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2269),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2269),
.Y(n_2794)
);

CKINVDCx5p33_ASAP7_75t_R g2795 ( 
.A(n_2021),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2123),
.Y(n_2796)
);

BUFx8_ASAP7_75t_SL g2797 ( 
.A(n_2046),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2009),
.B(n_156),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2009),
.B(n_156),
.Y(n_2799)
);

BUFx2_ASAP7_75t_L g2800 ( 
.A(n_2027),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2027),
.B(n_157),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2178),
.B(n_2239),
.Y(n_2802)
);

BUFx2_ASAP7_75t_L g2803 ( 
.A(n_2179),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2265),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2179),
.B(n_157),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2117),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2250),
.Y(n_2807)
);

OR2x6_ASAP7_75t_L g2808 ( 
.A(n_2259),
.B(n_159),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_1965),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2048),
.B(n_159),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_SL g2811 ( 
.A(n_1995),
.B(n_161),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_1994),
.B(n_837),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2122),
.B(n_161),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2048),
.B(n_162),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_1982),
.Y(n_2815)
);

OR2x6_ASAP7_75t_L g2816 ( 
.A(n_2104),
.B(n_162),
.Y(n_2816)
);

OR2x2_ASAP7_75t_L g2817 ( 
.A(n_1960),
.B(n_163),
.Y(n_2817)
);

AND2x4_ASAP7_75t_L g2818 ( 
.A(n_2120),
.B(n_163),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2122),
.B(n_164),
.Y(n_2819)
);

OR2x6_ASAP7_75t_L g2820 ( 
.A(n_2104),
.B(n_165),
.Y(n_2820)
);

OR2x2_ASAP7_75t_L g2821 ( 
.A(n_1960),
.B(n_165),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2120),
.B(n_166),
.Y(n_2822)
);

INVx1_ASAP7_75t_SL g2823 ( 
.A(n_1960),
.Y(n_2823)
);

BUFx6f_ASAP7_75t_L g2824 ( 
.A(n_1982),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2122),
.B(n_166),
.Y(n_2825)
);

BUFx12f_ASAP7_75t_L g2826 ( 
.A(n_2121),
.Y(n_2826)
);

CKINVDCx20_ASAP7_75t_R g2827 ( 
.A(n_1972),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2048),
.B(n_169),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_1965),
.Y(n_2829)
);

BUFx12f_ASAP7_75t_L g2830 ( 
.A(n_2121),
.Y(n_2830)
);

NAND2x1p5_ASAP7_75t_L g2831 ( 
.A(n_2120),
.B(n_170),
.Y(n_2831)
);

NAND2x1p5_ASAP7_75t_L g2832 ( 
.A(n_2120),
.B(n_170),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_1983),
.Y(n_2833)
);

BUFx5_ASAP7_75t_L g2834 ( 
.A(n_2261),
.Y(n_2834)
);

BUFx8_ASAP7_75t_SL g2835 ( 
.A(n_1972),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2048),
.B(n_169),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2291),
.Y(n_2837)
);

OR2x6_ASAP7_75t_L g2838 ( 
.A(n_2104),
.B(n_171),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_1994),
.B(n_826),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_1965),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_1964),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2048),
.B(n_171),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2122),
.B(n_172),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2120),
.B(n_172),
.Y(n_2844)
);

CKINVDCx16_ASAP7_75t_R g2845 ( 
.A(n_1972),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2048),
.B(n_173),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_1965),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2122),
.B(n_174),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2122),
.B(n_175),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_1982),
.Y(n_2850)
);

BUFx12f_ASAP7_75t_L g2851 ( 
.A(n_2121),
.Y(n_2851)
);

BUFx3_ASAP7_75t_L g2852 ( 
.A(n_2321),
.Y(n_2852)
);

BUFx3_ASAP7_75t_L g2853 ( 
.A(n_2321),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2835),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2310),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2310),
.Y(n_2856)
);

BUFx3_ASAP7_75t_L g2857 ( 
.A(n_2395),
.Y(n_2857)
);

BUFx3_ASAP7_75t_L g2858 ( 
.A(n_2312),
.Y(n_2858)
);

BUFx12f_ASAP7_75t_L g2859 ( 
.A(n_2826),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2368),
.A2(n_179),
.B1(n_176),
.B2(n_177),
.Y(n_2860)
);

INVx5_ASAP7_75t_L g2861 ( 
.A(n_2362),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2384),
.Y(n_2862)
);

BUFx2_ASAP7_75t_L g2863 ( 
.A(n_2326),
.Y(n_2863)
);

CKINVDCx20_ASAP7_75t_R g2864 ( 
.A(n_2827),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2319),
.A2(n_181),
.B1(n_176),
.B2(n_177),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2333),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_2830),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_L g2868 ( 
.A(n_2460),
.B(n_182),
.Y(n_2868)
);

INVx5_ASAP7_75t_L g2869 ( 
.A(n_2362),
.Y(n_2869)
);

BUFx8_ASAP7_75t_SL g2870 ( 
.A(n_2851),
.Y(n_2870)
);

BUFx5_ASAP7_75t_L g2871 ( 
.A(n_2314),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2314),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2841),
.Y(n_2873)
);

INVx8_ASAP7_75t_L g2874 ( 
.A(n_2320),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2457),
.B(n_182),
.Y(n_2875)
);

INVx4_ASAP7_75t_L g2876 ( 
.A(n_2312),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2351),
.Y(n_2877)
);

INVx4_ASAP7_75t_L g2878 ( 
.A(n_2326),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2779),
.B(n_183),
.Y(n_2879)
);

BUFx5_ASAP7_75t_L g2880 ( 
.A(n_2841),
.Y(n_2880)
);

BUFx6f_ASAP7_75t_L g2881 ( 
.A(n_2308),
.Y(n_2881)
);

CKINVDCx5p33_ASAP7_75t_R g2882 ( 
.A(n_2610),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_2308),
.Y(n_2883)
);

CKINVDCx8_ASAP7_75t_R g2884 ( 
.A(n_2320),
.Y(n_2884)
);

INVxp67_ASAP7_75t_SL g2885 ( 
.A(n_2337),
.Y(n_2885)
);

HB1xp67_ASAP7_75t_L g2886 ( 
.A(n_2353),
.Y(n_2886)
);

INVx1_ASAP7_75t_SL g2887 ( 
.A(n_2823),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2349),
.B(n_183),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2694),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2458),
.Y(n_2890)
);

CKINVDCx8_ASAP7_75t_R g2891 ( 
.A(n_2346),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2458),
.Y(n_2892)
);

INVx1_ASAP7_75t_SL g2893 ( 
.A(n_2694),
.Y(n_2893)
);

INVx5_ASAP7_75t_L g2894 ( 
.A(n_2362),
.Y(n_2894)
);

INVx5_ASAP7_75t_SL g2895 ( 
.A(n_2346),
.Y(n_2895)
);

OR2x6_ASAP7_75t_L g2896 ( 
.A(n_2600),
.B(n_184),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2337),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2375),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2464),
.Y(n_2899)
);

BUFx12f_ASAP7_75t_L g2900 ( 
.A(n_2393),
.Y(n_2900)
);

BUFx12f_ASAP7_75t_L g2901 ( 
.A(n_2340),
.Y(n_2901)
);

INVx5_ASAP7_75t_L g2902 ( 
.A(n_2367),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2543),
.Y(n_2903)
);

BUFx4f_ASAP7_75t_SL g2904 ( 
.A(n_2435),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2780),
.B(n_184),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2781),
.B(n_185),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2781),
.B(n_185),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2336),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2464),
.Y(n_2909)
);

BUFx4f_ASAP7_75t_L g2910 ( 
.A(n_2400),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2378),
.Y(n_2911)
);

BUFx3_ASAP7_75t_L g2912 ( 
.A(n_2833),
.Y(n_2912)
);

BUFx3_ASAP7_75t_L g2913 ( 
.A(n_2417),
.Y(n_2913)
);

INVx1_ASAP7_75t_SL g2914 ( 
.A(n_2307),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2364),
.Y(n_2915)
);

BUFx12f_ASAP7_75t_L g2916 ( 
.A(n_2340),
.Y(n_2916)
);

BUFx3_ASAP7_75t_L g2917 ( 
.A(n_2332),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_2364),
.Y(n_2918)
);

NAND2x1p5_ASAP7_75t_L g2919 ( 
.A(n_2407),
.B(n_186),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2809),
.Y(n_2920)
);

BUFx3_ASAP7_75t_L g2921 ( 
.A(n_2648),
.Y(n_2921)
);

BUFx3_ASAP7_75t_L g2922 ( 
.A(n_2707),
.Y(n_2922)
);

INVx8_ASAP7_75t_L g2923 ( 
.A(n_2318),
.Y(n_2923)
);

BUFx12f_ASAP7_75t_L g2924 ( 
.A(n_2517),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2470),
.Y(n_2925)
);

NAND2x1p5_ASAP7_75t_L g2926 ( 
.A(n_2407),
.B(n_187),
.Y(n_2926)
);

CKINVDCx6p67_ASAP7_75t_R g2927 ( 
.A(n_2400),
.Y(n_2927)
);

BUFx3_ASAP7_75t_L g2928 ( 
.A(n_2357),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2829),
.Y(n_2929)
);

BUFx3_ASAP7_75t_L g2930 ( 
.A(n_2439),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2443),
.Y(n_2931)
);

INVx1_ASAP7_75t_SL g2932 ( 
.A(n_2412),
.Y(n_2932)
);

INVx4_ASAP7_75t_L g2933 ( 
.A(n_2600),
.Y(n_2933)
);

CKINVDCx20_ASAP7_75t_R g2934 ( 
.A(n_2845),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2470),
.Y(n_2935)
);

BUFx12f_ASAP7_75t_L g2936 ( 
.A(n_2538),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2480),
.Y(n_2937)
);

BUFx12f_ASAP7_75t_L g2938 ( 
.A(n_2538),
.Y(n_2938)
);

INVx5_ASAP7_75t_L g2939 ( 
.A(n_2362),
.Y(n_2939)
);

BUFx2_ASAP7_75t_L g2940 ( 
.A(n_2415),
.Y(n_2940)
);

BUFx3_ASAP7_75t_L g2941 ( 
.A(n_2555),
.Y(n_2941)
);

INVx3_ASAP7_75t_SL g2942 ( 
.A(n_2845),
.Y(n_2942)
);

BUFx6f_ASAP7_75t_L g2943 ( 
.A(n_2308),
.Y(n_2943)
);

CKINVDCx16_ASAP7_75t_R g2944 ( 
.A(n_2419),
.Y(n_2944)
);

BUFx6f_ASAP7_75t_L g2945 ( 
.A(n_2328),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2480),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2510),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_2947)
);

AOI22xp33_ASAP7_75t_L g2948 ( 
.A1(n_2612),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_2948)
);

BUFx3_ASAP7_75t_L g2949 ( 
.A(n_2577),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2840),
.Y(n_2950)
);

BUFx12f_ASAP7_75t_L g2951 ( 
.A(n_2549),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2784),
.B(n_191),
.Y(n_2952)
);

CKINVDCx20_ASAP7_75t_R g2953 ( 
.A(n_2683),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2427),
.Y(n_2954)
);

BUFx12f_ASAP7_75t_L g2955 ( 
.A(n_2549),
.Y(n_2955)
);

INVx6_ASAP7_75t_SL g2956 ( 
.A(n_2318),
.Y(n_2956)
);

BUFx2_ASAP7_75t_SL g2957 ( 
.A(n_2633),
.Y(n_2957)
);

BUFx12f_ASAP7_75t_L g2958 ( 
.A(n_2567),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2482),
.Y(n_2959)
);

INVx5_ASAP7_75t_L g2960 ( 
.A(n_2367),
.Y(n_2960)
);

INVx1_ASAP7_75t_SL g2961 ( 
.A(n_2412),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2328),
.Y(n_2962)
);

INVx1_ASAP7_75t_SL g2963 ( 
.A(n_2541),
.Y(n_2963)
);

BUFx4_ASAP7_75t_SL g2964 ( 
.A(n_2567),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2847),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2427),
.Y(n_2966)
);

BUFx10_ASAP7_75t_L g2967 ( 
.A(n_2816),
.Y(n_2967)
);

INVx3_ASAP7_75t_L g2968 ( 
.A(n_2741),
.Y(n_2968)
);

CKINVDCx20_ASAP7_75t_R g2969 ( 
.A(n_2730),
.Y(n_2969)
);

CKINVDCx20_ASAP7_75t_R g2970 ( 
.A(n_2706),
.Y(n_2970)
);

BUFx3_ASAP7_75t_L g2971 ( 
.A(n_2389),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2482),
.Y(n_2972)
);

BUFx3_ASAP7_75t_L g2973 ( 
.A(n_2448),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2494),
.Y(n_2974)
);

CKINVDCx20_ASAP7_75t_R g2975 ( 
.A(n_2693),
.Y(n_2975)
);

INVxp67_ASAP7_75t_SL g2976 ( 
.A(n_2476),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2424),
.Y(n_2977)
);

CKINVDCx20_ASAP7_75t_R g2978 ( 
.A(n_2693),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2328),
.Y(n_2979)
);

BUFx12f_ASAP7_75t_L g2980 ( 
.A(n_2578),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2741),
.Y(n_2981)
);

INVx3_ASAP7_75t_L g2982 ( 
.A(n_2511),
.Y(n_2982)
);

BUFx6f_ASAP7_75t_L g2983 ( 
.A(n_2334),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2319),
.A2(n_2313),
.B1(n_2811),
.B2(n_2366),
.Y(n_2984)
);

BUFx12f_ASAP7_75t_L g2985 ( 
.A(n_2578),
.Y(n_2985)
);

INVx1_ASAP7_75t_SL g2986 ( 
.A(n_2459),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2533),
.B(n_192),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2733),
.B(n_192),
.Y(n_2988)
);

BUFx2_ASAP7_75t_SL g2989 ( 
.A(n_2367),
.Y(n_2989)
);

CKINVDCx16_ASAP7_75t_R g2990 ( 
.A(n_2434),
.Y(n_2990)
);

BUFx2_ASAP7_75t_L g2991 ( 
.A(n_2415),
.Y(n_2991)
);

CKINVDCx16_ASAP7_75t_R g2992 ( 
.A(n_2621),
.Y(n_2992)
);

OAI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2476),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_2993)
);

BUFx6f_ASAP7_75t_L g2994 ( 
.A(n_2334),
.Y(n_2994)
);

INVxp67_ASAP7_75t_SL g2995 ( 
.A(n_2495),
.Y(n_2995)
);

BUFx4f_ASAP7_75t_SL g2996 ( 
.A(n_2598),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2425),
.Y(n_2997)
);

INVx2_ASAP7_75t_SL g2998 ( 
.A(n_2495),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2595),
.Y(n_2999)
);

INVx1_ASAP7_75t_SL g3000 ( 
.A(n_2547),
.Y(n_3000)
);

BUFx3_ASAP7_75t_L g3001 ( 
.A(n_2360),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2494),
.Y(n_3002)
);

INVx8_ASAP7_75t_L g3003 ( 
.A(n_2621),
.Y(n_3003)
);

INVxp67_ASAP7_75t_SL g3004 ( 
.A(n_2652),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2334),
.Y(n_3005)
);

INVx1_ASAP7_75t_SL g3006 ( 
.A(n_2564),
.Y(n_3006)
);

NAND2x1p5_ASAP7_75t_L g3007 ( 
.A(n_2475),
.B(n_195),
.Y(n_3007)
);

BUFx6f_ASAP7_75t_L g3008 ( 
.A(n_2339),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2429),
.Y(n_3009)
);

BUFx6f_ASAP7_75t_SL g3010 ( 
.A(n_2816),
.Y(n_3010)
);

INVx3_ASAP7_75t_SL g3011 ( 
.A(n_2820),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2315),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2315),
.Y(n_3013)
);

BUFx2_ASAP7_75t_SL g3014 ( 
.A(n_2367),
.Y(n_3014)
);

INVx1_ASAP7_75t_SL g3015 ( 
.A(n_2418),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2733),
.B(n_196),
.Y(n_3016)
);

BUFx3_ASAP7_75t_L g3017 ( 
.A(n_2394),
.Y(n_3017)
);

NAND2x1p5_ASAP7_75t_L g3018 ( 
.A(n_2475),
.B(n_197),
.Y(n_3018)
);

INVx1_ASAP7_75t_SL g3019 ( 
.A(n_2418),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2784),
.B(n_2788),
.Y(n_3020)
);

BUFx2_ASAP7_75t_L g3021 ( 
.A(n_2449),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2477),
.B(n_198),
.Y(n_3022)
);

BUFx12f_ASAP7_75t_L g3023 ( 
.A(n_2820),
.Y(n_3023)
);

INVx5_ASAP7_75t_L g3024 ( 
.A(n_2585),
.Y(n_3024)
);

BUFx6f_ASAP7_75t_SL g3025 ( 
.A(n_2838),
.Y(n_3025)
);

INVx8_ASAP7_75t_L g3026 ( 
.A(n_2838),
.Y(n_3026)
);

INVx4_ASAP7_75t_L g3027 ( 
.A(n_2449),
.Y(n_3027)
);

INVxp67_ASAP7_75t_SL g3028 ( 
.A(n_2652),
.Y(n_3028)
);

NAND2x1p5_ASAP7_75t_L g3029 ( 
.A(n_2475),
.B(n_2498),
.Y(n_3029)
);

BUFx6f_ASAP7_75t_L g3030 ( 
.A(n_2339),
.Y(n_3030)
);

CKINVDCx6p67_ASAP7_75t_R g3031 ( 
.A(n_2595),
.Y(n_3031)
);

INVx2_ASAP7_75t_SL g3032 ( 
.A(n_2325),
.Y(n_3032)
);

BUFx3_ASAP7_75t_L g3033 ( 
.A(n_2430),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2456),
.Y(n_3034)
);

NAND2x1p5_ASAP7_75t_L g3035 ( 
.A(n_2498),
.B(n_198),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2339),
.Y(n_3036)
);

BUFx3_ASAP7_75t_L g3037 ( 
.A(n_2423),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2788),
.B(n_199),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2568),
.B(n_200),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2388),
.B(n_200),
.Y(n_3040)
);

INVx3_ASAP7_75t_L g3041 ( 
.A(n_2511),
.Y(n_3041)
);

INVx3_ASAP7_75t_L g3042 ( 
.A(n_2514),
.Y(n_3042)
);

BUFx6f_ASAP7_75t_L g3043 ( 
.A(n_2361),
.Y(n_3043)
);

INVx1_ASAP7_75t_SL g3044 ( 
.A(n_2626),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2373),
.B(n_201),
.Y(n_3045)
);

INVx1_ASAP7_75t_SL g3046 ( 
.A(n_2627),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2361),
.Y(n_3047)
);

INVx1_ASAP7_75t_SL g3048 ( 
.A(n_2632),
.Y(n_3048)
);

AOI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_2366),
.A2(n_2785),
.B1(n_2461),
.B2(n_2447),
.Y(n_3049)
);

BUFx5_ASAP7_75t_L g3050 ( 
.A(n_2591),
.Y(n_3050)
);

BUFx2_ASAP7_75t_SL g3051 ( 
.A(n_2585),
.Y(n_3051)
);

INVx6_ASAP7_75t_SL g3052 ( 
.A(n_2688),
.Y(n_3052)
);

BUFx3_ASAP7_75t_L g3053 ( 
.A(n_2504),
.Y(n_3053)
);

NAND2x1p5_ASAP7_75t_L g3054 ( 
.A(n_2498),
.B(n_202),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2519),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2462),
.Y(n_3056)
);

BUFx5_ASAP7_75t_L g3057 ( 
.A(n_2591),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_2666),
.B(n_203),
.Y(n_3058)
);

AOI22xp5_ASAP7_75t_L g3059 ( 
.A1(n_2785),
.A2(n_2461),
.B1(n_2468),
.B2(n_2309),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_L g3060 ( 
.A(n_2361),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2317),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2576),
.B(n_203),
.Y(n_3062)
);

INVx1_ASAP7_75t_SL g3063 ( 
.A(n_2405),
.Y(n_3063)
);

BUFx6f_ASAP7_75t_L g3064 ( 
.A(n_2392),
.Y(n_3064)
);

AOI22xp5_ASAP7_75t_L g3065 ( 
.A1(n_2776),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_L g3066 ( 
.A(n_2392),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_SL g3067 ( 
.A(n_2758),
.Y(n_3067)
);

INVx1_ASAP7_75t_SL g3068 ( 
.A(n_2405),
.Y(n_3068)
);

CKINVDCx20_ASAP7_75t_R g3069 ( 
.A(n_2797),
.Y(n_3069)
);

INVxp67_ASAP7_75t_SL g3070 ( 
.A(n_2754),
.Y(n_3070)
);

BUFx2_ASAP7_75t_L g3071 ( 
.A(n_2775),
.Y(n_3071)
);

INVx2_ASAP7_75t_SL g3072 ( 
.A(n_2748),
.Y(n_3072)
);

INVx3_ASAP7_75t_SL g3073 ( 
.A(n_2747),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2473),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2656),
.B(n_206),
.Y(n_3075)
);

BUFx3_ASAP7_75t_L g3076 ( 
.A(n_2581),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2647),
.Y(n_3077)
);

BUFx3_ASAP7_75t_L g3078 ( 
.A(n_2655),
.Y(n_3078)
);

BUFx6f_ASAP7_75t_L g3079 ( 
.A(n_2392),
.Y(n_3079)
);

INVx8_ASAP7_75t_L g3080 ( 
.A(n_2710),
.Y(n_3080)
);

INVx2_ASAP7_75t_SL g3081 ( 
.A(n_2631),
.Y(n_3081)
);

INVx4_ASAP7_75t_L g3082 ( 
.A(n_2502),
.Y(n_3082)
);

INVx2_ASAP7_75t_SL g3083 ( 
.A(n_2631),
.Y(n_3083)
);

BUFx4_ASAP7_75t_SL g3084 ( 
.A(n_2758),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2478),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2317),
.Y(n_3086)
);

INVx3_ASAP7_75t_L g3087 ( 
.A(n_2514),
.Y(n_3087)
);

BUFx4f_ASAP7_75t_SL g3088 ( 
.A(n_2775),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_2672),
.Y(n_3089)
);

BUFx6f_ASAP7_75t_L g3090 ( 
.A(n_2404),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2404),
.Y(n_3091)
);

HB1xp67_ASAP7_75t_L g3092 ( 
.A(n_2710),
.Y(n_3092)
);

NAND2x1p5_ASAP7_75t_L g3093 ( 
.A(n_2502),
.B(n_207),
.Y(n_3093)
);

INVx6_ASAP7_75t_L g3094 ( 
.A(n_2688),
.Y(n_3094)
);

INVx3_ASAP7_75t_L g3095 ( 
.A(n_2562),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2487),
.Y(n_3096)
);

HB1xp67_ASAP7_75t_L g3097 ( 
.A(n_2570),
.Y(n_3097)
);

INVx1_ASAP7_75t_SL g3098 ( 
.A(n_2372),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2348),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_2562),
.Y(n_3100)
);

BUFx3_ASAP7_75t_L g3101 ( 
.A(n_2687),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_2601),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2348),
.Y(n_3103)
);

BUFx2_ASAP7_75t_L g3104 ( 
.A(n_2391),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_2622),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2352),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2352),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2491),
.Y(n_3108)
);

BUFx3_ASAP7_75t_L g3109 ( 
.A(n_2372),
.Y(n_3109)
);

INVx8_ASAP7_75t_L g3110 ( 
.A(n_2585),
.Y(n_3110)
);

INVx6_ASAP7_75t_SL g3111 ( 
.A(n_2501),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2497),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2525),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_2329),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2354),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2354),
.Y(n_3116)
);

BUFx4f_ASAP7_75t_SL g3117 ( 
.A(n_2782),
.Y(n_3117)
);

BUFx3_ASAP7_75t_L g3118 ( 
.A(n_2715),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2722),
.Y(n_3119)
);

INVx1_ASAP7_75t_SL g3120 ( 
.A(n_2329),
.Y(n_3120)
);

AOI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2653),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_3121)
);

NOR2xp67_ASAP7_75t_SL g3122 ( 
.A(n_2651),
.B(n_209),
.Y(n_3122)
);

INVx6_ASAP7_75t_SL g3123 ( 
.A(n_2501),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2376),
.Y(n_3124)
);

AO22x2_ASAP7_75t_L g3125 ( 
.A1(n_2754),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2376),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2404),
.Y(n_3127)
);

BUFx3_ASAP7_75t_L g3128 ( 
.A(n_2311),
.Y(n_3128)
);

BUFx12f_ASAP7_75t_L g3129 ( 
.A(n_2771),
.Y(n_3129)
);

CKINVDCx20_ASAP7_75t_R g3130 ( 
.A(n_2341),
.Y(n_3130)
);

INVx4_ASAP7_75t_L g3131 ( 
.A(n_2502),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2311),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2399),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2709),
.B(n_211),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2670),
.B(n_212),
.Y(n_3135)
);

INVx3_ASAP7_75t_SL g3136 ( 
.A(n_2771),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2399),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2414),
.Y(n_3138)
);

INVxp67_ASAP7_75t_SL g3139 ( 
.A(n_2433),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2744),
.B(n_213),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2316),
.B(n_2323),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2667),
.B(n_214),
.Y(n_3142)
);

INVx5_ASAP7_75t_L g3143 ( 
.A(n_2585),
.Y(n_3143)
);

NAND2x1p5_ASAP7_75t_L g3144 ( 
.A(n_2685),
.B(n_214),
.Y(n_3144)
);

BUFx3_ASAP7_75t_L g3145 ( 
.A(n_2358),
.Y(n_3145)
);

INVx3_ASAP7_75t_SL g3146 ( 
.A(n_2508),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2381),
.B(n_216),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2582),
.Y(n_3148)
);

HB1xp67_ASAP7_75t_L g3149 ( 
.A(n_2614),
.Y(n_3149)
);

INVx3_ASAP7_75t_L g3150 ( 
.A(n_2622),
.Y(n_3150)
);

BUFx3_ASAP7_75t_L g3151 ( 
.A(n_2358),
.Y(n_3151)
);

BUFx6f_ASAP7_75t_L g3152 ( 
.A(n_2414),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2681),
.B(n_216),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2582),
.Y(n_3154)
);

BUFx3_ASAP7_75t_L g3155 ( 
.A(n_2837),
.Y(n_3155)
);

BUFx3_ASAP7_75t_L g3156 ( 
.A(n_2837),
.Y(n_3156)
);

INVx3_ASAP7_75t_L g3157 ( 
.A(n_2663),
.Y(n_3157)
);

AOI22xp33_ASAP7_75t_L g3158 ( 
.A1(n_2685),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_3158)
);

INVx6_ASAP7_75t_L g3159 ( 
.A(n_2345),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2575),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_2624),
.B(n_218),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2588),
.Y(n_3162)
);

INVx5_ASAP7_75t_L g3163 ( 
.A(n_2746),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2744),
.B(n_219),
.Y(n_3164)
);

BUFx6f_ASAP7_75t_L g3165 ( 
.A(n_2414),
.Y(n_3165)
);

BUFx2_ASAP7_75t_R g3166 ( 
.A(n_2795),
.Y(n_3166)
);

INVx4_ASAP7_75t_L g3167 ( 
.A(n_2746),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2588),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2724),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2421),
.B(n_223),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2689),
.Y(n_3171)
);

BUFx8_ASAP7_75t_L g3172 ( 
.A(n_2532),
.Y(n_3172)
);

INVxp67_ASAP7_75t_SL g3173 ( 
.A(n_2618),
.Y(n_3173)
);

BUFx6f_ASAP7_75t_L g3174 ( 
.A(n_2428),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2499),
.Y(n_3175)
);

BUFx24_ASAP7_75t_L g3176 ( 
.A(n_2474),
.Y(n_3176)
);

BUFx8_ASAP7_75t_L g3177 ( 
.A(n_2408),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2759),
.B(n_224),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2499),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2422),
.B(n_224),
.Y(n_3180)
);

INVx3_ASAP7_75t_L g3181 ( 
.A(n_2663),
.Y(n_3181)
);

BUFx2_ASAP7_75t_L g3182 ( 
.A(n_2729),
.Y(n_3182)
);

BUFx3_ASAP7_75t_L g3183 ( 
.A(n_2592),
.Y(n_3183)
);

CKINVDCx5p33_ASAP7_75t_R g3184 ( 
.A(n_2508),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2505),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2413),
.Y(n_3186)
);

INVx3_ASAP7_75t_L g3187 ( 
.A(n_2663),
.Y(n_3187)
);

INVx6_ASAP7_75t_L g3188 ( 
.A(n_2345),
.Y(n_3188)
);

INVx3_ASAP7_75t_L g3189 ( 
.A(n_2669),
.Y(n_3189)
);

BUFx3_ASAP7_75t_L g3190 ( 
.A(n_2438),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2505),
.Y(n_3191)
);

AOI22xp33_ASAP7_75t_L g3192 ( 
.A1(n_2751),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_3192)
);

BUFx3_ASAP7_75t_L g3193 ( 
.A(n_2438),
.Y(n_3193)
);

INVx1_ASAP7_75t_SL g3194 ( 
.A(n_2817),
.Y(n_3194)
);

CKINVDCx20_ASAP7_75t_R g3195 ( 
.A(n_2342),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2512),
.Y(n_3196)
);

BUFx3_ASAP7_75t_L g3197 ( 
.A(n_2674),
.Y(n_3197)
);

CKINVDCx5p33_ASAP7_75t_R g3198 ( 
.A(n_2637),
.Y(n_3198)
);

CKINVDCx20_ASAP7_75t_R g3199 ( 
.A(n_2420),
.Y(n_3199)
);

BUFx2_ASAP7_75t_SL g3200 ( 
.A(n_2717),
.Y(n_3200)
);

CKINVDCx5p33_ASAP7_75t_R g3201 ( 
.A(n_2637),
.Y(n_3201)
);

INVx1_ASAP7_75t_SL g3202 ( 
.A(n_2483),
.Y(n_3202)
);

CKINVDCx8_ASAP7_75t_R g3203 ( 
.A(n_2675),
.Y(n_3203)
);

BUFx2_ASAP7_75t_L g3204 ( 
.A(n_2675),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2674),
.Y(n_3205)
);

INVx5_ASAP7_75t_L g3206 ( 
.A(n_2428),
.Y(n_3206)
);

NAND2x1p5_ASAP7_75t_L g3207 ( 
.A(n_2705),
.B(n_225),
.Y(n_3207)
);

BUFx3_ASAP7_75t_L g3208 ( 
.A(n_2679),
.Y(n_3208)
);

BUFx8_ASAP7_75t_L g3209 ( 
.A(n_2408),
.Y(n_3209)
);

INVx5_ASAP7_75t_L g3210 ( 
.A(n_2428),
.Y(n_3210)
);

INVx3_ASAP7_75t_SL g3211 ( 
.A(n_2411),
.Y(n_3211)
);

BUFx3_ASAP7_75t_L g3212 ( 
.A(n_2679),
.Y(n_3212)
);

INVx3_ASAP7_75t_SL g3213 ( 
.A(n_2411),
.Y(n_3213)
);

INVx3_ASAP7_75t_L g3214 ( 
.A(n_2669),
.Y(n_3214)
);

INVx3_ASAP7_75t_SL g3215 ( 
.A(n_2818),
.Y(n_3215)
);

BUFx2_ASAP7_75t_L g3216 ( 
.A(n_2675),
.Y(n_3216)
);

INVx5_ASAP7_75t_L g3217 ( 
.A(n_2444),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2512),
.Y(n_3218)
);

AND2x4_ASAP7_75t_L g3219 ( 
.A(n_2624),
.B(n_226),
.Y(n_3219)
);

INVx2_ASAP7_75t_SL g3220 ( 
.A(n_2691),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2515),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2609),
.Y(n_3222)
);

INVx3_ASAP7_75t_L g3223 ( 
.A(n_2669),
.Y(n_3223)
);

BUFx2_ASAP7_75t_L g3224 ( 
.A(n_2675),
.Y(n_3224)
);

INVx5_ASAP7_75t_L g3225 ( 
.A(n_2444),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_2444),
.Y(n_3226)
);

CKINVDCx16_ASAP7_75t_R g3227 ( 
.A(n_2472),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2617),
.Y(n_3228)
);

AND2x4_ASAP7_75t_L g3229 ( 
.A(n_2625),
.B(n_227),
.Y(n_3229)
);

BUFx10_ASAP7_75t_L g3230 ( 
.A(n_2818),
.Y(n_3230)
);

INVx1_ASAP7_75t_SL g3231 ( 
.A(n_2821),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_L g3232 ( 
.A1(n_2751),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_3232)
);

BUFx5_ASAP7_75t_L g3233 ( 
.A(n_2594),
.Y(n_3233)
);

INVx3_ASAP7_75t_L g3234 ( 
.A(n_2724),
.Y(n_3234)
);

BUFx3_ASAP7_75t_L g3235 ( 
.A(n_2691),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2515),
.Y(n_3236)
);

OR2x2_ASAP7_75t_L g3237 ( 
.A(n_2436),
.B(n_229),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2454),
.B(n_230),
.Y(n_3238)
);

OR2x2_ASAP7_75t_L g3239 ( 
.A(n_2463),
.B(n_231),
.Y(n_3239)
);

BUFx2_ASAP7_75t_L g3240 ( 
.A(n_2761),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_SL g3241 ( 
.A(n_2507),
.Y(n_3241)
);

AND2x6_ASAP7_75t_L g3242 ( 
.A(n_2724),
.B(n_232),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_2815),
.Y(n_3243)
);

INVx1_ASAP7_75t_SL g3244 ( 
.A(n_2523),
.Y(n_3244)
);

INVx1_ASAP7_75t_SL g3245 ( 
.A(n_2583),
.Y(n_3245)
);

NAND2x1p5_ASAP7_75t_L g3246 ( 
.A(n_2705),
.B(n_2717),
.Y(n_3246)
);

CKINVDCx20_ASAP7_75t_R g3247 ( 
.A(n_2711),
.Y(n_3247)
);

BUFx3_ASAP7_75t_L g3248 ( 
.A(n_2496),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_2530),
.B(n_232),
.Y(n_3249)
);

CKINVDCx20_ASAP7_75t_R g3250 ( 
.A(n_2350),
.Y(n_3250)
);

BUFx2_ASAP7_75t_L g3251 ( 
.A(n_2761),
.Y(n_3251)
);

BUFx2_ASAP7_75t_SL g3252 ( 
.A(n_2717),
.Y(n_3252)
);

BUFx2_ASAP7_75t_L g3253 ( 
.A(n_2822),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2620),
.Y(n_3254)
);

BUFx3_ASAP7_75t_L g3255 ( 
.A(n_2465),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_2465),
.Y(n_3256)
);

INVx3_ASAP7_75t_L g3257 ( 
.A(n_2725),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2516),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2630),
.Y(n_3259)
);

BUFx2_ASAP7_75t_R g3260 ( 
.A(n_2755),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2636),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_2642),
.B(n_233),
.Y(n_3262)
);

BUFx3_ASAP7_75t_L g3263 ( 
.A(n_2493),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2516),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2518),
.Y(n_3265)
);

BUFx4f_ASAP7_75t_SL g3266 ( 
.A(n_2490),
.Y(n_3266)
);

BUFx12f_ASAP7_75t_SL g3267 ( 
.A(n_2474),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2725),
.Y(n_3268)
);

INVx5_ASAP7_75t_L g3269 ( 
.A(n_2815),
.Y(n_3269)
);

INVx3_ASAP7_75t_L g3270 ( 
.A(n_2725),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2518),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2528),
.Y(n_3272)
);

BUFx12f_ASAP7_75t_L g3273 ( 
.A(n_2509),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_2493),
.Y(n_3274)
);

OR2x2_ASAP7_75t_L g3275 ( 
.A(n_2539),
.B(n_234),
.Y(n_3275)
);

BUFx3_ASAP7_75t_L g3276 ( 
.A(n_2561),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2646),
.Y(n_3277)
);

OR2x6_ASAP7_75t_L g3278 ( 
.A(n_2645),
.B(n_235),
.Y(n_3278)
);

BUFx12f_ASAP7_75t_L g3279 ( 
.A(n_2822),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_2359),
.B(n_235),
.Y(n_3280)
);

AOI22xp5_ASAP7_75t_L g3281 ( 
.A1(n_2410),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3281)
);

BUFx3_ASAP7_75t_L g3282 ( 
.A(n_2561),
.Y(n_3282)
);

BUFx6f_ASAP7_75t_L g3283 ( 
.A(n_2815),
.Y(n_3283)
);

BUFx8_ASAP7_75t_L g3284 ( 
.A(n_2574),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2657),
.Y(n_3285)
);

NAND2x1p5_ASAP7_75t_L g3286 ( 
.A(n_2583),
.B(n_236),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2662),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2432),
.B(n_237),
.Y(n_3288)
);

BUFx4f_ASAP7_75t_L g3289 ( 
.A(n_2650),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2639),
.B(n_2528),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2605),
.Y(n_3291)
);

INVx2_ASAP7_75t_SL g3292 ( 
.A(n_2597),
.Y(n_3292)
);

BUFx2_ASAP7_75t_L g3293 ( 
.A(n_2844),
.Y(n_3293)
);

BUFx4f_ASAP7_75t_L g3294 ( 
.A(n_2831),
.Y(n_3294)
);

BUFx3_ASAP7_75t_L g3295 ( 
.A(n_2611),
.Y(n_3295)
);

BUFx12f_ASAP7_75t_L g3296 ( 
.A(n_2844),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2529),
.Y(n_3297)
);

INVx1_ASAP7_75t_SL g3298 ( 
.A(n_2597),
.Y(n_3298)
);

INVx1_ASAP7_75t_SL g3299 ( 
.A(n_2604),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2605),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_2824),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_2450),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_3302)
);

BUFx12f_ASAP7_75t_L g3303 ( 
.A(n_2387),
.Y(n_3303)
);

INVx5_ASAP7_75t_L g3304 ( 
.A(n_2824),
.Y(n_3304)
);

INVx5_ASAP7_75t_L g3305 ( 
.A(n_2824),
.Y(n_3305)
);

INVx3_ASAP7_75t_L g3306 ( 
.A(n_2726),
.Y(n_3306)
);

INVx5_ASAP7_75t_L g3307 ( 
.A(n_2850),
.Y(n_3307)
);

AND2x4_ASAP7_75t_L g3308 ( 
.A(n_2625),
.B(n_239),
.Y(n_3308)
);

NAND2x1p5_ASAP7_75t_L g3309 ( 
.A(n_2703),
.B(n_242),
.Y(n_3309)
);

INVx2_ASAP7_75t_SL g3310 ( 
.A(n_2387),
.Y(n_3310)
);

BUFx12f_ASAP7_75t_L g3311 ( 
.A(n_2398),
.Y(n_3311)
);

CKINVDCx5p33_ASAP7_75t_R g3312 ( 
.A(n_2409),
.Y(n_3312)
);

BUFx6f_ASAP7_75t_L g3313 ( 
.A(n_2850),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_2406),
.B(n_2431),
.Y(n_3314)
);

BUFx12f_ASAP7_75t_L g3315 ( 
.A(n_2398),
.Y(n_3315)
);

INVx4_ASAP7_75t_L g3316 ( 
.A(n_2726),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2529),
.Y(n_3317)
);

BUFx6f_ASAP7_75t_L g3318 ( 
.A(n_2850),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_2558),
.Y(n_3319)
);

INVx1_ASAP7_75t_SL g3320 ( 
.A(n_2607),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2558),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2571),
.Y(n_3322)
);

BUFx2_ASAP7_75t_L g3323 ( 
.A(n_2371),
.Y(n_3323)
);

OAI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3049),
.A2(n_2643),
.B1(n_2565),
.B2(n_2481),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3291),
.Y(n_3325)
);

CKINVDCx11_ASAP7_75t_R g3326 ( 
.A(n_2854),
.Y(n_3326)
);

BUFx2_ASAP7_75t_L g3327 ( 
.A(n_2956),
.Y(n_3327)
);

BUFx12f_ASAP7_75t_L g3328 ( 
.A(n_2859),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2890),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2890),
.Y(n_3330)
);

CKINVDCx16_ASAP7_75t_R g3331 ( 
.A(n_2975),
.Y(n_3331)
);

CKINVDCx11_ASAP7_75t_R g3332 ( 
.A(n_2924),
.Y(n_3332)
);

INVxp67_ASAP7_75t_SL g3333 ( 
.A(n_3070),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_2910),
.A2(n_2643),
.B1(n_2565),
.B2(n_2812),
.Y(n_3334)
);

CKINVDCx11_ASAP7_75t_R g3335 ( 
.A(n_2978),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_SL g3336 ( 
.A1(n_3003),
.A2(n_2628),
.B1(n_2472),
.B2(n_2756),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3175),
.B(n_2762),
.Y(n_3337)
);

AOI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_2910),
.A2(n_2839),
.B1(n_2534),
.B2(n_2757),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_SL g3339 ( 
.A1(n_3003),
.A2(n_2537),
.B1(n_2481),
.B2(n_2522),
.Y(n_3339)
);

CKINVDCx11_ASAP7_75t_R g3340 ( 
.A(n_2864),
.Y(n_3340)
);

BUFx4_ASAP7_75t_SL g3341 ( 
.A(n_2953),
.Y(n_3341)
);

OAI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3049),
.A2(n_2522),
.B1(n_2507),
.B2(n_2545),
.Y(n_3342)
);

INVxp67_ASAP7_75t_SL g3343 ( 
.A(n_3173),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_3300),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3175),
.B(n_2383),
.Y(n_3345)
);

NAND2x1p5_ASAP7_75t_L g3346 ( 
.A(n_2876),
.B(n_2703),
.Y(n_3346)
);

INVx5_ASAP7_75t_L g3347 ( 
.A(n_2896),
.Y(n_3347)
);

AOI22xp33_ASAP7_75t_L g3348 ( 
.A1(n_3067),
.A2(n_2764),
.B1(n_2800),
.B2(n_2745),
.Y(n_3348)
);

OAI22xp33_ASAP7_75t_L g3349 ( 
.A1(n_2992),
.A2(n_2790),
.B1(n_2799),
.B2(n_2789),
.Y(n_3349)
);

INVx2_ASAP7_75t_SL g3350 ( 
.A(n_2904),
.Y(n_3350)
);

INVx3_ASAP7_75t_L g3351 ( 
.A(n_3203),
.Y(n_3351)
);

OAI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_2992),
.A2(n_2832),
.B1(n_2769),
.B2(n_2380),
.Y(n_3352)
);

BUFx10_ASAP7_75t_L g3353 ( 
.A(n_3010),
.Y(n_3353)
);

BUFx8_ASAP7_75t_SL g3354 ( 
.A(n_2870),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3012),
.Y(n_3355)
);

INVx6_ASAP7_75t_L g3356 ( 
.A(n_2876),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_SL g3357 ( 
.A1(n_2984),
.A2(n_2783),
.B(n_2489),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3012),
.Y(n_3358)
);

BUFx12f_ASAP7_75t_L g3359 ( 
.A(n_2867),
.Y(n_3359)
);

BUFx10_ASAP7_75t_L g3360 ( 
.A(n_3010),
.Y(n_3360)
);

BUFx2_ASAP7_75t_L g3361 ( 
.A(n_2956),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3013),
.Y(n_3362)
);

BUFx3_ASAP7_75t_L g3363 ( 
.A(n_2857),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_2964),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3179),
.B(n_2639),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3013),
.Y(n_3366)
);

CKINVDCx11_ASAP7_75t_R g3367 ( 
.A(n_2884),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_3067),
.A2(n_2738),
.B1(n_2766),
.B2(n_2735),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3314),
.B(n_2441),
.Y(n_3369)
);

OAI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_2896),
.A2(n_2712),
.B1(n_2503),
.B2(n_2808),
.Y(n_3370)
);

INVx5_ASAP7_75t_L g3371 ( 
.A(n_2874),
.Y(n_3371)
);

INVx4_ASAP7_75t_L g3372 ( 
.A(n_3110),
.Y(n_3372)
);

BUFx12f_ASAP7_75t_L g3373 ( 
.A(n_2862),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2866),
.Y(n_3374)
);

OAI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_2944),
.A2(n_2808),
.B1(n_2485),
.B2(n_2521),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_2984),
.A2(n_2545),
.B1(n_2556),
.B2(n_2551),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_2933),
.A2(n_3240),
.B1(n_3251),
.B2(n_3027),
.Y(n_3377)
);

AOI22xp33_ASAP7_75t_L g3378 ( 
.A1(n_2933),
.A2(n_3027),
.B1(n_3025),
.B2(n_3129),
.Y(n_3378)
);

INVx2_ASAP7_75t_SL g3379 ( 
.A(n_2858),
.Y(n_3379)
);

INVx6_ASAP7_75t_L g3380 ( 
.A(n_3172),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_3025),
.A2(n_2770),
.B1(n_2638),
.B2(n_2641),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3061),
.Y(n_3382)
);

BUFx6f_ASAP7_75t_L g3383 ( 
.A(n_3029),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3059),
.A2(n_2644),
.B1(n_2608),
.B2(n_2696),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3059),
.A2(n_2551),
.B1(n_2560),
.B2(n_2556),
.Y(n_3385)
);

CKINVDCx20_ASAP7_75t_R g3386 ( 
.A(n_2969),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2877),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_SL g3388 ( 
.A1(n_2891),
.A2(n_2489),
.B1(n_2704),
.B2(n_2752),
.Y(n_3388)
);

INVx2_ASAP7_75t_SL g3389 ( 
.A(n_2874),
.Y(n_3389)
);

OAI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_2944),
.A2(n_2990),
.B1(n_2927),
.B2(n_3227),
.Y(n_3390)
);

BUFx8_ASAP7_75t_SL g3391 ( 
.A(n_2900),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_2963),
.B(n_2363),
.Y(n_3392)
);

INVx3_ASAP7_75t_L g3393 ( 
.A(n_3082),
.Y(n_3393)
);

HB1xp67_ASAP7_75t_L g3394 ( 
.A(n_3104),
.Y(n_3394)
);

BUFx3_ASAP7_75t_L g3395 ( 
.A(n_2973),
.Y(n_3395)
);

INVx1_ASAP7_75t_SL g3396 ( 
.A(n_3073),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_L g3397 ( 
.A1(n_3111),
.A2(n_3123),
.B1(n_3136),
.B2(n_3267),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3061),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3086),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_2898),
.Y(n_3400)
);

BUFx2_ASAP7_75t_L g3401 ( 
.A(n_3052),
.Y(n_3401)
);

AOI22xp5_ASAP7_75t_L g3402 ( 
.A1(n_2990),
.A2(n_2579),
.B1(n_2572),
.B2(n_2704),
.Y(n_3402)
);

AOI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3111),
.A2(n_3123),
.B1(n_3021),
.B2(n_2936),
.Y(n_3403)
);

CKINVDCx20_ASAP7_75t_R g3404 ( 
.A(n_3069),
.Y(n_3404)
);

AOI22xp33_ASAP7_75t_SL g3405 ( 
.A1(n_3080),
.A2(n_2560),
.B1(n_2580),
.B2(n_2603),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3086),
.Y(n_3406)
);

BUFx4f_ASAP7_75t_L g3407 ( 
.A(n_2923),
.Y(n_3407)
);

OAI22xp5_ASAP7_75t_SL g3408 ( 
.A1(n_3011),
.A2(n_2752),
.B1(n_2740),
.B2(n_2455),
.Y(n_3408)
);

INVx1_ASAP7_75t_SL g3409 ( 
.A(n_2986),
.Y(n_3409)
);

CKINVDCx20_ASAP7_75t_R g3410 ( 
.A(n_2970),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_2938),
.A2(n_2697),
.B1(n_2740),
.B2(n_2773),
.Y(n_3411)
);

OAI22xp33_ASAP7_75t_L g3412 ( 
.A1(n_3227),
.A2(n_2571),
.B1(n_2682),
.B2(n_2702),
.Y(n_3412)
);

AOI22xp33_ASAP7_75t_L g3413 ( 
.A1(n_2951),
.A2(n_2958),
.B1(n_2980),
.B2(n_2955),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2911),
.Y(n_3414)
);

AOI21xp33_ASAP7_75t_L g3415 ( 
.A1(n_3288),
.A2(n_2774),
.B(n_2767),
.Y(n_3415)
);

BUFx12f_ASAP7_75t_L g3416 ( 
.A(n_2882),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_SL g3417 ( 
.A1(n_3080),
.A2(n_2580),
.B1(n_2629),
.B2(n_2603),
.Y(n_3417)
);

AOI22xp33_ASAP7_75t_L g3418 ( 
.A1(n_2985),
.A2(n_2743),
.B1(n_2728),
.B2(n_2557),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2920),
.Y(n_3419)
);

AOI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3199),
.A2(n_2698),
.B1(n_2680),
.B2(n_2742),
.Y(n_3420)
);

AOI22xp33_ASAP7_75t_L g3421 ( 
.A1(n_2940),
.A2(n_2728),
.B1(n_2743),
.B2(n_2553),
.Y(n_3421)
);

INVx3_ASAP7_75t_L g3422 ( 
.A(n_3082),
.Y(n_3422)
);

BUFx2_ASAP7_75t_L g3423 ( 
.A(n_3052),
.Y(n_3423)
);

BUFx3_ASAP7_75t_L g3424 ( 
.A(n_2913),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_SL g3425 ( 
.A1(n_2923),
.A2(n_2629),
.B1(n_2755),
.B2(n_2810),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_2991),
.A2(n_2714),
.B1(n_2723),
.B2(n_2671),
.Y(n_3426)
);

AOI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3250),
.A2(n_3247),
.B1(n_3241),
.B2(n_3312),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3179),
.B(n_2718),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_2881),
.Y(n_3429)
);

OAI21xp33_ASAP7_75t_SL g3430 ( 
.A1(n_3004),
.A2(n_2768),
.B(n_2613),
.Y(n_3430)
);

OAI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_3241),
.A2(n_2713),
.B1(n_2768),
.B2(n_2377),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2892),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3131),
.Y(n_3433)
);

AOI22xp33_ASAP7_75t_SL g3434 ( 
.A1(n_2895),
.A2(n_2828),
.B1(n_2836),
.B2(n_2814),
.Y(n_3434)
);

CKINVDCx6p67_ASAP7_75t_R g3435 ( 
.A(n_3176),
.Y(n_3435)
);

AOI22xp33_ASAP7_75t_L g3436 ( 
.A1(n_3177),
.A2(n_2500),
.B1(n_2526),
.B2(n_2466),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_2929),
.Y(n_3437)
);

CKINVDCx11_ASAP7_75t_R g3438 ( 
.A(n_3031),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3099),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3099),
.Y(n_3440)
);

BUFx6f_ASAP7_75t_L g3441 ( 
.A(n_2881),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3141),
.B(n_2842),
.Y(n_3442)
);

INVx6_ASAP7_75t_L g3443 ( 
.A(n_3172),
.Y(n_3443)
);

AOI22xp5_ASAP7_75t_L g3444 ( 
.A1(n_3198),
.A2(n_2602),
.B1(n_2606),
.B2(n_2397),
.Y(n_3444)
);

BUFx3_ASAP7_75t_L g3445 ( 
.A(n_2908),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3103),
.Y(n_3446)
);

CKINVDCx11_ASAP7_75t_R g3447 ( 
.A(n_2942),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3177),
.A2(n_2324),
.B1(n_2677),
.B2(n_2673),
.Y(n_3448)
);

BUFx3_ASAP7_75t_L g3449 ( 
.A(n_2912),
.Y(n_3449)
);

CKINVDCx11_ASAP7_75t_R g3450 ( 
.A(n_2934),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_2950),
.Y(n_3451)
);

INVx1_ASAP7_75t_SL g3452 ( 
.A(n_3130),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_SL g3453 ( 
.A1(n_2895),
.A2(n_2846),
.B1(n_2734),
.B2(n_2726),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3103),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3084),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3106),
.Y(n_3456)
);

NAND2x1p5_ASAP7_75t_L g3457 ( 
.A(n_3163),
.B(n_2734),
.Y(n_3457)
);

INVx8_ASAP7_75t_L g3458 ( 
.A(n_3026),
.Y(n_3458)
);

INVx1_ASAP7_75t_SL g3459 ( 
.A(n_3211),
.Y(n_3459)
);

BUFx3_ASAP7_75t_L g3460 ( 
.A(n_2971),
.Y(n_3460)
);

BUFx2_ASAP7_75t_L g3461 ( 
.A(n_3209),
.Y(n_3461)
);

CKINVDCx5p33_ASAP7_75t_R g3462 ( 
.A(n_3023),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2965),
.Y(n_3463)
);

OAI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_3213),
.A2(n_2374),
.B1(n_2801),
.B2(n_2798),
.Y(n_3464)
);

INVx6_ASAP7_75t_L g3465 ( 
.A(n_3209),
.Y(n_3465)
);

OAI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3278),
.A2(n_2791),
.B1(n_2327),
.B2(n_2322),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3106),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3107),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3107),
.Y(n_3469)
);

INVx1_ASAP7_75t_SL g3470 ( 
.A(n_2887),
.Y(n_3470)
);

CKINVDCx11_ASAP7_75t_R g3471 ( 
.A(n_2901),
.Y(n_3471)
);

OAI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3278),
.A2(n_2796),
.B1(n_2792),
.B2(n_2452),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_2888),
.B(n_2563),
.Y(n_3473)
);

OAI21xp5_ASAP7_75t_SL g3474 ( 
.A1(n_3144),
.A2(n_2777),
.B(n_2613),
.Y(n_3474)
);

BUFx12f_ASAP7_75t_L g3475 ( 
.A(n_2999),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3185),
.B(n_2566),
.Y(n_3476)
);

BUFx3_ASAP7_75t_L g3477 ( 
.A(n_2921),
.Y(n_3477)
);

BUFx4_ASAP7_75t_R g3478 ( 
.A(n_2967),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_SL g3479 ( 
.A1(n_3026),
.A2(n_2734),
.B1(n_2355),
.B2(n_2787),
.Y(n_3479)
);

INVx6_ASAP7_75t_L g3480 ( 
.A(n_2916),
.Y(n_3480)
);

BUFx4_ASAP7_75t_SL g3481 ( 
.A(n_2922),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_SL g3482 ( 
.A1(n_3279),
.A2(n_2355),
.B1(n_2750),
.B2(n_2736),
.Y(n_3482)
);

CKINVDCx6p67_ASAP7_75t_R g3483 ( 
.A(n_2852),
.Y(n_3483)
);

INVx1_ASAP7_75t_SL g3484 ( 
.A(n_3094),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3146),
.A2(n_2677),
.B1(n_2678),
.B2(n_2673),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3115),
.Y(n_3486)
);

OAI22xp33_ASAP7_75t_L g3487 ( 
.A1(n_3065),
.A2(n_2796),
.B1(n_2792),
.B2(n_2731),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3115),
.Y(n_3488)
);

INVx3_ASAP7_75t_L g3489 ( 
.A(n_3131),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3116),
.Y(n_3490)
);

INVx2_ASAP7_75t_SL g3491 ( 
.A(n_3088),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_2881),
.Y(n_3492)
);

AOI22xp5_ASAP7_75t_SL g3493 ( 
.A1(n_3201),
.A2(n_2331),
.B1(n_2716),
.B2(n_2370),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_2892),
.Y(n_3494)
);

BUFx2_ASAP7_75t_SL g3495 ( 
.A(n_2861),
.Y(n_3495)
);

BUFx10_ASAP7_75t_L g3496 ( 
.A(n_3094),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3245),
.A2(n_2803),
.B1(n_2737),
.B2(n_2739),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_2855),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_2855),
.Y(n_3499)
);

CKINVDCx11_ASAP7_75t_R g3500 ( 
.A(n_2967),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2899),
.Y(n_3501)
);

BUFx2_ASAP7_75t_L g3502 ( 
.A(n_3303),
.Y(n_3502)
);

OAI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3245),
.A2(n_2763),
.B1(n_2765),
.B2(n_2732),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3296),
.A2(n_2690),
.B1(n_2678),
.B2(n_2708),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_L g3505 ( 
.A1(n_3289),
.A2(n_2690),
.B1(n_2720),
.B2(n_2708),
.Y(n_3505)
);

BUFx3_ASAP7_75t_L g3506 ( 
.A(n_2917),
.Y(n_3506)
);

OAI21xp5_ASAP7_75t_SL g3507 ( 
.A1(n_3065),
.A2(n_2589),
.B(n_2520),
.Y(n_3507)
);

BUFx3_ASAP7_75t_L g3508 ( 
.A(n_2928),
.Y(n_3508)
);

BUFx6f_ASAP7_75t_L g3509 ( 
.A(n_2883),
.Y(n_3509)
);

AOI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3142),
.A2(n_2720),
.B1(n_2437),
.B2(n_2330),
.Y(n_3510)
);

AOI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_2868),
.A2(n_2819),
.B1(n_2825),
.B2(n_2813),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_2856),
.Y(n_3512)
);

OAI22xp33_ASAP7_75t_L g3513 ( 
.A1(n_3289),
.A2(n_3309),
.B1(n_3286),
.B2(n_3121),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3294),
.A2(n_2586),
.B1(n_2590),
.B2(n_2587),
.Y(n_3514)
);

INVx6_ASAP7_75t_L g3515 ( 
.A(n_3273),
.Y(n_3515)
);

INVx1_ASAP7_75t_SL g3516 ( 
.A(n_3001),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3294),
.A2(n_2615),
.B1(n_2369),
.B2(n_2619),
.Y(n_3517)
);

BUFx10_ASAP7_75t_L g3518 ( 
.A(n_3242),
.Y(n_3518)
);

AOI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_2987),
.A2(n_2848),
.B1(n_2849),
.B2(n_2843),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3116),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_2856),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3124),
.Y(n_3522)
);

INVx8_ASAP7_75t_L g3523 ( 
.A(n_3311),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_2963),
.Y(n_3524)
);

BUFx2_ASAP7_75t_L g3525 ( 
.A(n_3315),
.Y(n_3525)
);

BUFx3_ASAP7_75t_L g3526 ( 
.A(n_3033),
.Y(n_3526)
);

BUFx4_ASAP7_75t_R g3527 ( 
.A(n_3171),
.Y(n_3527)
);

INVx3_ASAP7_75t_SL g3528 ( 
.A(n_2931),
.Y(n_3528)
);

OAI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_3298),
.A2(n_2778),
.B1(n_2654),
.B2(n_2658),
.Y(n_3529)
);

AOI22xp5_ASAP7_75t_SL g3530 ( 
.A1(n_3184),
.A2(n_3071),
.B1(n_2957),
.B2(n_3092),
.Y(n_3530)
);

INVxp67_ASAP7_75t_SL g3531 ( 
.A(n_3197),
.Y(n_3531)
);

CKINVDCx11_ASAP7_75t_R g3532 ( 
.A(n_2930),
.Y(n_3532)
);

INVxp67_ASAP7_75t_SL g3533 ( 
.A(n_3208),
.Y(n_3533)
);

AOI22xp33_ASAP7_75t_L g3534 ( 
.A1(n_3253),
.A2(n_2640),
.B1(n_2676),
.B2(n_2668),
.Y(n_3534)
);

INVx1_ASAP7_75t_SL g3535 ( 
.A(n_3017),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_2872),
.Y(n_3536)
);

HB1xp67_ASAP7_75t_L g3537 ( 
.A(n_3000),
.Y(n_3537)
);

BUFx8_ASAP7_75t_L g3538 ( 
.A(n_2853),
.Y(n_3538)
);

NAND2x1p5_ASAP7_75t_L g3539 ( 
.A(n_3163),
.B(n_2623),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3124),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3126),
.Y(n_3541)
);

AOI22xp33_ASAP7_75t_SL g3542 ( 
.A1(n_3125),
.A2(n_2716),
.B1(n_2356),
.B2(n_2760),
.Y(n_3542)
);

AOI21xp33_ASAP7_75t_L g3543 ( 
.A1(n_3075),
.A2(n_2542),
.B(n_2536),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3293),
.A2(n_2684),
.B1(n_2692),
.B2(n_2686),
.Y(n_3544)
);

INVx1_ASAP7_75t_SL g3545 ( 
.A(n_2903),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3298),
.A2(n_2727),
.B1(n_2721),
.B2(n_2589),
.Y(n_3546)
);

AOI22xp33_ASAP7_75t_SL g3547 ( 
.A1(n_3125),
.A2(n_2716),
.B1(n_2772),
.B2(n_2760),
.Y(n_3547)
);

INVx4_ASAP7_75t_L g3548 ( 
.A(n_3110),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3185),
.B(n_2616),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3126),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3133),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_2861),
.B(n_2869),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3190),
.A2(n_2546),
.B1(n_2347),
.B2(n_2446),
.Y(n_3553)
);

BUFx3_ASAP7_75t_L g3554 ( 
.A(n_3077),
.Y(n_3554)
);

CKINVDCx11_ASAP7_75t_R g3555 ( 
.A(n_2941),
.Y(n_3555)
);

AOI22xp33_ASAP7_75t_SL g3556 ( 
.A1(n_3159),
.A2(n_2716),
.B1(n_2772),
.B2(n_2760),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_SL g3557 ( 
.A1(n_3159),
.A2(n_2772),
.B1(n_2805),
.B2(n_2416),
.Y(n_3557)
);

INVx3_ASAP7_75t_L g3558 ( 
.A(n_3163),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_2899),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3133),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3137),
.Y(n_3561)
);

INVx1_ASAP7_75t_SL g3562 ( 
.A(n_3078),
.Y(n_3562)
);

CKINVDCx20_ASAP7_75t_R g3563 ( 
.A(n_2996),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_2872),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3193),
.A2(n_2440),
.B1(n_2531),
.B2(n_2467),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3137),
.Y(n_3566)
);

CKINVDCx20_ASAP7_75t_R g3567 ( 
.A(n_3117),
.Y(n_3567)
);

AOI21xp33_ASAP7_75t_L g3568 ( 
.A1(n_3134),
.A2(n_2573),
.B(n_2584),
.Y(n_3568)
);

OAI22xp5_ASAP7_75t_SL g3569 ( 
.A1(n_2919),
.A2(n_2700),
.B1(n_2338),
.B2(n_2343),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_2909),
.Y(n_3570)
);

INVx4_ASAP7_75t_L g3571 ( 
.A(n_2861),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2909),
.Y(n_3572)
);

OAI22x1_ASAP7_75t_L g3573 ( 
.A1(n_3215),
.A2(n_2616),
.B1(n_2426),
.B2(n_2442),
.Y(n_3573)
);

BUFx6f_ASAP7_75t_L g3574 ( 
.A(n_2883),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_2873),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_2873),
.Y(n_3576)
);

INVx2_ASAP7_75t_SL g3577 ( 
.A(n_2954),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_2977),
.Y(n_3578)
);

INVx6_ASAP7_75t_L g3579 ( 
.A(n_2878),
.Y(n_3579)
);

BUFx12f_ASAP7_75t_L g3580 ( 
.A(n_3055),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2925),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_L g3582 ( 
.A1(n_3195),
.A2(n_2344),
.B1(n_2486),
.B2(n_2479),
.Y(n_3582)
);

BUFx12f_ASAP7_75t_L g3583 ( 
.A(n_2949),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_2947),
.A2(n_2524),
.B1(n_2527),
.B2(n_2506),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_2925),
.Y(n_3585)
);

AOI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_2948),
.A2(n_2416),
.B1(n_2442),
.B2(n_2426),
.Y(n_3586)
);

INVx2_ASAP7_75t_SL g3587 ( 
.A(n_3076),
.Y(n_3587)
);

AOI22xp33_ASAP7_75t_L g3588 ( 
.A1(n_3147),
.A2(n_2453),
.B1(n_2335),
.B2(n_2382),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_2935),
.Y(n_3589)
);

CKINVDCx6p67_ASAP7_75t_R g3590 ( 
.A(n_2869),
.Y(n_3590)
);

INVx6_ASAP7_75t_L g3591 ( 
.A(n_2878),
.Y(n_3591)
);

AOI22xp33_ASAP7_75t_SL g3592 ( 
.A1(n_3188),
.A2(n_2453),
.B1(n_2834),
.B2(n_2634),
.Y(n_3592)
);

OAI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3121),
.A2(n_2385),
.B1(n_2390),
.B2(n_2386),
.Y(n_3593)
);

AOI22xp33_ASAP7_75t_L g3594 ( 
.A1(n_3170),
.A2(n_3188),
.B1(n_3022),
.B2(n_3284),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3191),
.B(n_2634),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3015),
.A2(n_2403),
.B1(n_2402),
.B2(n_2548),
.Y(n_3596)
);

OAI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3019),
.A2(n_2554),
.B1(n_2665),
.B2(n_2661),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2935),
.Y(n_3598)
);

INVxp67_ASAP7_75t_SL g3599 ( 
.A(n_3212),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_2937),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_2937),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_2946),
.Y(n_3602)
);

CKINVDCx11_ASAP7_75t_R g3603 ( 
.A(n_3037),
.Y(n_3603)
);

INVx6_ASAP7_75t_L g3604 ( 
.A(n_2915),
.Y(n_3604)
);

OAI22xp5_ASAP7_75t_L g3605 ( 
.A1(n_2865),
.A2(n_2661),
.B1(n_2665),
.B2(n_2599),
.Y(n_3605)
);

BUFx12f_ASAP7_75t_L g3606 ( 
.A(n_2915),
.Y(n_3606)
);

INVxp67_ASAP7_75t_L g3607 ( 
.A(n_2886),
.Y(n_3607)
);

INVx4_ASAP7_75t_L g3608 ( 
.A(n_2869),
.Y(n_3608)
);

AOI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3299),
.A2(n_2659),
.B1(n_2660),
.B2(n_2786),
.Y(n_3609)
);

INVx6_ASAP7_75t_L g3610 ( 
.A(n_3284),
.Y(n_3610)
);

BUFx2_ASAP7_75t_L g3611 ( 
.A(n_2863),
.Y(n_3611)
);

CKINVDCx20_ASAP7_75t_R g3612 ( 
.A(n_3266),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_2997),
.Y(n_3613)
);

BUFx3_ASAP7_75t_L g3614 ( 
.A(n_3089),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_SL g3615 ( 
.A1(n_2989),
.A2(n_2834),
.B1(n_2623),
.B2(n_2719),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_2946),
.Y(n_3616)
);

OAI22xp5_ASAP7_75t_L g3617 ( 
.A1(n_2865),
.A2(n_2659),
.B1(n_2794),
.B2(n_2793),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_2883),
.Y(n_3618)
);

AOI22xp33_ASAP7_75t_SL g3619 ( 
.A1(n_3014),
.A2(n_2834),
.B1(n_2719),
.B2(n_2701),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3280),
.B(n_2664),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_2959),
.Y(n_3621)
);

BUFx10_ASAP7_75t_L g3622 ( 
.A(n_3242),
.Y(n_3622)
);

OAI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_2894),
.A2(n_2660),
.B1(n_2611),
.B2(n_2396),
.Y(n_3623)
);

INVx6_ASAP7_75t_L g3624 ( 
.A(n_3101),
.Y(n_3624)
);

BUFx3_ASAP7_75t_L g3625 ( 
.A(n_3072),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3161),
.A2(n_2802),
.B1(n_2786),
.B2(n_2699),
.Y(n_3626)
);

AOI22xp33_ASAP7_75t_L g3627 ( 
.A1(n_3161),
.A2(n_2802),
.B1(n_2695),
.B2(n_2396),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_2959),
.Y(n_3628)
);

INVx6_ASAP7_75t_L g3629 ( 
.A(n_3183),
.Y(n_3629)
);

CKINVDCx20_ASAP7_75t_R g3630 ( 
.A(n_3248),
.Y(n_3630)
);

AOI22xp33_ASAP7_75t_L g3631 ( 
.A1(n_3219),
.A2(n_2401),
.B1(n_2451),
.B2(n_2365),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3219),
.A2(n_2401),
.B1(n_2451),
.B2(n_2365),
.Y(n_3632)
);

BUFx4_ASAP7_75t_SL g3633 ( 
.A(n_3109),
.Y(n_3633)
);

OR2x2_ASAP7_75t_L g3634 ( 
.A(n_3000),
.B(n_2552),
.Y(n_3634)
);

CKINVDCx16_ASAP7_75t_R g3635 ( 
.A(n_2897),
.Y(n_3635)
);

AOI22xp33_ASAP7_75t_L g3636 ( 
.A1(n_3229),
.A2(n_2807),
.B1(n_2749),
.B2(n_2552),
.Y(n_3636)
);

BUFx3_ASAP7_75t_L g3637 ( 
.A(n_3053),
.Y(n_3637)
);

INVxp67_ASAP7_75t_SL g3638 ( 
.A(n_3235),
.Y(n_3638)
);

CKINVDCx20_ASAP7_75t_R g3639 ( 
.A(n_2918),
.Y(n_3639)
);

AOI22xp5_ASAP7_75t_L g3640 ( 
.A1(n_3320),
.A2(n_2596),
.B1(n_2594),
.B2(n_2749),
.Y(n_3640)
);

BUFx8_ASAP7_75t_SL g3641 ( 
.A(n_3182),
.Y(n_3641)
);

CKINVDCx11_ASAP7_75t_R g3642 ( 
.A(n_3230),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_L g3643 ( 
.A1(n_3229),
.A2(n_2596),
.B1(n_2535),
.B2(n_2513),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3308),
.A2(n_2535),
.B1(n_2513),
.B2(n_2753),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_SL g3645 ( 
.A1(n_3204),
.A2(n_2834),
.B1(n_2719),
.B2(n_2701),
.Y(n_3645)
);

BUFx6f_ASAP7_75t_SL g3646 ( 
.A(n_3242),
.Y(n_3646)
);

BUFx12f_ASAP7_75t_L g3647 ( 
.A(n_2926),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3308),
.A2(n_2753),
.B1(n_2834),
.B2(n_2806),
.Y(n_3648)
);

BUFx10_ASAP7_75t_L g3649 ( 
.A(n_3242),
.Y(n_3649)
);

AOI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3063),
.A2(n_2379),
.B1(n_2753),
.B2(n_2471),
.Y(n_3650)
);

INVx3_ASAP7_75t_L g3651 ( 
.A(n_2894),
.Y(n_3651)
);

BUFx3_ASAP7_75t_L g3652 ( 
.A(n_3118),
.Y(n_3652)
);

AOI22xp33_ASAP7_75t_SL g3653 ( 
.A1(n_3216),
.A2(n_2701),
.B1(n_2469),
.B2(n_2484),
.Y(n_3653)
);

AOI22xp5_ASAP7_75t_SL g3654 ( 
.A1(n_3051),
.A2(n_2469),
.B1(n_2471),
.B2(n_2484),
.Y(n_3654)
);

BUFx8_ASAP7_75t_L g3655 ( 
.A(n_2998),
.Y(n_3655)
);

INVx2_ASAP7_75t_SL g3656 ( 
.A(n_2966),
.Y(n_3656)
);

AOI22xp33_ASAP7_75t_L g3657 ( 
.A1(n_3310),
.A2(n_2806),
.B1(n_2445),
.B2(n_2488),
.Y(n_3657)
);

OAI22xp5_ASAP7_75t_SL g3658 ( 
.A1(n_3098),
.A2(n_2540),
.B1(n_2559),
.B2(n_2550),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3009),
.Y(n_3659)
);

AOI22xp33_ASAP7_75t_SL g3660 ( 
.A1(n_3224),
.A2(n_2488),
.B1(n_2492),
.B2(n_2540),
.Y(n_3660)
);

AO22x1_ASAP7_75t_L g3661 ( 
.A1(n_2894),
.A2(n_2492),
.B1(n_2550),
.B2(n_2540),
.Y(n_3661)
);

INVx3_ASAP7_75t_L g3662 ( 
.A(n_2902),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_2972),
.Y(n_3663)
);

OAI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_2902),
.A2(n_2960),
.B1(n_2939),
.B2(n_3292),
.Y(n_3664)
);

CKINVDCx6p67_ASAP7_75t_R g3665 ( 
.A(n_2902),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3034),
.Y(n_3666)
);

OAI22xp33_ASAP7_75t_L g3667 ( 
.A1(n_3281),
.A2(n_2806),
.B1(n_2492),
.B2(n_2544),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_2988),
.B(n_242),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3056),
.Y(n_3669)
);

BUFx3_ASAP7_75t_L g3670 ( 
.A(n_3119),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3074),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_2972),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_2974),
.Y(n_3673)
);

CKINVDCx6p67_ASAP7_75t_R g3674 ( 
.A(n_2939),
.Y(n_3674)
);

CKINVDCx11_ASAP7_75t_R g3675 ( 
.A(n_3230),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3085),
.Y(n_3676)
);

CKINVDCx11_ASAP7_75t_R g3677 ( 
.A(n_3068),
.Y(n_3677)
);

AOI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3139),
.A2(n_2559),
.B1(n_2569),
.B2(n_2550),
.Y(n_3678)
);

BUFx8_ASAP7_75t_SL g3679 ( 
.A(n_3323),
.Y(n_3679)
);

BUFx12f_ASAP7_75t_L g3680 ( 
.A(n_3167),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_SL g3681 ( 
.A1(n_2939),
.A2(n_2569),
.B1(n_2593),
.B2(n_2559),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_2974),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3002),
.Y(n_3683)
);

INVx6_ASAP7_75t_L g3684 ( 
.A(n_3167),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3002),
.Y(n_3685)
);

BUFx12f_ASAP7_75t_L g3686 ( 
.A(n_3007),
.Y(n_3686)
);

AOI22xp33_ASAP7_75t_L g3687 ( 
.A1(n_3249),
.A2(n_2804),
.B1(n_2593),
.B2(n_2635),
.Y(n_3687)
);

INVx6_ASAP7_75t_L g3688 ( 
.A(n_2960),
.Y(n_3688)
);

INVx6_ASAP7_75t_L g3689 ( 
.A(n_2960),
.Y(n_3689)
);

INVxp67_ASAP7_75t_L g3690 ( 
.A(n_3097),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3096),
.Y(n_3691)
);

BUFx12f_ASAP7_75t_L g3692 ( 
.A(n_3018),
.Y(n_3692)
);

CKINVDCx20_ASAP7_75t_R g3693 ( 
.A(n_3102),
.Y(n_3693)
);

AOI22xp33_ASAP7_75t_L g3694 ( 
.A1(n_3114),
.A2(n_2804),
.B1(n_2593),
.B2(n_2635),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3148),
.Y(n_3695)
);

CKINVDCx5p33_ASAP7_75t_R g3696 ( 
.A(n_3166),
.Y(n_3696)
);

OAI21xp5_ASAP7_75t_SL g3697 ( 
.A1(n_3281),
.A2(n_2635),
.B(n_2569),
.Y(n_3697)
);

BUFx2_ASAP7_75t_L g3698 ( 
.A(n_2885),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3108),
.Y(n_3699)
);

INVx3_ASAP7_75t_L g3700 ( 
.A(n_2982),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3148),
.Y(n_3701)
);

BUFx2_ASAP7_75t_SL g3702 ( 
.A(n_3024),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3120),
.A2(n_2804),
.B1(n_2649),
.B2(n_246),
.Y(n_3703)
);

BUFx3_ASAP7_75t_L g3704 ( 
.A(n_3128),
.Y(n_3704)
);

BUFx8_ASAP7_75t_L g3705 ( 
.A(n_3016),
.Y(n_3705)
);

INVx6_ASAP7_75t_L g3706 ( 
.A(n_3206),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_L g3707 ( 
.A1(n_3062),
.A2(n_2649),
.B1(n_247),
.B2(n_244),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3154),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_SL g3709 ( 
.A1(n_2932),
.A2(n_2649),
.B1(n_247),
.B2(n_244),
.Y(n_3709)
);

AOI22xp33_ASAP7_75t_L g3710 ( 
.A1(n_3262),
.A2(n_249),
.B1(n_245),
.B2(n_248),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3154),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3191),
.B(n_245),
.Y(n_3712)
);

AOI22xp33_ASAP7_75t_L g3713 ( 
.A1(n_3081),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3162),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3162),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3168),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3083),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3168),
.Y(n_3718)
);

OAI22xp33_ASAP7_75t_L g3719 ( 
.A1(n_3006),
.A2(n_255),
.B1(n_252),
.B2(n_253),
.Y(n_3719)
);

CKINVDCx6p67_ASAP7_75t_R g3720 ( 
.A(n_3024),
.Y(n_3720)
);

INVx6_ASAP7_75t_L g3721 ( 
.A(n_3206),
.Y(n_3721)
);

BUFx4f_ASAP7_75t_SL g3722 ( 
.A(n_3202),
.Y(n_3722)
);

OAI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_2875),
.A2(n_253),
.B(n_255),
.Y(n_3723)
);

CKINVDCx11_ASAP7_75t_R g3724 ( 
.A(n_2961),
.Y(n_3724)
);

OAI22xp5_ASAP7_75t_SL g3725 ( 
.A1(n_2976),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_3725)
);

AOI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_3388),
.A2(n_2993),
.B1(n_2860),
.B2(n_3205),
.Y(n_3726)
);

AOI22xp33_ASAP7_75t_L g3727 ( 
.A1(n_3342),
.A2(n_3349),
.B1(n_3324),
.B2(n_3370),
.Y(n_3727)
);

BUFx3_ASAP7_75t_L g3728 ( 
.A(n_3630),
.Y(n_3728)
);

NAND3xp33_ASAP7_75t_L g3729 ( 
.A(n_3482),
.B(n_3418),
.C(n_3381),
.Y(n_3729)
);

AOI22xp33_ASAP7_75t_L g3730 ( 
.A1(n_3385),
.A2(n_3158),
.B1(n_3302),
.B2(n_3220),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_SL g3731 ( 
.A1(n_3347),
.A2(n_3143),
.B1(n_3024),
.B2(n_3028),
.Y(n_3731)
);

AOI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3347),
.A2(n_3231),
.B1(n_3194),
.B2(n_2880),
.Y(n_3732)
);

OAI21xp5_ASAP7_75t_SL g3733 ( 
.A1(n_3336),
.A2(n_3054),
.B(n_3035),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3329),
.Y(n_3734)
);

BUFx12f_ASAP7_75t_L g3735 ( 
.A(n_3332),
.Y(n_3735)
);

OAI22xp5_ASAP7_75t_L g3736 ( 
.A1(n_3339),
.A2(n_3143),
.B1(n_3207),
.B2(n_3006),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3374),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3329),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3330),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3330),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3369),
.B(n_3044),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3432),
.Y(n_3742)
);

INVx4_ASAP7_75t_L g3743 ( 
.A(n_3527),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_L g3744 ( 
.A1(n_3347),
.A2(n_2880),
.B1(n_2871),
.B2(n_3044),
.Y(n_3744)
);

INVx3_ASAP7_75t_L g3745 ( 
.A(n_3518),
.Y(n_3745)
);

AOI22xp33_ASAP7_75t_L g3746 ( 
.A1(n_3472),
.A2(n_2880),
.B1(n_2871),
.B2(n_3046),
.Y(n_3746)
);

OAI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3384),
.A2(n_3238),
.B(n_3180),
.Y(n_3747)
);

OAI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3405),
.A2(n_3143),
.B1(n_3046),
.B2(n_3093),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3387),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3466),
.A2(n_2880),
.B1(n_2871),
.B2(n_3192),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3376),
.A2(n_2880),
.B1(n_2871),
.B2(n_3232),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3442),
.B(n_3620),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3432),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3343),
.B(n_3196),
.Y(n_3754)
);

HB1xp67_ASAP7_75t_L g3755 ( 
.A(n_3394),
.Y(n_3755)
);

AOI222xp33_ASAP7_75t_L g3756 ( 
.A1(n_3513),
.A2(n_3040),
.B1(n_3045),
.B2(n_2995),
.C1(n_3039),
.C2(n_3196),
.Y(n_3756)
);

AOI22xp33_ASAP7_75t_L g3757 ( 
.A1(n_3464),
.A2(n_2871),
.B1(n_3221),
.B2(n_3218),
.Y(n_3757)
);

OAI21xp33_ASAP7_75t_L g3758 ( 
.A1(n_3542),
.A2(n_3260),
.B(n_3058),
.Y(n_3758)
);

AND2x2_ASAP7_75t_SL g3759 ( 
.A(n_3407),
.B(n_3237),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3355),
.B(n_3218),
.Y(n_3760)
);

AOI22xp33_ASAP7_75t_L g3761 ( 
.A1(n_3569),
.A2(n_3236),
.B1(n_3258),
.B2(n_3221),
.Y(n_3761)
);

OAI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3417),
.A2(n_3020),
.B1(n_3048),
.B2(n_3290),
.Y(n_3762)
);

BUFx5_ASAP7_75t_L g3763 ( 
.A(n_3518),
.Y(n_3763)
);

INVx5_ASAP7_75t_SL g3764 ( 
.A(n_3435),
.Y(n_3764)
);

INVx3_ASAP7_75t_L g3765 ( 
.A(n_3622),
.Y(n_3765)
);

AOI22xp33_ASAP7_75t_SL g3766 ( 
.A1(n_3646),
.A2(n_2982),
.B1(n_3042),
.B2(n_3041),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3358),
.B(n_3236),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3357),
.A2(n_3048),
.B1(n_3319),
.B2(n_3317),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3375),
.A2(n_3258),
.B1(n_3265),
.B2(n_3264),
.Y(n_3769)
);

OAI21xp5_ASAP7_75t_SL g3770 ( 
.A1(n_3474),
.A2(n_3100),
.B(n_3095),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3362),
.B(n_3264),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3494),
.Y(n_3772)
);

AOI22xp33_ASAP7_75t_L g3773 ( 
.A1(n_3593),
.A2(n_3265),
.B1(n_3272),
.B2(n_3271),
.Y(n_3773)
);

BUFx4f_ASAP7_75t_SL g3774 ( 
.A(n_3328),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3494),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3473),
.B(n_3149),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3366),
.B(n_3271),
.Y(n_3777)
);

OAI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3402),
.A2(n_3239),
.B1(n_3275),
.B2(n_2914),
.Y(n_3778)
);

OAI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3346),
.A2(n_3338),
.B1(n_3547),
.B2(n_3421),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3408),
.A2(n_3348),
.B1(n_3487),
.B2(n_3390),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3501),
.Y(n_3781)
);

AOI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_3725),
.A2(n_3272),
.B1(n_3317),
.B2(n_3297),
.Y(n_3782)
);

INVx1_ASAP7_75t_SL g3783 ( 
.A(n_3603),
.Y(n_3783)
);

OAI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_3722),
.A2(n_2914),
.B1(n_3319),
.B2(n_3297),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3501),
.Y(n_3785)
);

INVx1_ASAP7_75t_SL g3786 ( 
.A(n_3641),
.Y(n_3786)
);

AOI22xp33_ASAP7_75t_L g3787 ( 
.A1(n_3425),
.A2(n_3321),
.B1(n_3322),
.B2(n_3153),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3559),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3559),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3683),
.Y(n_3790)
);

INVx1_ASAP7_75t_SL g3791 ( 
.A(n_3679),
.Y(n_3791)
);

BUFx2_ASAP7_75t_L g3792 ( 
.A(n_3506),
.Y(n_3792)
);

AOI222xp33_ASAP7_75t_L g3793 ( 
.A1(n_3647),
.A2(n_3321),
.B1(n_3322),
.B2(n_3135),
.C1(n_3164),
.C2(n_3140),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3683),
.Y(n_3794)
);

INVx3_ASAP7_75t_L g3795 ( 
.A(n_3622),
.Y(n_3795)
);

OAI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3693),
.A2(n_3244),
.B1(n_3202),
.B2(n_2907),
.Y(n_3796)
);

BUFx4f_ASAP7_75t_SL g3797 ( 
.A(n_3567),
.Y(n_3797)
);

AOI22xp33_ASAP7_75t_L g3798 ( 
.A1(n_3646),
.A2(n_2952),
.B1(n_3038),
.B2(n_2906),
.Y(n_3798)
);

BUFx2_ASAP7_75t_L g3799 ( 
.A(n_3356),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3411),
.A2(n_3122),
.B1(n_3178),
.B2(n_2905),
.Y(n_3800)
);

OAI21xp33_ASAP7_75t_L g3801 ( 
.A1(n_3582),
.A2(n_3032),
.B(n_2879),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3596),
.A2(n_2893),
.B1(n_2889),
.B2(n_3244),
.Y(n_3802)
);

OAI22xp5_ASAP7_75t_L g3803 ( 
.A1(n_3505),
.A2(n_3042),
.B1(n_3087),
.B2(n_3041),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3382),
.B(n_3112),
.Y(n_3804)
);

CKINVDCx5p33_ASAP7_75t_R g3805 ( 
.A(n_3354),
.Y(n_3805)
);

BUFx6f_ASAP7_75t_L g3806 ( 
.A(n_3383),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3685),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3398),
.B(n_3113),
.Y(n_3808)
);

AOI22xp33_ASAP7_75t_L g3809 ( 
.A1(n_3497),
.A2(n_3431),
.B1(n_3568),
.B2(n_3352),
.Y(n_3809)
);

BUFx2_ASAP7_75t_L g3810 ( 
.A(n_3356),
.Y(n_3810)
);

OAI22xp5_ASAP7_75t_L g3811 ( 
.A1(n_3485),
.A2(n_3087),
.B1(n_3100),
.B2(n_3095),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3334),
.A2(n_3150),
.B1(n_3105),
.B2(n_2893),
.Y(n_3812)
);

AOI22xp33_ASAP7_75t_L g3813 ( 
.A1(n_3543),
.A2(n_2889),
.B1(n_3145),
.B2(n_3132),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3668),
.B(n_3160),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3685),
.Y(n_3815)
);

INVx4_ASAP7_75t_SL g3816 ( 
.A(n_3380),
.Y(n_3816)
);

BUFx4f_ASAP7_75t_SL g3817 ( 
.A(n_3563),
.Y(n_3817)
);

AOI22xp33_ASAP7_75t_L g3818 ( 
.A1(n_3686),
.A2(n_3692),
.B1(n_3415),
.B2(n_3586),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_SL g3819 ( 
.A1(n_3493),
.A2(n_3150),
.B1(n_3105),
.B2(n_3200),
.Y(n_3819)
);

AOI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3529),
.A2(n_3155),
.B1(n_3156),
.B2(n_3151),
.Y(n_3820)
);

NOR2xp33_ASAP7_75t_L g3821 ( 
.A(n_3452),
.B(n_3255),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_L g3822 ( 
.A1(n_3553),
.A2(n_3222),
.B1(n_3228),
.B2(n_3186),
.Y(n_3822)
);

OAI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3426),
.A2(n_2981),
.B1(n_2968),
.B2(n_3246),
.Y(n_3823)
);

INVxp67_ASAP7_75t_L g3824 ( 
.A(n_3379),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3399),
.B(n_3254),
.Y(n_3825)
);

AOI22xp33_ASAP7_75t_SL g3826 ( 
.A1(n_3649),
.A2(n_3252),
.B1(n_2981),
.B2(n_2968),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3565),
.A2(n_3259),
.B1(n_3277),
.B2(n_3261),
.Y(n_3827)
);

AOI222xp33_ASAP7_75t_L g3828 ( 
.A1(n_3407),
.A2(n_3461),
.B1(n_3723),
.B2(n_3367),
.C1(n_3345),
.C2(n_3465),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3406),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3439),
.Y(n_3830)
);

OAI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3511),
.A2(n_3287),
.B(n_3285),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_L g3832 ( 
.A1(n_3412),
.A2(n_3263),
.B1(n_3274),
.B2(n_3256),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3440),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3446),
.B(n_3157),
.Y(n_3834)
);

BUFx12f_ASAP7_75t_L g3835 ( 
.A(n_3438),
.Y(n_3835)
);

BUFx2_ASAP7_75t_L g3836 ( 
.A(n_3383),
.Y(n_3836)
);

OAI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3434),
.A2(n_3504),
.B1(n_3448),
.B2(n_3510),
.Y(n_3837)
);

BUFx12f_ASAP7_75t_L g3838 ( 
.A(n_3335),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3503),
.A2(n_3282),
.B1(n_3295),
.B2(n_3276),
.Y(n_3839)
);

OAI22xp5_ASAP7_75t_L g3840 ( 
.A1(n_3436),
.A2(n_3210),
.B1(n_3217),
.B2(n_3206),
.Y(n_3840)
);

AOI22xp33_ASAP7_75t_L g3841 ( 
.A1(n_3588),
.A2(n_3057),
.B1(n_3233),
.B2(n_3050),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3454),
.B(n_3157),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3584),
.A2(n_3057),
.B1(n_3233),
.B2(n_3050),
.Y(n_3843)
);

BUFx6f_ASAP7_75t_L g3844 ( 
.A(n_3383),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3594),
.A2(n_3057),
.B1(n_3233),
.B2(n_3050),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3524),
.Y(n_3846)
);

BUFx4f_ASAP7_75t_SL g3847 ( 
.A(n_3680),
.Y(n_3847)
);

AOI22xp33_ASAP7_75t_SL g3848 ( 
.A1(n_3649),
.A2(n_3057),
.B1(n_3233),
.B2(n_3050),
.Y(n_3848)
);

OAI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3368),
.A2(n_3217),
.B1(n_3225),
.B2(n_3210),
.Y(n_3849)
);

AOI22xp33_ASAP7_75t_L g3850 ( 
.A1(n_3534),
.A2(n_3057),
.B1(n_3233),
.B2(n_3050),
.Y(n_3850)
);

OAI21xp5_ASAP7_75t_SL g3851 ( 
.A1(n_3397),
.A2(n_3257),
.B(n_3234),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3544),
.A2(n_3181),
.B1(n_3189),
.B2(n_3187),
.Y(n_3852)
);

OAI22xp33_ASAP7_75t_L g3853 ( 
.A1(n_3371),
.A2(n_3316),
.B1(n_3169),
.B2(n_3225),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3400),
.Y(n_3854)
);

AND2x6_ASAP7_75t_L g3855 ( 
.A(n_3651),
.B(n_3234),
.Y(n_3855)
);

AOI22xp33_ASAP7_75t_L g3856 ( 
.A1(n_3597),
.A2(n_3181),
.B1(n_3189),
.B2(n_3187),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_L g3857 ( 
.A1(n_3626),
.A2(n_3210),
.B1(n_3225),
.B2(n_3217),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3537),
.B(n_256),
.Y(n_3858)
);

OAI22xp5_ASAP7_75t_L g3859 ( 
.A1(n_3627),
.A2(n_3269),
.B1(n_3305),
.B2(n_3304),
.Y(n_3859)
);

BUFx2_ASAP7_75t_L g3860 ( 
.A(n_3395),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_L g3861 ( 
.A1(n_3517),
.A2(n_3214),
.B1(n_3223),
.B2(n_3169),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_3690),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3456),
.B(n_3467),
.Y(n_3863)
);

AOI22xp33_ASAP7_75t_SL g3864 ( 
.A1(n_3698),
.A2(n_3316),
.B1(n_3214),
.B2(n_3223),
.Y(n_3864)
);

INVx2_ASAP7_75t_SL g3865 ( 
.A(n_3380),
.Y(n_3865)
);

AOI22xp33_ASAP7_75t_L g3866 ( 
.A1(n_3709),
.A2(n_3268),
.B1(n_3270),
.B2(n_3257),
.Y(n_3866)
);

OAI21xp5_ASAP7_75t_SL g3867 ( 
.A1(n_3697),
.A2(n_3270),
.B(n_3268),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3414),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3468),
.Y(n_3869)
);

OAI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_3631),
.A2(n_3304),
.B1(n_3305),
.B2(n_3269),
.Y(n_3870)
);

INVx3_ASAP7_75t_L g3871 ( 
.A(n_3571),
.Y(n_3871)
);

AOI22xp33_ASAP7_75t_L g3872 ( 
.A1(n_3677),
.A2(n_3306),
.B1(n_3304),
.B2(n_3305),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3419),
.Y(n_3873)
);

AOI22xp33_ASAP7_75t_L g3874 ( 
.A1(n_3514),
.A2(n_3306),
.B1(n_3307),
.B2(n_3269),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3652),
.B(n_257),
.Y(n_3875)
);

OAI22xp5_ASAP7_75t_L g3876 ( 
.A1(n_3632),
.A2(n_3307),
.B1(n_3127),
.B2(n_3138),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3724),
.A2(n_3307),
.B1(n_2945),
.B2(n_2962),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3469),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3486),
.Y(n_3879)
);

OAI21xp5_ASAP7_75t_SL g3880 ( 
.A1(n_3378),
.A2(n_2945),
.B(n_2943),
.Y(n_3880)
);

OAI222xp33_ASAP7_75t_L g3881 ( 
.A1(n_3479),
.A2(n_260),
.B1(n_262),
.B2(n_258),
.C1(n_259),
.C2(n_261),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_3393),
.B(n_2943),
.Y(n_3882)
);

NOR2xp33_ASAP7_75t_L g3883 ( 
.A(n_3516),
.B(n_259),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3670),
.B(n_261),
.Y(n_3884)
);

AOI22xp5_ASAP7_75t_L g3885 ( 
.A1(n_3420),
.A2(n_2945),
.B1(n_2962),
.B2(n_2943),
.Y(n_3885)
);

AOI22xp5_ASAP7_75t_SL g3886 ( 
.A1(n_3364),
.A2(n_2979),
.B1(n_2983),
.B2(n_2962),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_L g3887 ( 
.A1(n_3710),
.A2(n_2983),
.B1(n_2994),
.B2(n_2979),
.Y(n_3887)
);

OAI22xp5_ASAP7_75t_L g3888 ( 
.A1(n_3333),
.A2(n_3283),
.B1(n_3301),
.B2(n_3243),
.Y(n_3888)
);

INVx3_ASAP7_75t_SL g3889 ( 
.A(n_3515),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3488),
.Y(n_3890)
);

AOI222xp33_ASAP7_75t_L g3891 ( 
.A1(n_3465),
.A2(n_265),
.B1(n_268),
.B2(n_262),
.C1(n_263),
.C2(n_266),
.Y(n_3891)
);

BUFx4f_ASAP7_75t_SL g3892 ( 
.A(n_3359),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_SL g3893 ( 
.A1(n_3371),
.A2(n_2983),
.B1(n_2994),
.B2(n_2979),
.Y(n_3893)
);

CKINVDCx6p67_ASAP7_75t_R g3894 ( 
.A(n_3371),
.Y(n_3894)
);

AOI22xp5_ASAP7_75t_L g3895 ( 
.A1(n_3444),
.A2(n_3005),
.B1(n_3008),
.B2(n_2994),
.Y(n_3895)
);

BUFx6f_ASAP7_75t_L g3896 ( 
.A(n_3429),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3490),
.Y(n_3897)
);

NOR2x1_ASAP7_75t_L g3898 ( 
.A(n_3393),
.B(n_3005),
.Y(n_3898)
);

OAI21xp5_ASAP7_75t_SL g3899 ( 
.A1(n_3507),
.A2(n_3008),
.B(n_3005),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_L g3900 ( 
.A1(n_3705),
.A2(n_3030),
.B1(n_3036),
.B2(n_3008),
.Y(n_3900)
);

OAI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_3609),
.A2(n_3090),
.B1(n_3091),
.B2(n_3079),
.Y(n_3901)
);

BUFx5_ASAP7_75t_L g3902 ( 
.A(n_3695),
.Y(n_3902)
);

BUFx2_ASAP7_75t_L g3903 ( 
.A(n_3422),
.Y(n_3903)
);

OAI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3377),
.A2(n_3090),
.B1(n_3091),
.B2(n_3079),
.Y(n_3904)
);

CKINVDCx5p33_ASAP7_75t_R g3905 ( 
.A(n_3481),
.Y(n_3905)
);

AOI22xp33_ASAP7_75t_SL g3906 ( 
.A1(n_3495),
.A2(n_3036),
.B1(n_3043),
.B2(n_3030),
.Y(n_3906)
);

BUFx4f_ASAP7_75t_SL g3907 ( 
.A(n_3373),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3705),
.A2(n_3036),
.B1(n_3043),
.B2(n_3030),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3519),
.A2(n_3047),
.B1(n_3060),
.B2(n_3043),
.Y(n_3909)
);

AOI22xp33_ASAP7_75t_L g3910 ( 
.A1(n_3546),
.A2(n_3060),
.B1(n_3064),
.B2(n_3047),
.Y(n_3910)
);

AOI22xp33_ASAP7_75t_L g3911 ( 
.A1(n_3351),
.A2(n_3060),
.B1(n_3064),
.B2(n_3047),
.Y(n_3911)
);

INVx1_ASAP7_75t_SL g3912 ( 
.A(n_3562),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3437),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3520),
.B(n_3064),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3522),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3540),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3451),
.Y(n_3917)
);

NOR2xp33_ASAP7_75t_L g3918 ( 
.A(n_3535),
.B(n_3459),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3607),
.Y(n_3919)
);

CKINVDCx5p33_ASAP7_75t_R g3920 ( 
.A(n_3341),
.Y(n_3920)
);

AOI22xp33_ASAP7_75t_L g3921 ( 
.A1(n_3351),
.A2(n_3079),
.B1(n_3090),
.B2(n_3066),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3541),
.Y(n_3922)
);

HB1xp67_ASAP7_75t_L g3923 ( 
.A(n_3634),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3463),
.Y(n_3924)
);

BUFx6f_ASAP7_75t_L g3925 ( 
.A(n_3429),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3422),
.Y(n_3926)
);

BUFx4f_ASAP7_75t_SL g3927 ( 
.A(n_3612),
.Y(n_3927)
);

AOI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3719),
.A2(n_3091),
.B1(n_3127),
.B2(n_3066),
.Y(n_3928)
);

AOI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3707),
.A2(n_3127),
.B1(n_3138),
.B2(n_3066),
.Y(n_3929)
);

BUFx12f_ASAP7_75t_L g3930 ( 
.A(n_3340),
.Y(n_3930)
);

AOI22xp33_ASAP7_75t_L g3931 ( 
.A1(n_3617),
.A2(n_3152),
.B1(n_3165),
.B2(n_3138),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3550),
.Y(n_3932)
);

INVx4_ASAP7_75t_SL g3933 ( 
.A(n_3443),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3551),
.Y(n_3934)
);

BUFx2_ASAP7_75t_L g3935 ( 
.A(n_3433),
.Y(n_3935)
);

OAI222xp33_ASAP7_75t_L g3936 ( 
.A1(n_3557),
.A2(n_268),
.B1(n_270),
.B2(n_265),
.C1(n_266),
.C2(n_269),
.Y(n_3936)
);

BUFx4f_ASAP7_75t_SL g3937 ( 
.A(n_3386),
.Y(n_3937)
);

BUFx6f_ASAP7_75t_L g3938 ( 
.A(n_3429),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3430),
.A2(n_3165),
.B(n_3152),
.Y(n_3939)
);

AND2x4_ASAP7_75t_L g3940 ( 
.A(n_3695),
.B(n_3152),
.Y(n_3940)
);

OAI21xp33_ASAP7_75t_SL g3941 ( 
.A1(n_3552),
.A2(n_3489),
.B(n_3433),
.Y(n_3941)
);

INVx2_ASAP7_75t_SL g3942 ( 
.A(n_3443),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3560),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3561),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3325),
.Y(n_3945)
);

BUFx6f_ASAP7_75t_L g3946 ( 
.A(n_3441),
.Y(n_3946)
);

AOI22xp33_ASAP7_75t_L g3947 ( 
.A1(n_3392),
.A2(n_3174),
.B1(n_3226),
.B2(n_3165),
.Y(n_3947)
);

NOR2xp33_ASAP7_75t_L g3948 ( 
.A(n_3635),
.B(n_839),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3701),
.A2(n_3226),
.B1(n_3243),
.B2(n_3174),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3566),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3344),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3570),
.B(n_3174),
.Y(n_3952)
);

OAI22xp5_ASAP7_75t_L g3953 ( 
.A1(n_3643),
.A2(n_3243),
.B1(n_3283),
.B2(n_3226),
.Y(n_3953)
);

OAI22xp5_ASAP7_75t_L g3954 ( 
.A1(n_3636),
.A2(n_3301),
.B1(n_3313),
.B2(n_3283),
.Y(n_3954)
);

HB1xp67_ASAP7_75t_L g3955 ( 
.A(n_3573),
.Y(n_3955)
);

OAI21xp33_ASAP7_75t_L g3956 ( 
.A1(n_3713),
.A2(n_3313),
.B(n_3301),
.Y(n_3956)
);

AOI22xp33_ASAP7_75t_SL g3957 ( 
.A1(n_3610),
.A2(n_3318),
.B1(n_3313),
.B2(n_272),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3572),
.Y(n_3958)
);

CKINVDCx20_ASAP7_75t_R g3959 ( 
.A(n_3404),
.Y(n_3959)
);

OAI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3453),
.A2(n_3318),
.B1(n_272),
.B2(n_269),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3581),
.Y(n_3961)
);

INVx1_ASAP7_75t_SL g3962 ( 
.A(n_3477),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3585),
.B(n_3589),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_SL g3964 ( 
.A1(n_3610),
.A2(n_3318),
.B1(n_274),
.B2(n_271),
.Y(n_3964)
);

INVxp67_ASAP7_75t_L g3965 ( 
.A(n_3508),
.Y(n_3965)
);

INVx5_ASAP7_75t_SL g3966 ( 
.A(n_3483),
.Y(n_3966)
);

NAND2x1p5_ASAP7_75t_L g3967 ( 
.A(n_3350),
.B(n_3491),
.Y(n_3967)
);

OR2x2_ASAP7_75t_SL g3968 ( 
.A(n_3331),
.B(n_271),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3704),
.B(n_273),
.Y(n_3969)
);

OAI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3427),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_3970)
);

OAI21xp5_ASAP7_75t_SL g3971 ( 
.A1(n_3413),
.A2(n_276),
.B(n_279),
.Y(n_3971)
);

INVx3_ASAP7_75t_L g3972 ( 
.A(n_3571),
.Y(n_3972)
);

OAI222xp33_ASAP7_75t_L g3973 ( 
.A1(n_3530),
.A2(n_284),
.B1(n_286),
.B2(n_280),
.C1(n_283),
.C2(n_285),
.Y(n_3973)
);

CKINVDCx5p33_ASAP7_75t_R g3974 ( 
.A(n_3455),
.Y(n_3974)
);

OAI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3605),
.A2(n_280),
.B(n_283),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_L g3976 ( 
.A1(n_3701),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_3976)
);

AOI222xp33_ASAP7_75t_L g3977 ( 
.A1(n_3447),
.A2(n_290),
.B1(n_292),
.B2(n_288),
.C1(n_289),
.C2(n_291),
.Y(n_3977)
);

OAI21xp33_ASAP7_75t_L g3978 ( 
.A1(n_3717),
.A2(n_289),
.B(n_290),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3625),
.B(n_292),
.Y(n_3979)
);

OAI22xp5_ASAP7_75t_L g3980 ( 
.A1(n_3644),
.A2(n_3372),
.B1(n_3548),
.B2(n_3533),
.Y(n_3980)
);

BUFx2_ASAP7_75t_SL g3981 ( 
.A(n_3389),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3578),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3598),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3613),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_L g3985 ( 
.A1(n_3708),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3600),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_SL g3987 ( 
.A1(n_3696),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_3987)
);

OAI22xp33_ASAP7_75t_SL g3988 ( 
.A1(n_3531),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_3988)
);

BUFx6f_ASAP7_75t_L g3989 ( 
.A(n_3441),
.Y(n_3989)
);

INVx2_ASAP7_75t_SL g3990 ( 
.A(n_3515),
.Y(n_3990)
);

INVx4_ASAP7_75t_SL g3991 ( 
.A(n_3480),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3708),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_3992)
);

AOI22xp33_ASAP7_75t_SL g3993 ( 
.A1(n_3702),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3993)
);

OAI21xp33_ASAP7_75t_L g3994 ( 
.A1(n_3470),
.A2(n_300),
.B(n_301),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3711),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3711),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_3996)
);

BUFx6f_ASAP7_75t_L g3997 ( 
.A(n_3441),
.Y(n_3997)
);

OAI21xp33_ASAP7_75t_L g3998 ( 
.A1(n_3545),
.A2(n_306),
.B(n_307),
.Y(n_3998)
);

OAI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_3372),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_3999)
);

OAI21xp5_ASAP7_75t_SL g4000 ( 
.A1(n_3403),
.A2(n_309),
.B(n_310),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_SL g4001 ( 
.A1(n_3599),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3714),
.A2(n_315),
.B1(n_312),
.B2(n_314),
.Y(n_4002)
);

INVx3_ASAP7_75t_L g4003 ( 
.A(n_3608),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_SL g4004 ( 
.A1(n_3638),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_3611),
.B(n_316),
.Y(n_4005)
);

INVx3_ASAP7_75t_L g4006 ( 
.A(n_3608),
.Y(n_4006)
);

NOR2x1_ASAP7_75t_R g4007 ( 
.A(n_3471),
.B(n_317),
.Y(n_4007)
);

BUFx4f_ASAP7_75t_SL g4008 ( 
.A(n_3416),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3659),
.B(n_318),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3714),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_4010)
);

AOI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3337),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_3458),
.Y(n_4012)
);

HB1xp67_ASAP7_75t_L g4013 ( 
.A(n_3409),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_3666),
.Y(n_4014)
);

HB1xp67_ASAP7_75t_SL g4015 ( 
.A(n_3538),
.Y(n_4015)
);

AOI22xp33_ASAP7_75t_SL g4016 ( 
.A1(n_3548),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_4016)
);

AOI22xp33_ASAP7_75t_L g4017 ( 
.A1(n_3715),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_4017)
);

OAI22xp5_ASAP7_75t_L g4018 ( 
.A1(n_3590),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_4018)
);

OAI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3458),
.A2(n_328),
.B1(n_325),
.B2(n_327),
.Y(n_4019)
);

OAI21xp33_ASAP7_75t_L g4020 ( 
.A1(n_3712),
.A2(n_328),
.B(n_329),
.Y(n_4020)
);

INVx2_ASAP7_75t_SL g4021 ( 
.A(n_3523),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3715),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3601),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_3716),
.A2(n_333),
.B1(n_330),
.B2(n_331),
.Y(n_4024)
);

AOI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3716),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_4025)
);

OAI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3665),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_4026)
);

OAI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3674),
.A2(n_341),
.B1(n_337),
.B2(n_338),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3669),
.Y(n_4028)
);

OAI22xp5_ASAP7_75t_SL g4029 ( 
.A1(n_3639),
.A2(n_343),
.B1(n_338),
.B2(n_342),
.Y(n_4029)
);

OAI21xp5_ASAP7_75t_SL g4030 ( 
.A1(n_3558),
.A2(n_342),
.B(n_343),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3602),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_SL g4032 ( 
.A1(n_3700),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_4032)
);

AOI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_3718),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_SL g4034 ( 
.A1(n_3700),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3671),
.Y(n_4035)
);

CKINVDCx6p67_ASAP7_75t_R g4036 ( 
.A(n_3523),
.Y(n_4036)
);

BUFx2_ASAP7_75t_L g4037 ( 
.A(n_3489),
.Y(n_4037)
);

HB1xp67_ASAP7_75t_L g4038 ( 
.A(n_3676),
.Y(n_4038)
);

OAI22xp5_ASAP7_75t_L g4039 ( 
.A1(n_3428),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_4039)
);

AND2x4_ASAP7_75t_L g4040 ( 
.A(n_3718),
.B(n_350),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3691),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3500),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_3326),
.Y(n_4043)
);

AOI222xp33_ASAP7_75t_L g4044 ( 
.A1(n_3476),
.A2(n_356),
.B1(n_358),
.B2(n_353),
.C1(n_354),
.C2(n_357),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3616),
.Y(n_4045)
);

AOI222xp33_ASAP7_75t_L g4046 ( 
.A1(n_3353),
.A2(n_3360),
.B1(n_3675),
.B2(n_3642),
.C1(n_3450),
.C2(n_3525),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3621),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3502),
.A2(n_358),
.B1(n_354),
.B2(n_357),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3699),
.Y(n_4049)
);

AOI22xp33_ASAP7_75t_SL g4050 ( 
.A1(n_3688),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_4050)
);

OAI22xp33_ASAP7_75t_L g4051 ( 
.A1(n_3558),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_4051)
);

OAI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3720),
.A2(n_365),
.B1(n_362),
.B2(n_363),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_SL g4053 ( 
.A1(n_3688),
.A2(n_365),
.B1(n_362),
.B2(n_363),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_3391),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3327),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_4055)
);

OAI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_3556),
.A2(n_369),
.B1(n_366),
.B2(n_368),
.Y(n_4056)
);

AOI22xp33_ASAP7_75t_L g4057 ( 
.A1(n_3727),
.A2(n_3837),
.B1(n_3780),
.B2(n_3729),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_4038),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3923),
.B(n_3628),
.Y(n_4059)
);

NAND3xp33_ASAP7_75t_L g4060 ( 
.A(n_3828),
.B(n_3656),
.C(n_3703),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3752),
.B(n_3498),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_4030),
.A2(n_3648),
.B1(n_3640),
.B2(n_3689),
.Y(n_4062)
);

OAI221xp5_ASAP7_75t_L g4063 ( 
.A1(n_3971),
.A2(n_3484),
.B1(n_3361),
.B2(n_3396),
.C(n_3423),
.Y(n_4063)
);

OAI22xp5_ASAP7_75t_L g4064 ( 
.A1(n_3743),
.A2(n_3689),
.B1(n_3592),
.B2(n_3687),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3743),
.A2(n_3672),
.B1(n_3673),
.B2(n_3663),
.Y(n_4065)
);

OAI221xp5_ASAP7_75t_L g4066 ( 
.A1(n_3733),
.A2(n_3401),
.B1(n_3577),
.B2(n_3684),
.C(n_3591),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3741),
.B(n_3682),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3756),
.A2(n_3499),
.B1(n_3521),
.B2(n_3512),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3829),
.Y(n_4069)
);

AOI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_4029),
.A2(n_3536),
.B1(n_3575),
.B2(n_3564),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3977),
.A2(n_3576),
.B1(n_3365),
.B2(n_3360),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3762),
.A2(n_3353),
.B1(n_3480),
.B2(n_3579),
.Y(n_4072)
);

AOI221xp5_ASAP7_75t_SL g4073 ( 
.A1(n_3968),
.A2(n_3410),
.B1(n_3667),
.B2(n_3478),
.C(n_3664),
.Y(n_4073)
);

AOI221xp5_ASAP7_75t_L g4074 ( 
.A1(n_3778),
.A2(n_3595),
.B1(n_3549),
.B2(n_3526),
.C(n_3587),
.Y(n_4074)
);

OAI22xp33_ASAP7_75t_L g4075 ( 
.A1(n_3768),
.A2(n_3651),
.B1(n_3662),
.B2(n_3591),
.Y(n_4075)
);

AOI22xp5_ASAP7_75t_SL g4076 ( 
.A1(n_3905),
.A2(n_3462),
.B1(n_3424),
.B2(n_3445),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3779),
.A2(n_3579),
.B1(n_3604),
.B2(n_3532),
.Y(n_4077)
);

OAI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_3809),
.A2(n_3604),
.B1(n_3684),
.B2(n_3662),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3758),
.A2(n_3637),
.B1(n_3721),
.B2(n_3706),
.Y(n_4079)
);

AOI22xp33_ASAP7_75t_L g4080 ( 
.A1(n_3793),
.A2(n_3706),
.B1(n_3721),
.B2(n_3624),
.Y(n_4080)
);

OAI22xp33_ASAP7_75t_L g4081 ( 
.A1(n_4000),
.A2(n_3623),
.B1(n_3539),
.B2(n_3606),
.Y(n_4081)
);

AOI22xp33_ASAP7_75t_L g4082 ( 
.A1(n_4044),
.A2(n_3624),
.B1(n_3614),
.B2(n_3554),
.Y(n_4082)
);

CKINVDCx20_ASAP7_75t_R g4083 ( 
.A(n_3847),
.Y(n_4083)
);

AOI22xp33_ASAP7_75t_L g4084 ( 
.A1(n_3964),
.A2(n_3629),
.B1(n_3449),
.B2(n_3460),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_3891),
.A2(n_3629),
.B1(n_3363),
.B2(n_3580),
.Y(n_4085)
);

NAND3xp33_ASAP7_75t_L g4086 ( 
.A(n_3955),
.B(n_3655),
.C(n_3694),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_SL g4087 ( 
.A(n_3941),
.B(n_3654),
.Y(n_4087)
);

AOI22xp33_ASAP7_75t_L g4088 ( 
.A1(n_3801),
.A2(n_3658),
.B1(n_3555),
.B2(n_3496),
.Y(n_4088)
);

OAI222xp33_ASAP7_75t_L g4089 ( 
.A1(n_3761),
.A2(n_3615),
.B1(n_3660),
.B2(n_3653),
.C1(n_3645),
.C2(n_3619),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3759),
.A2(n_3496),
.B1(n_3583),
.B2(n_3655),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3755),
.B(n_3492),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3830),
.B(n_3492),
.Y(n_4092)
);

AOI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_3787),
.A2(n_3657),
.B1(n_3538),
.B2(n_3681),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3833),
.B(n_3869),
.Y(n_4094)
);

AOI22xp33_ASAP7_75t_SL g4095 ( 
.A1(n_3736),
.A2(n_3492),
.B1(n_3574),
.B2(n_3509),
.Y(n_4095)
);

OAI211xp5_ASAP7_75t_L g4096 ( 
.A1(n_3770),
.A2(n_3650),
.B(n_3678),
.C(n_3633),
.Y(n_4096)
);

OAI22xp5_ASAP7_75t_L g4097 ( 
.A1(n_3782),
.A2(n_3457),
.B1(n_3528),
.B2(n_3509),
.Y(n_4097)
);

AOI22xp33_ASAP7_75t_L g4098 ( 
.A1(n_3970),
.A2(n_3509),
.B1(n_3618),
.B2(n_3574),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3878),
.Y(n_4099)
);

OAI22xp5_ASAP7_75t_SL g4100 ( 
.A1(n_3889),
.A2(n_3475),
.B1(n_3618),
.B2(n_3574),
.Y(n_4100)
);

AOI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_3726),
.A2(n_3661),
.B1(n_3618),
.B2(n_371),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_SL g4102 ( 
.A1(n_3748),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_4102)
);

AOI22xp33_ASAP7_75t_SL g4103 ( 
.A1(n_3764),
.A2(n_373),
.B1(n_370),
.B2(n_372),
.Y(n_4103)
);

AOI221xp5_ASAP7_75t_L g4104 ( 
.A1(n_3747),
.A2(n_376),
.B1(n_373),
.B2(n_375),
.C(n_377),
.Y(n_4104)
);

AOI22xp33_ASAP7_75t_L g4105 ( 
.A1(n_4018),
.A2(n_378),
.B1(n_375),
.B2(n_376),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3776),
.B(n_379),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3879),
.B(n_379),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_4026),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_L g4109 ( 
.A1(n_4027),
.A2(n_385),
.B1(n_381),
.B2(n_384),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_4052),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_4110)
);

AOI22xp33_ASAP7_75t_SL g4111 ( 
.A1(n_3764),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_4111)
);

AOI22xp33_ASAP7_75t_L g4112 ( 
.A1(n_3978),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3890),
.B(n_389),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3994),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3897),
.B(n_3915),
.Y(n_4115)
);

AOI22xp33_ASAP7_75t_L g4116 ( 
.A1(n_3998),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_SL g4117 ( 
.A1(n_3903),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_4117)
);

OAI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_3769),
.A2(n_3957),
.B1(n_3819),
.B2(n_3746),
.Y(n_4118)
);

AOI22xp33_ASAP7_75t_L g4119 ( 
.A1(n_3730),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_4119)
);

AOI22xp33_ASAP7_75t_L g4120 ( 
.A1(n_3987),
.A2(n_4019),
.B1(n_4040),
.B2(n_4001),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_3814),
.B(n_852),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_4040),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_4004),
.A2(n_4016),
.B1(n_3975),
.B2(n_4050),
.Y(n_4123)
);

AOI22xp33_ASAP7_75t_L g4124 ( 
.A1(n_4053),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_4124)
);

AOI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_3993),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3916),
.B(n_403),
.Y(n_4126)
);

AOI22xp33_ASAP7_75t_L g4127 ( 
.A1(n_3999),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3773),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_L g4129 ( 
.A1(n_4020),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_4129)
);

AOI22xp33_ASAP7_75t_L g4130 ( 
.A1(n_4056),
.A2(n_410),
.B1(n_407),
.B2(n_409),
.Y(n_4130)
);

AOI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_3751),
.A2(n_413),
.B1(n_410),
.B2(n_412),
.Y(n_4131)
);

AOI22xp33_ASAP7_75t_L g4132 ( 
.A1(n_4032),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4132)
);

OAI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_3818),
.A2(n_417),
.B1(n_414),
.B2(n_415),
.Y(n_4133)
);

AOI22xp33_ASAP7_75t_SL g4134 ( 
.A1(n_3926),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_3757),
.A2(n_421),
.B1(n_418),
.B2(n_420),
.Y(n_4135)
);

OAI22xp5_ASAP7_75t_L g4136 ( 
.A1(n_3766),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_4136)
);

OAI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_3802),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_4137)
);

AOI22xp33_ASAP7_75t_L g4138 ( 
.A1(n_4034),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4138)
);

NAND2xp33_ASAP7_75t_SL g4139 ( 
.A(n_3920),
.B(n_3935),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3945),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3922),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_3960),
.A2(n_430),
.B1(n_426),
.B2(n_429),
.Y(n_4142)
);

OAI22xp5_ASAP7_75t_L g4143 ( 
.A1(n_3885),
.A2(n_431),
.B1(n_426),
.B2(n_430),
.Y(n_4143)
);

OAI21xp5_ASAP7_75t_SL g4144 ( 
.A1(n_4046),
.A2(n_432),
.B(n_433),
.Y(n_4144)
);

AOI22xp33_ASAP7_75t_L g4145 ( 
.A1(n_3750),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_4145)
);

AOI22xp33_ASAP7_75t_SL g4146 ( 
.A1(n_4037),
.A2(n_437),
.B1(n_434),
.B2(n_436),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_SL g4147 ( 
.A1(n_3792),
.A2(n_3811),
.B1(n_3763),
.B2(n_3803),
.Y(n_4147)
);

AOI22xp33_ASAP7_75t_L g4148 ( 
.A1(n_3800),
.A2(n_439),
.B1(n_436),
.B2(n_438),
.Y(n_4148)
);

NAND3xp33_ASAP7_75t_SL g4149 ( 
.A(n_3791),
.B(n_438),
.C(n_439),
.Y(n_4149)
);

AOI22xp33_ASAP7_75t_L g4150 ( 
.A1(n_3796),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_4150)
);

OAI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3754),
.A2(n_444),
.B1(n_441),
.B2(n_443),
.Y(n_4151)
);

AOI22xp33_ASAP7_75t_SL g4152 ( 
.A1(n_3763),
.A2(n_3745),
.B1(n_3795),
.B2(n_3765),
.Y(n_4152)
);

AOI22xp33_ASAP7_75t_SL g4153 ( 
.A1(n_3763),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_4153)
);

AND2x2_ASAP7_75t_L g4154 ( 
.A(n_3846),
.B(n_852),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3932),
.B(n_446),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_3862),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_4156)
);

AOI22xp33_ASAP7_75t_SL g4157 ( 
.A1(n_3763),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_4157)
);

AOI22xp5_ASAP7_75t_L g4158 ( 
.A1(n_4039),
.A2(n_453),
.B1(n_450),
.B2(n_451),
.Y(n_4158)
);

AOI22xp33_ASAP7_75t_L g4159 ( 
.A1(n_4051),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_4159)
);

AOI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_4042),
.A2(n_459),
.B1(n_456),
.B2(n_457),
.Y(n_4160)
);

AOI22xp33_ASAP7_75t_L g4161 ( 
.A1(n_3919),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_4161)
);

OAI221xp5_ASAP7_75t_SL g4162 ( 
.A1(n_4048),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.C(n_464),
.Y(n_4162)
);

AOI22xp33_ASAP7_75t_SL g4163 ( 
.A1(n_3763),
.A2(n_465),
.B1(n_462),
.B2(n_464),
.Y(n_4163)
);

OAI222xp33_ASAP7_75t_L g4164 ( 
.A1(n_3784),
.A2(n_4015),
.B1(n_3912),
.B2(n_3732),
.C1(n_3783),
.C2(n_3786),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_SL g4165 ( 
.A1(n_4007),
.A2(n_465),
.B(n_466),
.Y(n_4165)
);

OAI221xp5_ASAP7_75t_SL g4166 ( 
.A1(n_4055),
.A2(n_470),
.B1(n_466),
.B2(n_467),
.C(n_471),
.Y(n_4166)
);

AOI22xp33_ASAP7_75t_L g4167 ( 
.A1(n_4013),
.A2(n_472),
.B1(n_467),
.B2(n_470),
.Y(n_4167)
);

OAI222xp33_ASAP7_75t_L g4168 ( 
.A1(n_3980),
.A2(n_476),
.B1(n_479),
.B2(n_473),
.C1(n_474),
.C2(n_478),
.Y(n_4168)
);

OAI22xp5_ASAP7_75t_L g4169 ( 
.A1(n_3820),
.A2(n_480),
.B1(n_473),
.B2(n_479),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_L g4170 ( 
.A1(n_3988),
.A2(n_483),
.B1(n_480),
.B2(n_481),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_L g4171 ( 
.A1(n_3798),
.A2(n_484),
.B1(n_481),
.B2(n_483),
.Y(n_4171)
);

AOI22xp5_ASAP7_75t_SL g4172 ( 
.A1(n_3805),
.A2(n_488),
.B1(n_486),
.B2(n_487),
.Y(n_4172)
);

NOR3xp33_ASAP7_75t_L g4173 ( 
.A(n_3973),
.B(n_486),
.C(n_487),
.Y(n_4173)
);

OAI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_3894),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_3948),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_4175)
);

AOI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_3812),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_4005),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3934),
.B(n_494),
.Y(n_4178)
);

AOI222xp33_ASAP7_75t_L g4179 ( 
.A1(n_4007),
.A2(n_498),
.B1(n_502),
.B2(n_496),
.C1(n_497),
.C2(n_501),
.Y(n_4179)
);

OAI222xp33_ASAP7_75t_L g4180 ( 
.A1(n_3860),
.A2(n_501),
.B1(n_503),
.B2(n_497),
.C1(n_498),
.C2(n_502),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3943),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_L g4182 ( 
.A1(n_3852),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_3865),
.A2(n_508),
.B1(n_505),
.B2(n_506),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3944),
.B(n_508),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3951),
.Y(n_4185)
);

OAI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_3826),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_3950),
.B(n_511),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3958),
.B(n_513),
.Y(n_4188)
);

AOI22xp33_ASAP7_75t_L g4189 ( 
.A1(n_3942),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_3858),
.A2(n_518),
.B1(n_515),
.B2(n_517),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3961),
.B(n_519),
.Y(n_4191)
);

OAI22xp33_ASAP7_75t_L g4192 ( 
.A1(n_4011),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_4192)
);

OAI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_3845),
.A2(n_3866),
.B1(n_3744),
.B2(n_3900),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_SL g4194 ( 
.A1(n_3745),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_4194)
);

AOI22xp33_ASAP7_75t_L g4195 ( 
.A1(n_3875),
.A2(n_527),
.B1(n_524),
.B2(n_525),
.Y(n_4195)
);

AOI22xp33_ASAP7_75t_L g4196 ( 
.A1(n_3884),
.A2(n_528),
.B1(n_524),
.B2(n_527),
.Y(n_4196)
);

OA21x2_ASAP7_75t_L g4197 ( 
.A1(n_3899),
.A2(n_528),
.B(n_529),
.Y(n_4197)
);

AOI22xp33_ASAP7_75t_SL g4198 ( 
.A1(n_3765),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_4198)
);

AOI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_3823),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3908),
.A2(n_3813),
.B1(n_3824),
.B2(n_3822),
.Y(n_4200)
);

AOI221xp5_ASAP7_75t_L g4201 ( 
.A1(n_3881),
.A2(n_539),
.B1(n_535),
.B2(n_537),
.C(n_540),
.Y(n_4201)
);

AOI221xp5_ASAP7_75t_SL g4202 ( 
.A1(n_3883),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.C(n_542),
.Y(n_4202)
);

AOI22xp33_ASAP7_75t_L g4203 ( 
.A1(n_3979),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_4203)
);

AOI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_3969),
.A2(n_546),
.B1(n_544),
.B2(n_545),
.Y(n_4204)
);

AOI22xp33_ASAP7_75t_L g4205 ( 
.A1(n_3902),
.A2(n_547),
.B1(n_545),
.B2(n_546),
.Y(n_4205)
);

OAI221xp5_ASAP7_75t_L g4206 ( 
.A1(n_3839),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.C(n_550),
.Y(n_4206)
);

AOI22xp33_ASAP7_75t_L g4207 ( 
.A1(n_3902),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3983),
.B(n_551),
.Y(n_4208)
);

OAI222xp33_ASAP7_75t_L g4209 ( 
.A1(n_3962),
.A2(n_552),
.B1(n_553),
.B2(n_555),
.C1(n_556),
.C2(n_557),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_3902),
.A2(n_560),
.B1(n_552),
.B2(n_559),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_3965),
.B(n_850),
.Y(n_4211)
);

AOI22xp33_ASAP7_75t_L g4212 ( 
.A1(n_3902),
.A2(n_562),
.B1(n_559),
.B2(n_560),
.Y(n_4212)
);

AOI22xp33_ASAP7_75t_L g4213 ( 
.A1(n_3902),
.A2(n_3940),
.B1(n_3856),
.B2(n_3976),
.Y(n_4213)
);

OAI221xp5_ASAP7_75t_L g4214 ( 
.A1(n_3832),
.A2(n_565),
.B1(n_562),
.B2(n_563),
.C(n_566),
.Y(n_4214)
);

OAI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_4036),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_4215)
);

AOI22xp33_ASAP7_75t_L g4216 ( 
.A1(n_3940),
.A2(n_571),
.B1(n_567),
.B2(n_569),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3986),
.B(n_569),
.Y(n_4217)
);

NAND3xp33_ASAP7_75t_L g4218 ( 
.A(n_3985),
.B(n_571),
.C(n_572),
.Y(n_4218)
);

AOI22xp33_ASAP7_75t_SL g4219 ( 
.A1(n_3795),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_4219)
);

AOI22xp33_ASAP7_75t_L g4220 ( 
.A1(n_3992),
.A2(n_576),
.B1(n_573),
.B2(n_575),
.Y(n_4220)
);

BUFx2_ASAP7_75t_L g4221 ( 
.A(n_3799),
.Y(n_4221)
);

OAI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_3827),
.A2(n_578),
.B1(n_575),
.B2(n_576),
.Y(n_4222)
);

AOI22xp33_ASAP7_75t_L g4223 ( 
.A1(n_3995),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4223)
);

NOR3xp33_ASAP7_75t_L g4224 ( 
.A(n_3936),
.B(n_579),
.C(n_580),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_3737),
.B(n_581),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_3996),
.A2(n_584),
.B1(n_581),
.B2(n_582),
.Y(n_4226)
);

AOI221xp5_ASAP7_75t_SL g4227 ( 
.A1(n_3918),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.C(n_589),
.Y(n_4227)
);

NAND4xp25_ASAP7_75t_L g4228 ( 
.A(n_4002),
.B(n_591),
.C(n_589),
.D(n_590),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_4023),
.B(n_590),
.Y(n_4229)
);

OAI22xp5_ASAP7_75t_L g4230 ( 
.A1(n_3874),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_4230)
);

AND2x2_ASAP7_75t_L g4231 ( 
.A(n_3749),
.B(n_843),
.Y(n_4231)
);

OAI222xp33_ASAP7_75t_L g4232 ( 
.A1(n_3864),
.A2(n_593),
.B1(n_594),
.B2(n_595),
.C1(n_596),
.C2(n_597),
.Y(n_4232)
);

AOI22xp33_ASAP7_75t_SL g4233 ( 
.A1(n_3871),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_4233)
);

AOI22xp5_ASAP7_75t_L g4234 ( 
.A1(n_3840),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3928),
.A2(n_601),
.B1(n_598),
.B2(n_599),
.Y(n_4235)
);

AOI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_4010),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_4236)
);

AOI22xp33_ASAP7_75t_L g4237 ( 
.A1(n_4017),
.A2(n_608),
.B1(n_603),
.B2(n_605),
.Y(n_4237)
);

AOI22xp33_ASAP7_75t_L g4238 ( 
.A1(n_4022),
.A2(n_611),
.B1(n_608),
.B2(n_610),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3854),
.Y(n_4239)
);

AOI21xp33_ASAP7_75t_SL g4240 ( 
.A1(n_4021),
.A2(n_610),
.B(n_613),
.Y(n_4240)
);

AOI22xp33_ASAP7_75t_L g4241 ( 
.A1(n_4031),
.A2(n_616),
.B1(n_613),
.B2(n_615),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4045),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_4242)
);

OAI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_3850),
.A2(n_619),
.B1(n_617),
.B2(n_618),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_4047),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_4244)
);

AOI22xp33_ASAP7_75t_L g4245 ( 
.A1(n_4024),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_4245)
);

AOI22xp5_ASAP7_75t_L g4246 ( 
.A1(n_3861),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_4246)
);

AOI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_4025),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_4247)
);

AOI22xp33_ASAP7_75t_L g4248 ( 
.A1(n_4033),
.A2(n_630),
.B1(n_625),
.B2(n_629),
.Y(n_4248)
);

OAI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_3880),
.A2(n_632),
.B1(n_630),
.B2(n_631),
.Y(n_4249)
);

NAND3xp33_ASAP7_75t_L g4250 ( 
.A(n_3909),
.B(n_3831),
.C(n_3895),
.Y(n_4250)
);

AOI22xp33_ASAP7_75t_L g4251 ( 
.A1(n_4009),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.Y(n_4251)
);

NOR2x1_ASAP7_75t_SL g4252 ( 
.A(n_3981),
.B(n_633),
.Y(n_4252)
);

INVxp67_ASAP7_75t_L g4253 ( 
.A(n_3810),
.Y(n_4253)
);

AOI22xp33_ASAP7_75t_L g4254 ( 
.A1(n_3956),
.A2(n_637),
.B1(n_634),
.B2(n_636),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_3931),
.A2(n_638),
.B1(n_636),
.B2(n_637),
.Y(n_4255)
);

AOI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_3821),
.A2(n_641),
.B1(n_638),
.B2(n_639),
.Y(n_4256)
);

AOI22xp33_ASAP7_75t_SL g4257 ( 
.A1(n_3871),
.A2(n_642),
.B1(n_639),
.B2(n_641),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_3734),
.B(n_642),
.Y(n_4258)
);

OAI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_3841),
.A2(n_645),
.B1(n_643),
.B2(n_644),
.Y(n_4259)
);

NAND3xp33_ASAP7_75t_L g4260 ( 
.A(n_3910),
.B(n_643),
.C(n_644),
.Y(n_4260)
);

CKINVDCx5p33_ASAP7_75t_R g4261 ( 
.A(n_3774),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_3886),
.B(n_645),
.Y(n_4262)
);

OAI22xp5_ASAP7_75t_L g4263 ( 
.A1(n_3848),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_4263)
);

AOI22xp33_ASAP7_75t_L g4264 ( 
.A1(n_3843),
.A2(n_649),
.B1(n_646),
.B2(n_648),
.Y(n_4264)
);

AOI22xp33_ASAP7_75t_L g4265 ( 
.A1(n_3887),
.A2(n_652),
.B1(n_649),
.B2(n_650),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_3738),
.B(n_3739),
.Y(n_4266)
);

AOI22xp33_ASAP7_75t_L g4267 ( 
.A1(n_3740),
.A2(n_655),
.B1(n_650),
.B2(n_654),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3742),
.B(n_654),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_3868),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_3873),
.Y(n_4270)
);

AOI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_3753),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.Y(n_4271)
);

OAI22xp5_ASAP7_75t_L g4272 ( 
.A1(n_4072),
.A2(n_3972),
.B1(n_4006),
.B2(n_4003),
.Y(n_4272)
);

AND2x4_ASAP7_75t_L g4273 ( 
.A(n_4058),
.B(n_3772),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_SL g4274 ( 
.A(n_4075),
.B(n_3972),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_R g4275 ( 
.A(n_4083),
.B(n_3735),
.Y(n_4275)
);

OAI21xp5_ASAP7_75t_SL g4276 ( 
.A1(n_4144),
.A2(n_3731),
.B(n_3872),
.Y(n_4276)
);

OAI221xp5_ASAP7_75t_SL g4277 ( 
.A1(n_4057),
.A2(n_3851),
.B1(n_3867),
.B2(n_3877),
.C(n_3929),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4061),
.B(n_4067),
.Y(n_4278)
);

NOR2xp33_ASAP7_75t_L g4279 ( 
.A(n_4253),
.B(n_3990),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_4221),
.B(n_3775),
.Y(n_4280)
);

NAND3xp33_ASAP7_75t_L g4281 ( 
.A(n_4073),
.B(n_3947),
.C(n_3949),
.Y(n_4281)
);

NOR3xp33_ASAP7_75t_L g4282 ( 
.A(n_4149),
.B(n_4006),
.C(n_4003),
.Y(n_4282)
);

NAND3xp33_ASAP7_75t_SL g4283 ( 
.A(n_4179),
.B(n_3959),
.C(n_4043),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4059),
.B(n_3781),
.Y(n_4284)
);

AOI22xp33_ASAP7_75t_L g4285 ( 
.A1(n_4173),
.A2(n_4224),
.B1(n_4077),
.B2(n_4071),
.Y(n_4285)
);

OAI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4072),
.A2(n_3966),
.B1(n_3906),
.B2(n_3836),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4140),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4069),
.B(n_3785),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4099),
.B(n_3788),
.Y(n_4289)
);

NOR3xp33_ASAP7_75t_L g4290 ( 
.A(n_4060),
.B(n_4063),
.C(n_4209),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4141),
.B(n_3789),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4181),
.B(n_3790),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4094),
.B(n_3794),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_4091),
.B(n_3807),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4185),
.B(n_3815),
.Y(n_4295)
);

NAND3xp33_ASAP7_75t_L g4296 ( 
.A(n_4202),
.B(n_3904),
.C(n_3842),
.Y(n_4296)
);

NAND3xp33_ASAP7_75t_L g4297 ( 
.A(n_4227),
.B(n_3834),
.C(n_3863),
.Y(n_4297)
);

OAI211xp5_ASAP7_75t_L g4298 ( 
.A1(n_4165),
.A2(n_4068),
.B(n_4085),
.C(n_4080),
.Y(n_4298)
);

AND2x2_ASAP7_75t_SL g4299 ( 
.A(n_4197),
.B(n_3816),
.Y(n_4299)
);

AOI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4081),
.A2(n_3882),
.B(n_3939),
.Y(n_4300)
);

OR2x2_ASAP7_75t_L g4301 ( 
.A(n_4115),
.B(n_3963),
.Y(n_4301)
);

OAI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4249),
.A2(n_3898),
.B(n_3849),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4239),
.B(n_4269),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4068),
.B(n_3913),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4266),
.B(n_3917),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4270),
.B(n_3924),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4065),
.B(n_3982),
.Y(n_4307)
);

NAND3xp33_ASAP7_75t_L g4308 ( 
.A(n_4250),
.B(n_3952),
.C(n_3914),
.Y(n_4308)
);

OAI22xp5_ASAP7_75t_L g4309 ( 
.A1(n_4070),
.A2(n_3966),
.B1(n_3893),
.B2(n_3937),
.Y(n_4309)
);

AND2x2_ASAP7_75t_L g4310 ( 
.A(n_4106),
.B(n_3984),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4154),
.B(n_4014),
.Y(n_4311)
);

OAI21xp5_ASAP7_75t_SL g4312 ( 
.A1(n_4081),
.A2(n_3967),
.B(n_3870),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4065),
.B(n_4028),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4074),
.B(n_4121),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4092),
.B(n_4035),
.Y(n_4315)
);

NAND4xp25_ASAP7_75t_L g4316 ( 
.A(n_4071),
.B(n_4012),
.C(n_3728),
.D(n_3767),
.Y(n_4316)
);

OAI221xp5_ASAP7_75t_SL g4317 ( 
.A1(n_4120),
.A2(n_3777),
.B1(n_3771),
.B2(n_3760),
.C(n_3804),
.Y(n_4317)
);

AND2x2_ASAP7_75t_L g4318 ( 
.A(n_4200),
.B(n_4041),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4225),
.B(n_4049),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4231),
.B(n_3808),
.Y(n_4320)
);

AOI22xp33_ASAP7_75t_L g4321 ( 
.A1(n_4118),
.A2(n_3930),
.B1(n_3855),
.B2(n_3901),
.Y(n_4321)
);

OA21x2_ASAP7_75t_L g4322 ( 
.A1(n_4087),
.A2(n_3825),
.B(n_3888),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4107),
.B(n_3806),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4113),
.B(n_4126),
.Y(n_4324)
);

OAI221xp5_ASAP7_75t_L g4325 ( 
.A1(n_4082),
.A2(n_3911),
.B1(n_3921),
.B2(n_3954),
.C(n_3953),
.Y(n_4325)
);

OAI221xp5_ASAP7_75t_SL g4326 ( 
.A1(n_4070),
.A2(n_3853),
.B1(n_3933),
.B2(n_3816),
.C(n_3991),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4155),
.B(n_3806),
.Y(n_4327)
);

OAI21xp5_ASAP7_75t_SL g4328 ( 
.A1(n_4164),
.A2(n_4147),
.B(n_4084),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4178),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4184),
.B(n_3806),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4213),
.B(n_3844),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4187),
.B(n_3844),
.Y(n_4332)
);

NAND3xp33_ASAP7_75t_L g4333 ( 
.A(n_4102),
.B(n_3844),
.C(n_3876),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4188),
.B(n_3855),
.Y(n_4334)
);

NAND4xp25_ASAP7_75t_L g4335 ( 
.A(n_4172),
.B(n_3857),
.C(n_3859),
.D(n_3933),
.Y(n_4335)
);

OAI22xp5_ASAP7_75t_L g4336 ( 
.A1(n_4123),
.A2(n_3817),
.B1(n_3797),
.B2(n_3892),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_SL g4337 ( 
.A(n_4075),
.B(n_3991),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4191),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_4208),
.B(n_3855),
.Y(n_4339)
);

OAI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4249),
.A2(n_3855),
.B(n_3974),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4217),
.B(n_3896),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4211),
.B(n_4197),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4088),
.A2(n_3907),
.B1(n_4008),
.B2(n_3927),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_4229),
.B(n_3896),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_4258),
.B(n_3896),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4268),
.Y(n_4346)
);

OAI221xp5_ASAP7_75t_L g4347 ( 
.A1(n_4103),
.A2(n_4054),
.B1(n_3997),
.B2(n_3989),
.C(n_3946),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4151),
.B(n_3997),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4151),
.B(n_3997),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_4193),
.B(n_3925),
.Y(n_4350)
);

NOR2xp33_ASAP7_75t_L g4351 ( 
.A(n_4066),
.B(n_3838),
.Y(n_4351)
);

NAND4xp25_ASAP7_75t_L g4352 ( 
.A(n_4111),
.B(n_3835),
.C(n_660),
.D(n_656),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_L g4353 ( 
.A(n_4076),
.B(n_659),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4101),
.B(n_3989),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4079),
.B(n_3989),
.Y(n_4355)
);

NAND4xp25_ASAP7_75t_SL g4356 ( 
.A(n_4090),
.B(n_661),
.C(n_659),
.D(n_660),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4064),
.B(n_4097),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4197),
.B(n_3925),
.Y(n_4358)
);

AOI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_4228),
.A2(n_3938),
.B1(n_3946),
.B2(n_3925),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_4252),
.B(n_3946),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4093),
.B(n_4176),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4095),
.B(n_3938),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4139),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4152),
.B(n_3938),
.Y(n_4364)
);

AOI21xp5_ASAP7_75t_L g4365 ( 
.A1(n_4089),
.A2(n_661),
.B(n_662),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4271),
.B(n_662),
.Y(n_4366)
);

OAI22xp5_ASAP7_75t_L g4367 ( 
.A1(n_4262),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4086),
.B(n_663),
.Y(n_4368)
);

OAI22xp5_ASAP7_75t_L g4369 ( 
.A1(n_4117),
.A2(n_669),
.B1(n_666),
.B2(n_667),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_SL g4370 ( 
.A(n_4100),
.B(n_670),
.Y(n_4370)
);

NAND3xp33_ASAP7_75t_L g4371 ( 
.A(n_4254),
.B(n_671),
.C(n_672),
.Y(n_4371)
);

OAI21xp5_ASAP7_75t_L g4372 ( 
.A1(n_4215),
.A2(n_671),
.B(n_672),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_4215),
.B(n_673),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_4280),
.B(n_4098),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_4294),
.B(n_4078),
.Y(n_4375)
);

NOR3xp33_ASAP7_75t_L g4376 ( 
.A(n_4283),
.B(n_4168),
.C(n_4180),
.Y(n_4376)
);

AOI22xp5_ASAP7_75t_L g4377 ( 
.A1(n_4316),
.A2(n_4174),
.B1(n_4146),
.B2(n_4134),
.Y(n_4377)
);

NOR3xp33_ASAP7_75t_L g4378 ( 
.A(n_4328),
.B(n_4232),
.C(n_4260),
.Y(n_4378)
);

OR2x2_ASAP7_75t_L g4379 ( 
.A(n_4278),
.B(n_4301),
.Y(n_4379)
);

OAI221xp5_ASAP7_75t_L g4380 ( 
.A1(n_4328),
.A2(n_4175),
.B1(n_4219),
.B2(n_4198),
.C(n_4194),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4303),
.B(n_4062),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4318),
.B(n_4199),
.Y(n_4382)
);

OAI21xp33_ASAP7_75t_L g4383 ( 
.A1(n_4290),
.A2(n_4316),
.B(n_4312),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4273),
.Y(n_4384)
);

AOI211xp5_ASAP7_75t_L g4385 ( 
.A1(n_4312),
.A2(n_4096),
.B(n_4240),
.C(n_4133),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_4315),
.B(n_4234),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4273),
.B(n_4271),
.Y(n_4387)
);

NOR3xp33_ASAP7_75t_L g4388 ( 
.A(n_4298),
.B(n_4214),
.C(n_4206),
.Y(n_4388)
);

HB1xp67_ASAP7_75t_L g4389 ( 
.A(n_4287),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4306),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_4310),
.B(n_4246),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4295),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_L g4393 ( 
.A1(n_4357),
.A2(n_4201),
.B1(n_4263),
.B2(n_4186),
.Y(n_4393)
);

OR2x2_ASAP7_75t_L g4394 ( 
.A(n_4284),
.B(n_4143),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4331),
.B(n_4265),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4311),
.B(n_4150),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4288),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4346),
.B(n_4304),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4363),
.B(n_4122),
.Y(n_4399)
);

NOR2x1_ASAP7_75t_L g4400 ( 
.A(n_4337),
.B(n_4136),
.Y(n_4400)
);

NAND3xp33_ASAP7_75t_L g4401 ( 
.A(n_4350),
.B(n_4116),
.C(n_4114),
.Y(n_4401)
);

NOR2xp67_ASAP7_75t_L g4402 ( 
.A(n_4335),
.B(n_4261),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_SL g4403 ( 
.A(n_4299),
.B(n_4153),
.Y(n_4403)
);

NAND4xp75_ASAP7_75t_L g4404 ( 
.A(n_4340),
.B(n_4351),
.C(n_4322),
.D(n_4365),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4279),
.B(n_4205),
.Y(n_4405)
);

OR2x2_ASAP7_75t_L g4406 ( 
.A(n_4293),
.B(n_4241),
.Y(n_4406)
);

INVxp67_ASAP7_75t_SL g4407 ( 
.A(n_4274),
.Y(n_4407)
);

OR2x2_ASAP7_75t_L g4408 ( 
.A(n_4305),
.B(n_4241),
.Y(n_4408)
);

NAND3xp33_ASAP7_75t_L g4409 ( 
.A(n_4322),
.B(n_4244),
.C(n_4242),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4329),
.B(n_4242),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_4338),
.B(n_4342),
.Y(n_4411)
);

NOR2xp33_ASAP7_75t_L g4412 ( 
.A(n_4343),
.B(n_4160),
.Y(n_4412)
);

OR2x2_ASAP7_75t_L g4413 ( 
.A(n_4289),
.B(n_4244),
.Y(n_4413)
);

NAND3xp33_ASAP7_75t_L g4414 ( 
.A(n_4321),
.B(n_4170),
.C(n_4163),
.Y(n_4414)
);

AOI221xp5_ASAP7_75t_L g4415 ( 
.A1(n_4317),
.A2(n_4192),
.B1(n_4137),
.B2(n_4162),
.C(n_4166),
.Y(n_4415)
);

OR2x2_ASAP7_75t_L g4416 ( 
.A(n_4291),
.B(n_4255),
.Y(n_4416)
);

AOI221xp5_ASAP7_75t_L g4417 ( 
.A1(n_4285),
.A2(n_4192),
.B1(n_4169),
.B2(n_4128),
.C(n_4104),
.Y(n_4417)
);

AO22x1_ASAP7_75t_L g4418 ( 
.A1(n_4309),
.A2(n_4235),
.B1(n_4230),
.B2(n_4135),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4364),
.B(n_4158),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4362),
.B(n_4207),
.Y(n_4420)
);

NAND3xp33_ASAP7_75t_L g4421 ( 
.A(n_4281),
.B(n_4157),
.C(n_4129),
.Y(n_4421)
);

NAND3xp33_ASAP7_75t_L g4422 ( 
.A(n_4308),
.B(n_4257),
.C(n_4233),
.Y(n_4422)
);

NOR3xp33_ASAP7_75t_SL g4423 ( 
.A(n_4326),
.B(n_4243),
.C(n_4259),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4292),
.Y(n_4424)
);

HB1xp67_ASAP7_75t_L g4425 ( 
.A(n_4319),
.Y(n_4425)
);

OR2x2_ASAP7_75t_L g4426 ( 
.A(n_4320),
.B(n_4222),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4307),
.B(n_4119),
.Y(n_4427)
);

INVxp67_ASAP7_75t_L g4428 ( 
.A(n_4353),
.Y(n_4428)
);

CKINVDCx5p33_ASAP7_75t_R g4429 ( 
.A(n_4275),
.Y(n_4429)
);

OR2x2_ASAP7_75t_L g4430 ( 
.A(n_4313),
.B(n_4210),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4314),
.B(n_4190),
.Y(n_4431)
);

NAND3xp33_ASAP7_75t_L g4432 ( 
.A(n_4282),
.B(n_4112),
.C(n_4212),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4324),
.B(n_4177),
.Y(n_4433)
);

OR2x2_ASAP7_75t_L g4434 ( 
.A(n_4355),
.B(n_674),
.Y(n_4434)
);

NAND3xp33_ASAP7_75t_L g4435 ( 
.A(n_4296),
.B(n_4171),
.C(n_4148),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4358),
.B(n_4145),
.Y(n_4436)
);

NOR2x1_ASAP7_75t_L g4437 ( 
.A(n_4335),
.B(n_4218),
.Y(n_4437)
);

OR2x2_ASAP7_75t_L g4438 ( 
.A(n_4345),
.B(n_674),
.Y(n_4438)
);

NAND3xp33_ASAP7_75t_L g4439 ( 
.A(n_4276),
.B(n_4182),
.C(n_4131),
.Y(n_4439)
);

AOI211xp5_ASAP7_75t_L g4440 ( 
.A1(n_4352),
.A2(n_4125),
.B(n_4124),
.C(n_4108),
.Y(n_4440)
);

NAND4xp75_ASAP7_75t_L g4441 ( 
.A(n_4300),
.B(n_4370),
.C(n_4368),
.D(n_4302),
.Y(n_4441)
);

NAND4xp75_ASAP7_75t_L g4442 ( 
.A(n_4361),
.B(n_4196),
.C(n_4204),
.D(n_4195),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4341),
.Y(n_4443)
);

NOR3xp33_ASAP7_75t_L g4444 ( 
.A(n_4352),
.B(n_4336),
.C(n_4356),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_4297),
.B(n_4348),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4334),
.B(n_4216),
.Y(n_4446)
);

AOI22xp5_ASAP7_75t_L g4447 ( 
.A1(n_4276),
.A2(n_4203),
.B1(n_4109),
.B2(n_4110),
.Y(n_4447)
);

AND2x2_ASAP7_75t_L g4448 ( 
.A(n_4339),
.B(n_4323),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4344),
.Y(n_4449)
);

AOI22xp33_ASAP7_75t_L g4450 ( 
.A1(n_4373),
.A2(n_4142),
.B1(n_4105),
.B2(n_4159),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4327),
.B(n_4264),
.Y(n_4451)
);

NOR2xp33_ASAP7_75t_L g4452 ( 
.A(n_4347),
.B(n_4156),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4389),
.Y(n_4453)
);

NOR2xp33_ASAP7_75t_L g4454 ( 
.A(n_4428),
.B(n_4277),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4411),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_4429),
.B(n_4286),
.Y(n_4456)
);

INVxp67_ASAP7_75t_SL g4457 ( 
.A(n_4402),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4443),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4398),
.B(n_4349),
.Y(n_4459)
);

AOI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_4403),
.A2(n_4383),
.B(n_4402),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4397),
.Y(n_4461)
);

NAND4xp75_ASAP7_75t_SL g4462 ( 
.A(n_4452),
.B(n_4360),
.C(n_4372),
.D(n_4359),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4448),
.B(n_4330),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4424),
.Y(n_4464)
);

NAND3xp33_ASAP7_75t_SL g4465 ( 
.A(n_4383),
.B(n_4272),
.C(n_4333),
.Y(n_4465)
);

OR2x2_ASAP7_75t_L g4466 ( 
.A(n_4379),
.B(n_4332),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4392),
.Y(n_4467)
);

XNOR2xp5_ASAP7_75t_L g4468 ( 
.A(n_4441),
.B(n_4367),
.Y(n_4468)
);

XNOR2x2_ASAP7_75t_L g4469 ( 
.A(n_4404),
.B(n_4325),
.Y(n_4469)
);

AND2x4_ASAP7_75t_L g4470 ( 
.A(n_4407),
.B(n_4354),
.Y(n_4470)
);

BUFx3_ASAP7_75t_L g4471 ( 
.A(n_4390),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4425),
.Y(n_4472)
);

XNOR2xp5_ASAP7_75t_L g4473 ( 
.A(n_4381),
.B(n_4369),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4449),
.Y(n_4474)
);

AND2x2_ASAP7_75t_L g4475 ( 
.A(n_4374),
.B(n_4366),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4384),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4445),
.Y(n_4477)
);

NAND3xp33_ASAP7_75t_L g4478 ( 
.A(n_4378),
.B(n_4371),
.C(n_4167),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4375),
.B(n_4251),
.Y(n_4479)
);

NAND2xp33_ASAP7_75t_SL g4480 ( 
.A(n_4423),
.B(n_4132),
.Y(n_4480)
);

AND2x2_ASAP7_75t_L g4481 ( 
.A(n_4419),
.B(n_4161),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_4387),
.B(n_4267),
.Y(n_4482)
);

NAND4xp75_ASAP7_75t_SL g4483 ( 
.A(n_4412),
.B(n_4256),
.C(n_4138),
.D(n_4189),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4419),
.B(n_4127),
.Y(n_4484)
);

XOR2x2_ASAP7_75t_L g4485 ( 
.A(n_4444),
.B(n_4183),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4399),
.Y(n_4486)
);

OR2x2_ASAP7_75t_L g4487 ( 
.A(n_4408),
.B(n_4430),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_L g4488 ( 
.A(n_4431),
.B(n_675),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4413),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_4406),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_4386),
.Y(n_4491)
);

OR2x2_ASAP7_75t_L g4492 ( 
.A(n_4410),
.B(n_675),
.Y(n_4492)
);

XNOR2xp5_ASAP7_75t_L g4493 ( 
.A(n_4437),
.B(n_4130),
.Y(n_4493)
);

INVx1_ASAP7_75t_SL g4494 ( 
.A(n_4438),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4416),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4394),
.Y(n_4496)
);

AND2x4_ASAP7_75t_L g4497 ( 
.A(n_4436),
.B(n_676),
.Y(n_4497)
);

OR2x2_ASAP7_75t_L g4498 ( 
.A(n_4426),
.B(n_4382),
.Y(n_4498)
);

INVx4_ASAP7_75t_L g4499 ( 
.A(n_4434),
.Y(n_4499)
);

INVx2_ASAP7_75t_SL g4500 ( 
.A(n_4400),
.Y(n_4500)
);

NOR4xp25_ASAP7_75t_L g4501 ( 
.A(n_4409),
.B(n_4223),
.C(n_4226),
.D(n_4220),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4420),
.B(n_4236),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4427),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4391),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4395),
.B(n_4237),
.Y(n_4505)
);

INVx2_ASAP7_75t_SL g4506 ( 
.A(n_4396),
.Y(n_4506)
);

NAND3xp33_ASAP7_75t_L g4507 ( 
.A(n_4376),
.B(n_4248),
.C(n_4245),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4446),
.Y(n_4508)
);

AOI211xp5_ASAP7_75t_SL g4509 ( 
.A1(n_4385),
.A2(n_4247),
.B(n_4238),
.C(n_678),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4451),
.Y(n_4510)
);

AO22x2_ASAP7_75t_L g4511 ( 
.A1(n_4421),
.A2(n_4439),
.B1(n_4414),
.B2(n_4442),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_4433),
.B(n_4405),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4401),
.B(n_676),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4432),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4377),
.B(n_677),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_L g4516 ( 
.A(n_4380),
.B(n_677),
.Y(n_4516)
);

INVx2_ASAP7_75t_SL g4517 ( 
.A(n_4422),
.Y(n_4517)
);

OR2x2_ASAP7_75t_L g4518 ( 
.A(n_4435),
.B(n_840),
.Y(n_4518)
);

BUFx3_ASAP7_75t_L g4519 ( 
.A(n_4377),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4418),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4447),
.Y(n_4521)
);

OR2x2_ASAP7_75t_L g4522 ( 
.A(n_4489),
.B(n_4447),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4496),
.Y(n_4523)
);

XOR2x2_ASAP7_75t_L g4524 ( 
.A(n_4469),
.B(n_4388),
.Y(n_4524)
);

OAI22x1_ASAP7_75t_L g4525 ( 
.A1(n_4500),
.A2(n_4440),
.B1(n_4415),
.B2(n_4417),
.Y(n_4525)
);

INVxp67_ASAP7_75t_L g4526 ( 
.A(n_4456),
.Y(n_4526)
);

NAND2xp33_ASAP7_75t_R g4527 ( 
.A(n_4460),
.B(n_678),
.Y(n_4527)
);

XNOR2xp5_ASAP7_75t_L g4528 ( 
.A(n_4511),
.B(n_4440),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4521),
.B(n_4503),
.Y(n_4529)
);

XNOR2xp5_ASAP7_75t_L g4530 ( 
.A(n_4511),
.B(n_4393),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4471),
.Y(n_4531)
);

OR2x2_ASAP7_75t_L g4532 ( 
.A(n_4490),
.B(n_4450),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4453),
.Y(n_4533)
);

OR2x2_ASAP7_75t_L g4534 ( 
.A(n_4487),
.B(n_679),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4495),
.Y(n_4535)
);

INVx1_ASAP7_75t_SL g4536 ( 
.A(n_4494),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4472),
.Y(n_4537)
);

AO22x2_ASAP7_75t_L g4538 ( 
.A1(n_4520),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4503),
.B(n_680),
.Y(n_4539)
);

XOR2x2_ASAP7_75t_L g4540 ( 
.A(n_4519),
.B(n_682),
.Y(n_4540)
);

OA22x2_ASAP7_75t_L g4541 ( 
.A1(n_4517),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4510),
.Y(n_4542)
);

XOR2x1_ASAP7_75t_L g4543 ( 
.A(n_4485),
.B(n_683),
.Y(n_4543)
);

OR2x2_ASAP7_75t_L g4544 ( 
.A(n_4477),
.B(n_684),
.Y(n_4544)
);

INVxp67_ASAP7_75t_L g4545 ( 
.A(n_4513),
.Y(n_4545)
);

XOR2xp5_ASAP7_75t_L g4546 ( 
.A(n_4473),
.B(n_686),
.Y(n_4546)
);

XNOR2x1_ASAP7_75t_L g4547 ( 
.A(n_4468),
.B(n_686),
.Y(n_4547)
);

XOR2x2_ASAP7_75t_L g4548 ( 
.A(n_4454),
.B(n_687),
.Y(n_4548)
);

XOR2x2_ASAP7_75t_L g4549 ( 
.A(n_4465),
.B(n_688),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4470),
.B(n_689),
.Y(n_4550)
);

XNOR2x2_ASAP7_75t_L g4551 ( 
.A(n_4493),
.B(n_4514),
.Y(n_4551)
);

XNOR2x1_ASAP7_75t_L g4552 ( 
.A(n_4462),
.B(n_689),
.Y(n_4552)
);

XNOR2x1_ASAP7_75t_L g4553 ( 
.A(n_4515),
.B(n_690),
.Y(n_4553)
);

BUFx3_ASAP7_75t_L g4554 ( 
.A(n_4453),
.Y(n_4554)
);

INVxp67_ASAP7_75t_L g4555 ( 
.A(n_4518),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4510),
.Y(n_4556)
);

AOI22xp5_ASAP7_75t_L g4557 ( 
.A1(n_4480),
.A2(n_690),
.B1(n_691),
.B2(n_692),
.Y(n_4557)
);

XNOR2x2_ASAP7_75t_L g4558 ( 
.A(n_4478),
.B(n_691),
.Y(n_4558)
);

NOR2x1_ASAP7_75t_L g4559 ( 
.A(n_4497),
.B(n_692),
.Y(n_4559)
);

XNOR2xp5_ASAP7_75t_L g4560 ( 
.A(n_4497),
.B(n_693),
.Y(n_4560)
);

NOR2xp33_ASAP7_75t_L g4561 ( 
.A(n_4512),
.B(n_4498),
.Y(n_4561)
);

XNOR2xp5_ASAP7_75t_L g4562 ( 
.A(n_4457),
.B(n_693),
.Y(n_4562)
);

INVxp67_ASAP7_75t_L g4563 ( 
.A(n_4516),
.Y(n_4563)
);

XNOR2x2_ASAP7_75t_L g4564 ( 
.A(n_4507),
.B(n_694),
.Y(n_4564)
);

HB1xp67_ASAP7_75t_L g4565 ( 
.A(n_4532),
.Y(n_4565)
);

INVxp67_ASAP7_75t_L g4566 ( 
.A(n_4538),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4554),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4533),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4542),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4531),
.Y(n_4570)
);

OA22x2_ASAP7_75t_L g4571 ( 
.A1(n_4528),
.A2(n_4499),
.B1(n_4508),
.B2(n_4506),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4556),
.Y(n_4572)
);

XNOR2xp5_ASAP7_75t_L g4573 ( 
.A(n_4524),
.B(n_4483),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4537),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4555),
.B(n_4470),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4523),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4535),
.Y(n_4577)
);

OA22x2_ASAP7_75t_L g4578 ( 
.A1(n_4528),
.A2(n_4499),
.B1(n_4508),
.B2(n_4504),
.Y(n_4578)
);

AOI22x1_ASAP7_75t_L g4579 ( 
.A1(n_4525),
.A2(n_4509),
.B1(n_4481),
.B2(n_4484),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4536),
.Y(n_4580)
);

OA22x2_ASAP7_75t_L g4581 ( 
.A1(n_4530),
.A2(n_4504),
.B1(n_4486),
.B2(n_4459),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4529),
.Y(n_4582)
);

OA22x2_ASAP7_75t_L g4583 ( 
.A1(n_4526),
.A2(n_4491),
.B1(n_4475),
.B2(n_4461),
.Y(n_4583)
);

OAI22xp5_ASAP7_75t_L g4584 ( 
.A1(n_4559),
.A2(n_4482),
.B1(n_4466),
.B2(n_4455),
.Y(n_4584)
);

BUFx3_ASAP7_75t_L g4585 ( 
.A(n_4550),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4538),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4522),
.Y(n_4587)
);

XNOR2xp5_ASAP7_75t_L g4588 ( 
.A(n_4547),
.B(n_4502),
.Y(n_4588)
);

XNOR2x1_ASAP7_75t_L g4589 ( 
.A(n_4543),
.B(n_4551),
.Y(n_4589)
);

HB1xp67_ASAP7_75t_L g4590 ( 
.A(n_4545),
.Y(n_4590)
);

INVx1_ASAP7_75t_SL g4591 ( 
.A(n_4560),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4561),
.Y(n_4592)
);

HB1xp67_ASAP7_75t_L g4593 ( 
.A(n_4534),
.Y(n_4593)
);

BUFx2_ASAP7_75t_L g4594 ( 
.A(n_4562),
.Y(n_4594)
);

AOI22xp5_ASAP7_75t_L g4595 ( 
.A1(n_4527),
.A2(n_4488),
.B1(n_4505),
.B2(n_4479),
.Y(n_4595)
);

OA22x2_ASAP7_75t_L g4596 ( 
.A1(n_4546),
.A2(n_4464),
.B1(n_4455),
.B2(n_4474),
.Y(n_4596)
);

OAI22xp5_ASAP7_75t_L g4597 ( 
.A1(n_4553),
.A2(n_4492),
.B1(n_4467),
.B2(n_4476),
.Y(n_4597)
);

HB1xp67_ASAP7_75t_L g4598 ( 
.A(n_4539),
.Y(n_4598)
);

XOR2x2_ASAP7_75t_L g4599 ( 
.A(n_4548),
.B(n_4463),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4544),
.Y(n_4600)
);

OA22x2_ASAP7_75t_L g4601 ( 
.A1(n_4563),
.A2(n_4458),
.B1(n_4501),
.B2(n_696),
.Y(n_4601)
);

INVx2_ASAP7_75t_SL g4602 ( 
.A(n_4540),
.Y(n_4602)
);

INVx2_ASAP7_75t_SL g4603 ( 
.A(n_4541),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4549),
.Y(n_4604)
);

INVxp33_ASAP7_75t_L g4605 ( 
.A(n_4552),
.Y(n_4605)
);

OAI22xp33_ASAP7_75t_L g4606 ( 
.A1(n_4557),
.A2(n_694),
.B1(n_695),
.B2(n_696),
.Y(n_4606)
);

XNOR2xp5_ASAP7_75t_L g4607 ( 
.A(n_4564),
.B(n_4558),
.Y(n_4607)
);

INVx2_ASAP7_75t_L g4608 ( 
.A(n_4554),
.Y(n_4608)
);

CKINVDCx5p33_ASAP7_75t_R g4609 ( 
.A(n_4540),
.Y(n_4609)
);

OA22x2_ASAP7_75t_L g4610 ( 
.A1(n_4528),
.A2(n_697),
.B1(n_698),
.B2(n_699),
.Y(n_4610)
);

XOR2x2_ASAP7_75t_L g4611 ( 
.A(n_4524),
.B(n_697),
.Y(n_4611)
);

AOI322xp5_ASAP7_75t_L g4612 ( 
.A1(n_4565),
.A2(n_698),
.A3(n_700),
.B1(n_701),
.B2(n_702),
.C1(n_703),
.C2(n_704),
.Y(n_4612)
);

OAI322xp33_ASAP7_75t_L g4613 ( 
.A1(n_4578),
.A2(n_701),
.A3(n_703),
.B1(n_704),
.B2(n_706),
.C1(n_707),
.C2(n_708),
.Y(n_4613)
);

INVxp67_ASAP7_75t_SL g4614 ( 
.A(n_4610),
.Y(n_4614)
);

INVx2_ASAP7_75t_L g4615 ( 
.A(n_4580),
.Y(n_4615)
);

AND2x4_ASAP7_75t_L g4616 ( 
.A(n_4567),
.B(n_706),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4590),
.Y(n_4617)
);

CKINVDCx20_ASAP7_75t_R g4618 ( 
.A(n_4594),
.Y(n_4618)
);

BUFx3_ASAP7_75t_L g4619 ( 
.A(n_4570),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4608),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4587),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4575),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4576),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4592),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4577),
.Y(n_4625)
);

HB1xp67_ASAP7_75t_L g4626 ( 
.A(n_4574),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4569),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4571),
.B(n_707),
.Y(n_4628)
);

OAI322xp33_ASAP7_75t_L g4629 ( 
.A1(n_4578),
.A2(n_709),
.A3(n_711),
.B1(n_712),
.B2(n_713),
.C1(n_714),
.C2(n_716),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4582),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4600),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4593),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4566),
.B(n_709),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4572),
.Y(n_4634)
);

INVxp67_ASAP7_75t_L g4635 ( 
.A(n_4604),
.Y(n_4635)
);

HB1xp67_ASAP7_75t_L g4636 ( 
.A(n_4566),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4598),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4586),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4584),
.B(n_713),
.Y(n_4639)
);

AOI322xp5_ASAP7_75t_L g4640 ( 
.A1(n_4602),
.A2(n_4603),
.A3(n_4591),
.B1(n_4595),
.B2(n_4609),
.C1(n_4589),
.C2(n_4585),
.Y(n_4640)
);

CKINVDCx6p67_ASAP7_75t_R g4641 ( 
.A(n_4591),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4568),
.Y(n_4642)
);

AND4x1_ASAP7_75t_L g4643 ( 
.A(n_4633),
.B(n_4595),
.C(n_4573),
.D(n_4579),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4615),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4617),
.Y(n_4645)
);

AOI22xp5_ASAP7_75t_SL g4646 ( 
.A1(n_4614),
.A2(n_4601),
.B1(n_4596),
.B2(n_4607),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4621),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4620),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4622),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_SL g4650 ( 
.A(n_4616),
.Y(n_4650)
);

OA22x2_ASAP7_75t_L g4651 ( 
.A1(n_4614),
.A2(n_4635),
.B1(n_4636),
.B2(n_4638),
.Y(n_4651)
);

AO22x1_ASAP7_75t_L g4652 ( 
.A1(n_4628),
.A2(n_4605),
.B1(n_4584),
.B2(n_4597),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4633),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4619),
.Y(n_4654)
);

AOI22xp5_ASAP7_75t_L g4655 ( 
.A1(n_4618),
.A2(n_4601),
.B1(n_4596),
.B2(n_4571),
.Y(n_4655)
);

INVxp67_ASAP7_75t_L g4656 ( 
.A(n_4639),
.Y(n_4656)
);

AOI22xp5_ASAP7_75t_L g4657 ( 
.A1(n_4635),
.A2(n_4581),
.B1(n_4597),
.B2(n_4583),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_4641),
.B(n_4588),
.Y(n_4658)
);

AOI22x1_ASAP7_75t_L g4659 ( 
.A1(n_4637),
.A2(n_4611),
.B1(n_4581),
.B2(n_4610),
.Y(n_4659)
);

OA22x2_ASAP7_75t_SL g4660 ( 
.A1(n_4632),
.A2(n_4583),
.B1(n_4599),
.B2(n_4606),
.Y(n_4660)
);

AOI22xp33_ASAP7_75t_L g4661 ( 
.A1(n_4624),
.A2(n_840),
.B1(n_718),
.B2(n_719),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4626),
.Y(n_4662)
);

AOI22xp5_ASAP7_75t_L g4663 ( 
.A1(n_4639),
.A2(n_717),
.B1(n_718),
.B2(n_720),
.Y(n_4663)
);

AOI31xp33_ASAP7_75t_L g4664 ( 
.A1(n_4640),
.A2(n_717),
.A3(n_721),
.B(n_722),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4630),
.Y(n_4665)
);

AOI221xp5_ASAP7_75t_L g4666 ( 
.A1(n_4613),
.A2(n_722),
.B1(n_723),
.B2(n_724),
.C(n_725),
.Y(n_4666)
);

OAI22xp33_ASAP7_75t_L g4667 ( 
.A1(n_4655),
.A2(n_4631),
.B1(n_4625),
.B2(n_4642),
.Y(n_4667)
);

INVx2_ASAP7_75t_L g4668 ( 
.A(n_4654),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4648),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4662),
.Y(n_4670)
);

AOI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4657),
.A2(n_4658),
.B1(n_4652),
.B2(n_4656),
.Y(n_4671)
);

AOI22xp5_ASAP7_75t_L g4672 ( 
.A1(n_4651),
.A2(n_4616),
.B1(n_4623),
.B2(n_4627),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4644),
.Y(n_4673)
);

OAI22xp5_ASAP7_75t_L g4674 ( 
.A1(n_4659),
.A2(n_4634),
.B1(n_4629),
.B2(n_4612),
.Y(n_4674)
);

O2A1O1Ixp5_ASAP7_75t_SL g4675 ( 
.A1(n_4645),
.A2(n_724),
.B(n_725),
.C(n_726),
.Y(n_4675)
);

AOI311xp33_ASAP7_75t_L g4676 ( 
.A1(n_4660),
.A2(n_727),
.A3(n_728),
.B(n_729),
.C(n_730),
.Y(n_4676)
);

AOI22xp33_ASAP7_75t_SL g4677 ( 
.A1(n_4646),
.A2(n_730),
.B1(n_731),
.B2(n_732),
.Y(n_4677)
);

AOI22xp33_ASAP7_75t_SL g4678 ( 
.A1(n_4649),
.A2(n_4643),
.B1(n_4653),
.B2(n_4647),
.Y(n_4678)
);

AOI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4650),
.A2(n_732),
.B1(n_733),
.B2(n_735),
.Y(n_4679)
);

INVxp67_ASAP7_75t_L g4680 ( 
.A(n_4664),
.Y(n_4680)
);

A2O1A1Ixp33_ASAP7_75t_SL g4681 ( 
.A1(n_4665),
.A2(n_733),
.B(n_735),
.C(n_737),
.Y(n_4681)
);

AO22x2_ASAP7_75t_L g4682 ( 
.A1(n_4643),
.A2(n_737),
.B1(n_738),
.B2(n_739),
.Y(n_4682)
);

O2A1O1Ixp33_ASAP7_75t_SL g4683 ( 
.A1(n_4666),
.A2(n_739),
.B(n_740),
.C(n_741),
.Y(n_4683)
);

A2O1A1Ixp33_ASAP7_75t_SL g4684 ( 
.A1(n_4663),
.A2(n_741),
.B(n_742),
.C(n_743),
.Y(n_4684)
);

HB1xp67_ASAP7_75t_L g4685 ( 
.A(n_4661),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4648),
.Y(n_4686)
);

OA22x2_ASAP7_75t_L g4687 ( 
.A1(n_4671),
.A2(n_839),
.B1(n_743),
.B2(n_744),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4668),
.Y(n_4688)
);

NOR4xp25_ASAP7_75t_L g4689 ( 
.A(n_4676),
.B(n_742),
.C(n_745),
.D(n_746),
.Y(n_4689)
);

NOR2x1_ASAP7_75t_L g4690 ( 
.A(n_4667),
.B(n_745),
.Y(n_4690)
);

AO22x2_ASAP7_75t_L g4691 ( 
.A1(n_4674),
.A2(n_746),
.B1(n_748),
.B2(n_749),
.Y(n_4691)
);

INVxp67_ASAP7_75t_SL g4692 ( 
.A(n_4679),
.Y(n_4692)
);

AO22x2_ASAP7_75t_L g4693 ( 
.A1(n_4680),
.A2(n_748),
.B1(n_749),
.B2(n_750),
.Y(n_4693)
);

AOI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4677),
.A2(n_751),
.B1(n_752),
.B2(n_753),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4682),
.B(n_751),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4670),
.Y(n_4696)
);

NOR4xp25_ASAP7_75t_L g4697 ( 
.A(n_4669),
.B(n_752),
.C(n_754),
.D(n_755),
.Y(n_4697)
);

OA22x2_ASAP7_75t_L g4698 ( 
.A1(n_4672),
.A2(n_836),
.B1(n_755),
.B2(n_756),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_SL g4699 ( 
.A(n_4678),
.B(n_754),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4673),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4688),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4693),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4695),
.Y(n_4703)
);

AOI22xp5_ASAP7_75t_L g4704 ( 
.A1(n_4691),
.A2(n_4682),
.B1(n_4685),
.B2(n_4686),
.Y(n_4704)
);

AOI22xp5_ASAP7_75t_L g4705 ( 
.A1(n_4692),
.A2(n_4683),
.B1(n_4684),
.B2(n_4681),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4696),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4687),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4700),
.Y(n_4708)
);

INVxp67_ASAP7_75t_L g4709 ( 
.A(n_4690),
.Y(n_4709)
);

AOI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4699),
.A2(n_4675),
.B1(n_758),
.B2(n_759),
.Y(n_4710)
);

INVxp67_ASAP7_75t_L g4711 ( 
.A(n_4694),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4698),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4707),
.Y(n_4713)
);

AOI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4712),
.A2(n_4689),
.B1(n_4697),
.B2(n_760),
.Y(n_4714)
);

OAI22xp5_ASAP7_75t_L g4715 ( 
.A1(n_4705),
.A2(n_757),
.B1(n_759),
.B2(n_760),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4701),
.Y(n_4716)
);

HB1xp67_ASAP7_75t_L g4717 ( 
.A(n_4706),
.Y(n_4717)
);

AO22x2_ASAP7_75t_L g4718 ( 
.A1(n_4702),
.A2(n_761),
.B1(n_762),
.B2(n_763),
.Y(n_4718)
);

NOR2xp67_ASAP7_75t_L g4719 ( 
.A(n_4709),
.B(n_763),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4704),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4713),
.Y(n_4721)
);

AO22x2_ASAP7_75t_L g4722 ( 
.A1(n_4720),
.A2(n_4703),
.B1(n_4708),
.B2(n_4711),
.Y(n_4722)
);

HB1xp67_ASAP7_75t_L g4723 ( 
.A(n_4719),
.Y(n_4723)
);

AOI22xp5_ASAP7_75t_L g4724 ( 
.A1(n_4722),
.A2(n_4714),
.B1(n_4715),
.B2(n_4710),
.Y(n_4724)
);

AOI22xp33_ASAP7_75t_L g4725 ( 
.A1(n_4721),
.A2(n_4716),
.B1(n_4717),
.B2(n_4718),
.Y(n_4725)
);

OAI22x1_ASAP7_75t_L g4726 ( 
.A1(n_4723),
.A2(n_836),
.B1(n_765),
.B2(n_766),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4726),
.Y(n_4727)
);

AOI211xp5_ASAP7_75t_L g4728 ( 
.A1(n_4727),
.A2(n_4724),
.B(n_4725),
.C(n_766),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4728),
.Y(n_4729)
);

AOI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4729),
.A2(n_764),
.B1(n_765),
.B2(n_767),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4730),
.Y(n_4731)
);

AOI221xp5_ASAP7_75t_L g4732 ( 
.A1(n_4731),
.A2(n_768),
.B1(n_769),
.B2(n_770),
.C(n_771),
.Y(n_4732)
);

AOI211xp5_ASAP7_75t_L g4733 ( 
.A1(n_4732),
.A2(n_768),
.B(n_769),
.C(n_770),
.Y(n_4733)
);


endmodule