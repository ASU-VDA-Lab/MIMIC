module real_jpeg_27825_n_8 (n_5, n_4, n_0, n_54, n_1, n_51, n_2, n_6, n_50, n_7, n_55, n_53, n_3, n_49, n_52, n_8);

input n_5;
input n_4;
input n_0;
input n_54;
input n_1;
input n_51;
input n_2;
input n_6;
input n_50;
input n_7;
input n_55;
input n_53;
input n_3;
input n_49;
input n_52;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_0),
.B(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_1),
.B(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_4),
.B(n_19),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_17),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_15),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_12),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B(n_47),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_42),
.B(n_46),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_38),
.B(n_41),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B(n_37),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_32),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_40),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_49),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_50),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_51),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_52),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_53),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_54),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_55),
.Y(n_45)
);


endmodule