module fake_jpeg_4548_n_235 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_32),
.B(n_34),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_6),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_11),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_26),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_27),
.B1(n_25),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_22),
.B1(n_26),
.B2(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_60),
.B1(n_61),
.B2(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_62),
.Y(n_90)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_81),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_20),
.B1(n_23),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_27),
.B1(n_17),
.B2(n_23),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_63),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_31),
.B1(n_21),
.B2(n_20),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_82),
.B1(n_75),
.B2(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_35),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_29),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_77),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_23),
.B1(n_21),
.B2(n_2),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_5),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_79),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_5),
.B(n_12),
.C(n_10),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_6),
.B1(n_10),
.B2(n_7),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_36),
.B(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_0),
.C(n_1),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_58),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_62),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_70),
.B(n_86),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_54),
.B1(n_80),
.B2(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_73),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_113),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_2),
.A3(n_13),
.B1(n_79),
.B2(n_48),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_58),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_2),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_84),
.B1(n_56),
.B2(n_55),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_80),
.B(n_74),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_49),
.C(n_55),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_88),
.B1(n_75),
.B2(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_89),
.B1(n_88),
.B2(n_52),
.Y(n_121)
);

BUFx4f_ASAP7_75t_SL g118 ( 
.A(n_92),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_92),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_137),
.B1(n_140),
.B2(n_116),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_132),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_R g124 ( 
.A(n_96),
.B(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_104),
.B1(n_102),
.B2(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_63),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_135),
.Y(n_154)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_83),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_55),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_138),
.Y(n_149)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_63),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_146),
.B1(n_140),
.B2(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_145),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_158),
.B1(n_160),
.B2(n_165),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_97),
.B(n_110),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_163),
.B(n_164),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_145),
.C(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_121),
.C(n_100),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_105),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_93),
.B1(n_107),
.B2(n_108),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_93),
.B1(n_107),
.B2(n_108),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_131),
.B(n_126),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_96),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_117),
.B(n_111),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_133),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_181),
.C(n_188),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_154),
.A3(n_157),
.B1(n_147),
.B2(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_180),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_150),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_133),
.B(n_111),
.C(n_90),
.D(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_137),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_100),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_99),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_99),
.B1(n_94),
.B2(n_118),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_72),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_72),
.C(n_120),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_73),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_164),
.A3(n_156),
.B1(n_154),
.B2(n_147),
.C1(n_169),
.C2(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_171),
.B1(n_162),
.B2(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_158),
.B1(n_160),
.B2(n_149),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_170),
.C(n_169),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_155),
.B(n_167),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_155),
.B(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_205),
.A2(n_177),
.B1(n_172),
.B2(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_196),
.B1(n_203),
.B2(n_194),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_196),
.B(n_195),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_204),
.B(n_200),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_209),
.B1(n_206),
.B2(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_213),
.B1(n_202),
.B2(n_151),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_220),
.A2(n_215),
.B1(n_206),
.B2(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_193),
.C(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_213),
.C(n_166),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_223),
.A2(n_212),
.B1(n_218),
.B2(n_219),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.C(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_161),
.C(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_230),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_222),
.C(n_225),
.Y(n_230)
);

OA21x2_ASAP7_75t_SL g233 ( 
.A1(n_231),
.A2(n_201),
.B(n_226),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_232),
.Y(n_235)
);


endmodule