module real_jpeg_3170_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_32),
.B1(n_34),
.B2(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_3),
.A2(n_32),
.B1(n_39),
.B2(n_47),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.C(n_39),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_34),
.B1(n_61),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_58),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_6),
.B(n_26),
.C(n_48),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_39),
.B1(n_47),
.B2(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_6),
.B(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_6),
.B(n_72),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_39),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_54),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_39),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_11),
.A2(n_34),
.B1(n_52),
.B2(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_11),
.A2(n_24),
.B1(n_26),
.B2(n_52),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_66),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_18),
.B(n_66),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.C(n_55),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_19),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_19)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_42),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_21),
.A2(n_23),
.B1(n_30),
.B2(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_21),
.A2(n_30),
.B1(n_98),
.B2(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_22),
.A2(n_29),
.B(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_26),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_26),
.B(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_30),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_38),
.B1(n_59),
.B2(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_34),
.A2(n_61),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_39),
.B(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_43),
.B(n_55),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_44),
.A2(n_71),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_45),
.B(n_73),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_51),
.B(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_64),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_63),
.A2(n_100),
.B(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_75),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_134),
.B(n_138),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_115),
.B(n_133),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_109),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_104),
.C(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_127),
.B(n_132),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_122),
.B(n_126),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_125),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);


endmodule