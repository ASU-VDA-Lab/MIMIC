module fake_jpeg_25108_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_70),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_0),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_61),
.B1(n_66),
.B2(n_63),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_SL g77 ( 
.A(n_74),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_63),
.B1(n_67),
.B2(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_61),
.B1(n_55),
.B2(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_54),
.B(n_45),
.C(n_64),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_60),
.B1(n_57),
.B2(n_47),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_49),
.B(n_57),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_86),
.B1(n_1),
.B2(n_2),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_67),
.B1(n_53),
.B2(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_59),
.B1(n_65),
.B2(n_52),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_96),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_95),
.B1(n_81),
.B2(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_3),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_4),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_7),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_4),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_110),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_111),
.B1(n_9),
.B2(n_12),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_22),
.B(n_40),
.C(n_38),
.D(n_11),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_13),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_31),
.B(n_32),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_122),
.B(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_111),
.C(n_109),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_126),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_21),
.B(n_27),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_33),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_128),
.B(n_119),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_127),
.B(n_132),
.C(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_131),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_120),
.B(n_36),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_34),
.Y(n_140)
);


endmodule