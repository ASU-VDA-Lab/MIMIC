module real_aes_6352_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_528;
wire n_372;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_0), .A2(n_245), .B1(n_453), .B2(n_696), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_1), .A2(n_120), .B1(n_771), .B2(n_824), .Y(n_899) );
AOI22xp5_ASAP7_75t_SL g604 ( .A1(n_2), .A2(n_238), .B1(n_354), .B2(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_3), .A2(n_16), .B1(n_614), .B2(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_4), .A2(n_112), .B1(n_488), .B2(n_785), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_5), .A2(n_57), .B1(n_397), .B2(n_398), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_6), .Y(n_360) );
INVx1_ASAP7_75t_L g376 ( .A(n_7), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_8), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_9), .A2(n_131), .B1(n_508), .B2(n_675), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_10), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_11), .A2(n_138), .B1(n_742), .B2(n_776), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_12), .A2(n_148), .B1(n_422), .B2(n_423), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g721 ( .A1(n_13), .A2(n_128), .B1(n_217), .B2(n_435), .C1(n_488), .C2(n_540), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_14), .A2(n_226), .B1(n_418), .B2(n_769), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_15), .A2(n_220), .B1(n_771), .B2(n_773), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_17), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_18), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_19), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_20), .A2(n_168), .B1(n_502), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_21), .A2(n_76), .B1(n_696), .B2(n_697), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_22), .A2(n_103), .B1(n_462), .B2(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_23), .B(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_24), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_25), .B(n_666), .Y(n_665) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_26), .A2(n_90), .B1(n_308), .B2(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g849 ( .A(n_26), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_27), .A2(n_162), .B1(n_448), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_28), .A2(n_194), .B1(n_531), .B2(n_675), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_29), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_30), .A2(n_210), .B1(n_344), .B2(n_614), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_31), .A2(n_157), .B1(n_419), .B2(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_32), .A2(n_284), .B1(n_422), .B2(n_582), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_33), .A2(n_259), .B1(n_409), .B2(n_410), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_34), .B(n_390), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_35), .A2(n_515), .B1(n_552), .B2(n_553), .Y(n_514) );
INVx1_ASAP7_75t_L g552 ( .A(n_35), .Y(n_552) );
INVx1_ASAP7_75t_L g402 ( .A(n_36), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_37), .Y(n_816) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_38), .A2(n_176), .B1(n_398), .B2(n_668), .Y(n_667) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_39), .A2(n_94), .B1(n_308), .B2(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g850 ( .A(n_39), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_40), .A2(n_135), .B1(n_319), .B2(n_323), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_41), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_42), .A2(n_267), .B1(n_394), .B2(n_445), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_43), .A2(n_163), .B1(n_419), .B2(n_528), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_44), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_45), .A2(n_110), .B1(n_457), .B2(n_459), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_46), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_47), .A2(n_93), .B1(n_459), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_48), .A2(n_72), .B1(n_453), .B2(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_49), .B(n_544), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_50), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_51), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_52), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_53), .A2(n_160), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_54), .A2(n_853), .B1(n_854), .B2(n_868), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_54), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_55), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_56), .A2(n_115), .B1(n_459), .B2(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g866 ( .A1(n_58), .A2(n_188), .B1(n_264), .B2(n_344), .C1(n_486), .C2(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_59), .A2(n_61), .B1(n_414), .B2(n_466), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_60), .A2(n_77), .B1(n_415), .B2(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_62), .Y(n_519) );
AOI22xp5_ASAP7_75t_SL g601 ( .A1(n_63), .A2(n_161), .B1(n_499), .B2(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_64), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_64), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_65), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_66), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_67), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_68), .A2(n_277), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_69), .A2(n_150), .B1(n_450), .B2(n_614), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_70), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_71), .A2(n_192), .B1(n_672), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_73), .A2(n_186), .B1(n_422), .B2(n_528), .Y(n_864) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_74), .B(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_75), .A2(n_196), .B1(n_422), .B2(n_505), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_78), .A2(n_167), .B1(n_531), .B2(n_584), .Y(n_778) );
AOI22xp5_ASAP7_75t_SL g599 ( .A1(n_79), .A2(n_143), .B1(n_410), .B2(n_600), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_80), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_81), .A2(n_224), .B1(n_395), .B2(n_445), .Y(n_615) );
AO22x2_ASAP7_75t_L g470 ( .A1(n_82), .A2(n_471), .B1(n_509), .B2(n_510), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_82), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_83), .A2(n_235), .B1(n_501), .B2(n_502), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_84), .Y(n_535) );
INVx1_ASAP7_75t_L g637 ( .A(n_85), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g807 ( .A1(n_86), .A2(n_483), .B(n_808), .C(n_813), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_87), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_88), .A2(n_149), .B1(n_582), .B2(n_675), .Y(n_792) );
INVx1_ASAP7_75t_L g424 ( .A(n_89), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_91), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_92), .Y(n_684) );
INVx1_ASAP7_75t_L g633 ( .A(n_95), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_96), .A2(n_202), .B1(n_350), .B2(n_460), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_97), .Y(n_541) );
AND2x2_ASAP7_75t_L g293 ( .A(n_98), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g743 ( .A(n_99), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_100), .A2(n_152), .B1(n_579), .B2(n_582), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_101), .A2(n_136), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_102), .A2(n_199), .B1(n_418), .B2(n_422), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_104), .A2(n_203), .B1(n_423), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_105), .A2(n_140), .B1(n_466), .B2(n_579), .Y(n_646) );
INVx1_ASAP7_75t_L g290 ( .A(n_106), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_107), .A2(n_147), .B1(n_319), .B2(n_344), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_108), .A2(n_169), .B1(n_531), .B2(n_593), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_109), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g328 ( .A(n_111), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_113), .A2(n_244), .B1(n_414), .B2(n_508), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_114), .A2(n_156), .B1(n_668), .B2(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_116), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_117), .A2(n_219), .B1(n_344), .B2(n_614), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_118), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_119), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_121), .B(n_390), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_122), .A2(n_257), .B1(n_579), .B2(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_123), .A2(n_178), .B1(n_507), .B2(n_675), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_124), .A2(n_208), .B1(n_414), .B2(n_589), .Y(n_588) );
XNOR2xp5_ASAP7_75t_L g430 ( .A(n_125), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_126), .B(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_127), .Y(n_537) );
INVx1_ASAP7_75t_L g733 ( .A(n_129), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_130), .A2(n_246), .B1(n_589), .B2(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g380 ( .A(n_132), .Y(n_380) );
AOI22xp5_ASAP7_75t_SL g627 ( .A1(n_133), .A2(n_628), .B1(n_654), .B2(n_655), .Y(n_627) );
INVx1_ASAP7_75t_L g655 ( .A(n_133), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_134), .A2(n_236), .B1(n_460), .B2(n_593), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_137), .A2(n_181), .B1(n_323), .B2(n_488), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_139), .A2(n_213), .B1(n_447), .B2(n_448), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_141), .A2(n_225), .B1(n_579), .B2(n_651), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_142), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_144), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_145), .B(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g294 ( .A(n_146), .Y(n_294) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_151), .A2(n_222), .B1(n_438), .B2(n_439), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_153), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_154), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_155), .A2(n_206), .B1(n_459), .B2(n_592), .Y(n_698) );
AND2x6_ASAP7_75t_L g289 ( .A(n_158), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_158), .Y(n_843) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_159), .A2(n_232), .B1(n_308), .B2(n_312), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_164), .A2(n_255), .B1(n_418), .B2(n_504), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g805 ( .A(n_165), .Y(n_805) );
INVx1_ASAP7_75t_L g631 ( .A(n_166), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_170), .A2(n_200), .B1(n_409), .B2(n_600), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_171), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_172), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_173), .A2(n_261), .B1(n_418), .B2(n_419), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_174), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_175), .B(n_571), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_177), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_179), .A2(n_195), .B1(n_453), .B2(n_593), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_180), .Y(n_797) );
INVx1_ASAP7_75t_L g643 ( .A(n_182), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_183), .A2(n_205), .B1(n_531), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_184), .A2(n_260), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_185), .A2(n_252), .B1(n_582), .B2(n_675), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_187), .Y(n_677) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_189), .A2(n_248), .B1(n_308), .B2(n_309), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_190), .A2(n_269), .B1(n_488), .B2(n_668), .Y(n_734) );
INVx1_ASAP7_75t_L g638 ( .A(n_191), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_193), .A2(n_253), .B1(n_485), .B2(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g303 ( .A(n_197), .Y(n_303) );
INVx1_ASAP7_75t_L g832 ( .A(n_198), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_201), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_204), .A2(n_278), .B1(n_405), .B2(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g373 ( .A(n_207), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_209), .B(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_211), .A2(n_254), .B1(n_499), .B2(n_600), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_212), .A2(n_231), .B1(n_462), .B2(n_464), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_214), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_215), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g764 ( .A(n_216), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_218), .A2(n_251), .B1(n_460), .B2(n_501), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_221), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_223), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_227), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_228), .A2(n_237), .B1(n_414), .B2(n_415), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_229), .Y(n_573) );
INVx1_ASAP7_75t_L g760 ( .A(n_230), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_232), .B(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_233), .B(n_394), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_234), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_239), .A2(n_281), .B1(n_584), .B2(n_585), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_240), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_241), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_242), .A2(n_258), .B1(n_394), .B2(n_811), .Y(n_860) );
INVx1_ASAP7_75t_L g641 ( .A(n_243), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_247), .A2(n_263), .B1(n_592), .B2(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g846 ( .A(n_248), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_249), .A2(n_250), .B1(n_768), .B2(n_769), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_256), .Y(n_692) );
OA22x2_ASAP7_75t_L g555 ( .A1(n_262), .A2(n_556), .B1(n_557), .B2(n_595), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_262), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_265), .Y(n_883) );
INVx1_ASAP7_75t_L g308 ( .A(n_266), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_268), .Y(n_436) );
INVx1_ASAP7_75t_L g757 ( .A(n_270), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_271), .Y(n_892) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_272), .A2(n_287), .B(n_295), .C(n_851), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_273), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_274), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_275), .A2(n_285), .B1(n_344), .B2(n_439), .Y(n_761) );
INVx1_ASAP7_75t_L g756 ( .A(n_276), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_279), .Y(n_783) );
INVx1_ASAP7_75t_L g763 ( .A(n_280), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_282), .A2(n_681), .B1(n_704), .B2(n_705), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_282), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_283), .Y(n_561) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_290), .Y(n_842) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_291), .A2(n_841), .B(n_877), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_620), .B1(n_836), .B2(n_837), .C(n_838), .Y(n_295) );
INVx1_ASAP7_75t_L g837 ( .A(n_296), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_381), .B2(n_382), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
XNOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_380), .Y(n_299) );
AND3x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_347), .C(n_364), .Y(n_300) );
NOR3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_327), .C(n_336), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_318), .Y(n_302) );
INVx2_ASAP7_75t_L g476 ( .A(n_304), .Y(n_476) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_304), .Y(n_632) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_313), .Y(n_304) );
INVx2_ASAP7_75t_L g379 ( .A(n_305), .Y(n_379) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_311), .Y(n_305) );
AND2x2_ASAP7_75t_L g331 ( .A(n_306), .B(n_311), .Y(n_331) );
AND2x2_ASAP7_75t_L g351 ( .A(n_306), .B(n_335), .Y(n_351) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g322 ( .A(n_307), .B(n_317), .Y(n_322) );
AND2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_311), .Y(n_326) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_310), .Y(n_312) );
INVx2_ASAP7_75t_L g335 ( .A(n_311), .Y(n_335) );
INVx1_ASAP7_75t_L g400 ( .A(n_311), .Y(n_400) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_314), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g350 ( .A(n_314), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g392 ( .A(n_314), .B(n_379), .Y(n_392) );
AND2x6_ASAP7_75t_L g395 ( .A(n_314), .B(n_331), .Y(n_395) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g321 ( .A(n_315), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_315), .Y(n_325) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_315), .B(n_317), .Y(n_356) );
AND2x2_ASAP7_75t_L g340 ( .A(n_316), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g371 ( .A(n_317), .B(n_325), .Y(n_371) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_319), .Y(n_405) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_319), .Y(n_439) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_319), .Y(n_488) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g346 ( .A(n_321), .B(n_335), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_322), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g345 ( .A(n_322), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g398 ( .A(n_322), .B(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_SL g406 ( .A(n_323), .Y(n_406) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_323), .Y(n_450) );
BUFx3_ASAP7_75t_L g668 ( .A(n_323), .Y(n_668) );
BUFx2_ASAP7_75t_SL g785 ( .A(n_323), .Y(n_785) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g496 ( .A(n_324), .Y(n_496) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x6_ASAP7_75t_L g339 ( .A(n_326), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g495 ( .A(n_326), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B1(n_332), .B2(n_333), .Y(n_327) );
INVx2_ASAP7_75t_L g563 ( .A(n_329), .Y(n_563) );
OA211x2_ASAP7_75t_L g717 ( .A1(n_329), .A2(n_718), .B(n_719), .C(n_720), .Y(n_717) );
BUFx3_ASAP7_75t_L g758 ( .A(n_329), .Y(n_758) );
OAI22xp5_ASAP7_75t_SL g882 ( .A1(n_329), .A2(n_632), .B1(n_883), .B2(n_884), .Y(n_882) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g479 ( .A(n_330), .Y(n_479) );
AND2x4_ASAP7_75t_L g362 ( .A(n_331), .B(n_340), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_331), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_331), .B(n_371), .Y(n_412) );
INVx4_ASAP7_75t_L g492 ( .A(n_333), .Y(n_492) );
BUFx3_ASAP7_75t_L g548 ( .A(n_333), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_333), .A2(n_575), .B1(n_763), .B2(n_764), .Y(n_762) );
AND2x2_ASAP7_75t_L g354 ( .A(n_334), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_342), .B2(n_343), .Y(n_336) );
OAI222xp33_ASAP7_75t_L g885 ( .A1(n_338), .A2(n_886), .B1(n_888), .B2(n_889), .C1(n_890), .C2(n_892), .Y(n_885) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_339), .Y(n_435) );
BUFx3_ASAP7_75t_L g483 ( .A(n_339), .Y(n_483) );
INVx4_ASAP7_75t_L g566 ( .A(n_339), .Y(n_566) );
INVx2_ASAP7_75t_L g610 ( .A(n_339), .Y(n_610) );
AND2x2_ASAP7_75t_L g359 ( .A(n_340), .B(n_351), .Y(n_359) );
AND2x6_ASAP7_75t_L g378 ( .A(n_340), .B(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g438 ( .A(n_343), .Y(n_438) );
INVx4_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_345), .Y(n_397) );
BUFx2_ASAP7_75t_L g485 ( .A(n_345), .Y(n_485) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_345), .Y(n_540) );
BUFx4f_ASAP7_75t_SL g788 ( .A(n_345), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_357), .Y(n_347) );
OAI21xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_352), .B(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g697 ( .A(n_349), .Y(n_697) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
BUFx3_ASAP7_75t_L g505 ( .A(n_350), .Y(n_505) );
BUFx3_ASAP7_75t_L g528 ( .A(n_350), .Y(n_528) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_350), .Y(n_742) );
AND2x4_ASAP7_75t_L g368 ( .A(n_351), .B(n_355), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_351), .B(n_371), .Y(n_374) );
AND2x2_ASAP7_75t_L g420 ( .A(n_351), .B(n_371), .Y(n_420) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x6_ASAP7_75t_L g416 ( .A(n_356), .B(n_400), .Y(n_416) );
OAI22xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_360), .B1(n_361), .B2(n_363), .Y(n_357) );
INVx3_ASAP7_75t_L g422 ( .A(n_358), .Y(n_422) );
INVx3_ASAP7_75t_L g504 ( .A(n_358), .Y(n_504) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_359), .Y(n_463) );
BUFx2_ASAP7_75t_SL g602 ( .A(n_359), .Y(n_602) );
INVx2_ASAP7_75t_L g409 ( .A(n_361), .Y(n_409) );
INVx3_ASAP7_75t_L g531 ( .A(n_361), .Y(n_531) );
INVx2_ASAP7_75t_L g701 ( .A(n_361), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_361), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_825) );
INVx6_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g453 ( .A(n_362), .Y(n_453) );
BUFx3_ASAP7_75t_L g499 ( .A(n_362), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_372), .C(n_375), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_369), .B2(n_370), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g423 ( .A(n_368), .Y(n_423) );
BUFx3_ASAP7_75t_L g468 ( .A(n_368), .Y(n_468) );
BUFx3_ASAP7_75t_L g508 ( .A(n_368), .Y(n_508) );
BUFx3_ASAP7_75t_L g582 ( .A(n_368), .Y(n_582) );
BUFx3_ASAP7_75t_L g605 ( .A(n_368), .Y(n_605) );
BUFx2_ASAP7_75t_SL g769 ( .A(n_368), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g834 ( .A(n_374), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx5_ASAP7_75t_SL g418 ( .A(n_377), .Y(n_418) );
INVx4_ASAP7_75t_L g464 ( .A(n_377), .Y(n_464) );
INVx2_ASAP7_75t_SL g507 ( .A(n_377), .Y(n_507) );
INVx2_ASAP7_75t_L g648 ( .A(n_377), .Y(n_648) );
INVx11_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx11_ASAP7_75t_L g518 ( .A(n_378), .Y(n_518) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_511), .B1(n_618), .B2(n_619), .Y(n_382) );
INVx1_ASAP7_75t_L g619 ( .A(n_383), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_425), .B2(n_426), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
XOR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_424), .Y(n_385) );
NAND4xp75_ASAP7_75t_SL g386 ( .A(n_387), .B(n_407), .C(n_417), .D(n_421), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g387 ( .A(n_388), .B(n_401), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .C(n_396), .Y(n_388) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx5_ASAP7_75t_L g445 ( .A(n_391), .Y(n_445) );
INVx2_ASAP7_75t_L g666 ( .A(n_391), .Y(n_666) );
INVx2_ASAP7_75t_L g811 ( .A(n_391), .Y(n_811) );
INVx4_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
BUFx4f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g729 ( .A(n_395), .Y(n_729) );
INVx1_ASAP7_75t_L g815 ( .A(n_397), .Y(n_815) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_397), .Y(n_887) );
BUFx2_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
BUFx3_ASAP7_75t_L g614 ( .A(n_398), .Y(n_614) );
INVx1_ASAP7_75t_L g688 ( .A(n_398), .Y(n_688) );
BUFx2_ASAP7_75t_L g862 ( .A(n_398), .Y(n_862) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_404), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_403), .A2(n_661), .B(n_662), .Y(n_660) );
OAI222xp33_ASAP7_75t_L g689 ( .A1(n_403), .A2(n_539), .B1(n_543), .B2(n_690), .C1(n_691), .C2(n_692), .Y(n_689) );
OAI21xp5_ASAP7_75t_SL g732 ( .A1(n_403), .A2(n_733), .B(n_734), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_403), .A2(n_783), .B(n_784), .Y(n_782) );
BUFx3_ASAP7_75t_L g544 ( .A(n_405), .Y(n_544) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_413), .Y(n_407) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx4_ASAP7_75t_L g458 ( .A(n_411), .Y(n_458) );
INVx2_ASAP7_75t_L g501 ( .A(n_411), .Y(n_501) );
INVx5_ASAP7_75t_L g593 ( .A(n_411), .Y(n_593) );
INVx1_ASAP7_75t_L g672 ( .A(n_411), .Y(n_672) );
INVx8_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g651 ( .A(n_414), .Y(n_651) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx6_ASAP7_75t_SL g460 ( .A(n_416), .Y(n_460) );
INVx1_ASAP7_75t_L g594 ( .A(n_416), .Y(n_594) );
INVx1_ASAP7_75t_SL g824 ( .A(n_416), .Y(n_824) );
INVx1_ASAP7_75t_L g777 ( .A(n_418), .Y(n_777) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
BUFx2_ASAP7_75t_L g532 ( .A(n_419), .Y(n_532) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g581 ( .A(n_420), .Y(n_581) );
BUFx3_ASAP7_75t_L g675 ( .A(n_420), .Y(n_675) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AO22x1_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_469), .B2(n_470), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND4xp75_ASAP7_75t_SL g431 ( .A(n_432), .B(n_451), .C(n_461), .D(n_465), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g432 ( .A(n_433), .B(n_440), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_436), .B(n_437), .Y(n_433) );
OAI222xp33_ASAP7_75t_L g538 ( .A1(n_434), .A2(n_539), .B1(n_541), .B2(n_542), .C1(n_543), .C2(n_545), .Y(n_538) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g636 ( .A(n_435), .Y(n_636) );
INVx1_ASAP7_75t_L g568 ( .A(n_438), .Y(n_568) );
BUFx4f_ASAP7_75t_L g891 ( .A(n_439), .Y(n_891) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .C(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g586 ( .A(n_453), .Y(n_586) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g772 ( .A(n_458), .Y(n_772) );
BUFx4f_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
BUFx2_ASAP7_75t_L g773 ( .A(n_460), .Y(n_773) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_463), .Y(n_584) );
BUFx3_ASAP7_75t_L g696 ( .A(n_463), .Y(n_696) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI221xp5_ASAP7_75t_SL g517 ( .A1(n_467), .A2(n_518), .B1(n_519), .B2(n_520), .C(n_521), .Y(n_517) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g509 ( .A(n_471), .Y(n_509) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_472), .B(n_497), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .C(n_489), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_477), .B2(n_478), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_475), .A2(n_562), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_683) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g536 ( .A(n_476), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_478), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_534) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g634 ( .A(n_479), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_484), .Y(n_480) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g817 ( .A(n_486), .Y(n_817) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx4f_ASAP7_75t_SL g571 ( .A(n_488), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_493), .B2(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_SL g642 ( .A(n_492), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_494), .Y(n_551) );
BUFx2_ASAP7_75t_L g575 ( .A(n_494), .Y(n_575) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
AND4x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .C(n_503), .D(n_506), .Y(n_497) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_501), .Y(n_522) );
INVx1_ASAP7_75t_L g590 ( .A(n_507), .Y(n_590) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_512), .Y(n_618) );
XOR2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_554), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
AND2x2_ASAP7_75t_SL g515 ( .A(n_516), .B(n_533), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
INVx3_ASAP7_75t_L g600 ( .A(n_518), .Y(n_600) );
OAI221xp5_ASAP7_75t_SL g523 ( .A1(n_524), .A2(n_525), .B1(n_526), .B2(n_529), .C(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .C(n_546), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_536), .A2(n_560), .B1(n_561), .B2(n_562), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_536), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_548), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
OAI22xp5_ASAP7_75t_SL g893 ( .A1(n_548), .A2(n_550), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_596), .B1(n_597), .B2(n_617), .Y(n_554) );
INVx1_ASAP7_75t_L g617 ( .A(n_555), .Y(n_617) );
INVx1_ASAP7_75t_L g595 ( .A(n_557), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_576), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .C(n_572), .Y(n_558) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_562), .A2(n_809), .B(n_810), .C(n_812), .Y(n_808) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B1(n_568), .B2(n_569), .C(n_570), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx4_ASAP7_75t_L g867 ( .A(n_566), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_568), .A2(n_636), .B1(n_637), .B2(n_638), .C(n_639), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_575), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_640) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_577), .B(n_587), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx4f_ASAP7_75t_SL g768 ( .A(n_581), .Y(n_768) );
BUFx2_ASAP7_75t_L g703 ( .A(n_582), .Y(n_703) );
INVx1_ASAP7_75t_SL g831 ( .A(n_584), .Y(n_831) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_593), .Y(n_653) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
XOR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_616), .Y(n_597) );
NAND4xp75_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .C(n_603), .D(n_607), .Y(n_598) );
INVx1_ASAP7_75t_L g827 ( .A(n_600), .Y(n_827) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g836 ( .A(n_620), .Y(n_836) );
AOI22xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_801), .B1(n_802), .B2(n_835), .Y(n_620) );
INVx1_ASAP7_75t_L g835 ( .A(n_621), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_706), .B1(n_799), .B2(n_800), .Y(n_621) );
INVx1_ASAP7_75t_L g799 ( .A(n_622), .Y(n_799) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B1(n_679), .B2(n_680), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
OA22x2_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_656), .B1(n_657), .B2(n_678), .Y(n_626) );
INVx1_ASAP7_75t_L g678 ( .A(n_627), .Y(n_678) );
INVx2_ASAP7_75t_SL g654 ( .A(n_628), .Y(n_654) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_644), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_635), .C(n_640), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
OAI21xp33_ASAP7_75t_SL g759 ( .A1(n_636), .A2(n_760), .B(n_761), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_649), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx4_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
XOR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_677), .Y(n_657) );
NAND3x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_669), .C(n_673), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .C(n_667), .Y(n_663) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g705 ( .A(n_681), .Y(n_705) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_693), .Y(n_681) );
NOR2xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_689), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_699), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g800 ( .A(n_706), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_746), .B2(n_747), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_723), .B1(n_744), .B2(n_745), .Y(n_708) );
INVx2_ASAP7_75t_SL g744 ( .A(n_709), .Y(n_744) );
XOR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_722), .Y(n_709) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .C(n_717), .D(n_721), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_SL g745 ( .A(n_723), .Y(n_745) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
XOR2x2_ASAP7_75t_SL g724 ( .A(n_725), .B(n_743), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g725 ( .A(n_726), .B(n_735), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_732), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .C(n_731), .Y(n_727) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx4_ASAP7_75t_L g822 ( .A(n_742), .Y(n_822) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AO22x1_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_779), .B2(n_798), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_765), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_759), .C(n_762), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_774), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
INVx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_778), .Y(n_774) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_SL g798 ( .A(n_779), .Y(n_798) );
XOR2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_797), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_781), .B(n_790), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_786), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
XNOR2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_818), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_813) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_825), .C(n_829), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_823), .Y(n_819) );
INVx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_829) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
OR2x2_ASAP7_75t_SL g905 ( .A(n_840), .B(n_845), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_841), .Y(n_871) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_842), .B(n_874), .Y(n_877) );
CKINVDCx16_ASAP7_75t_R g874 ( .A(n_843), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
OAI322xp33_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_869), .A3(n_872), .B1(n_875), .B2(n_878), .C1(n_879), .C2(n_903), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_854), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND4xp75_ASAP7_75t_L g855 ( .A(n_856), .B(n_859), .C(n_863), .D(n_866), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
AND2x2_ASAP7_75t_SL g859 ( .A(n_860), .B(n_861), .Y(n_859) );
AND2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
CKINVDCx16_ASAP7_75t_R g875 ( .A(n_876), .Y(n_875) );
XNOR2x2_ASAP7_75t_L g879 ( .A(n_878), .B(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_896), .Y(n_880) );
NOR3xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .C(n_893), .Y(n_881) );
INVx2_ASAP7_75t_SL g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_904), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_905), .Y(n_904) );
endmodule