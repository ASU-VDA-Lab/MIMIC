module fake_jpeg_5608_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_30),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_15),
.B1(n_26),
.B2(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_63),
.B1(n_19),
.B2(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_16),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_75),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_39),
.B(n_37),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_43),
.B(n_52),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_18),
.B1(n_34),
.B2(n_25),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_34),
.B1(n_49),
.B2(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_80),
.B1(n_51),
.B2(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_87),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_64),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_16),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_106),
.B1(n_67),
.B2(n_85),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_94),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_100),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_98),
.B(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_112),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_35),
.C(n_47),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_76),
.C(n_82),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_113),
.B1(n_66),
.B2(n_75),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_21),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_80),
.B(n_83),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_116),
.B(n_128),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_97),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_116),
.C(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_135),
.B1(n_139),
.B2(n_103),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_65),
.B(n_45),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_108),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_81),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_32),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_86),
.B(n_82),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_65),
.B1(n_42),
.B2(n_68),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_131),
.B1(n_92),
.B2(n_68),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_87),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_67),
.B(n_73),
.C(n_47),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_153),
.C(n_163),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_138),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_144),
.B1(n_119),
.B2(n_122),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_111),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_96),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_164),
.Y(n_172)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_150),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_72),
.B1(n_106),
.B2(n_92),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_95),
.B1(n_103),
.B2(n_110),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_161),
.B1(n_139),
.B2(n_121),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_95),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_72),
.B1(n_26),
.B2(n_24),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_16),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_158),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_115),
.B(n_107),
.C(n_47),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_114),
.B(n_131),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_121),
.B1(n_123),
.B2(n_117),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_32),
.C(n_33),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_165),
.B1(n_156),
.B2(n_161),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_171),
.B(n_187),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_119),
.B1(n_122),
.B2(n_134),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_180),
.B(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_183),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_176),
.C(n_166),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NAND4xp25_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_134),
.C(n_126),
.D(n_32),
.Y(n_182)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_199),
.B1(n_200),
.B2(n_185),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_165),
.B1(n_154),
.B2(n_151),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_183),
.A2(n_151),
.B1(n_125),
.B2(n_162),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_170),
.B1(n_33),
.B2(n_27),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_151),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_180),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_190),
.B1(n_171),
.B2(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_137),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_215),
.C(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_126),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_32),
.C(n_134),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_196),
.B(n_191),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_231),
.B(n_233),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_176),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_186),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_170),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_33),
.C(n_31),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_195),
.B1(n_192),
.B2(n_200),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_193),
.B(n_17),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_234),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_210),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_230),
.B(n_197),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_240),
.B1(n_242),
.B2(n_248),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_210),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_235),
.B1(n_231),
.B2(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_211),
.B1(n_212),
.B2(n_192),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_245),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_202),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_224),
.B1(n_218),
.B2(n_209),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_195),
.B1(n_203),
.B2(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_27),
.B1(n_24),
.B2(n_102),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_204),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_253),
.C(n_17),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_204),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_0),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_96),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_256),
.B(n_263),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_235),
.B(n_216),
.C(n_29),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_10),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_102),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_260),
.B(n_265),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_256),
.B1(n_263),
.B2(n_266),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_246),
.C(n_258),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_251),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_239),
.A2(n_23),
.B1(n_30),
.B2(n_8),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_10),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_0),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_276),
.C(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_274),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_281),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_246),
.B1(n_244),
.B2(n_10),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_262),
.Y(n_277)
);

NAND5xp2_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_0),
.C(n_1),
.D(n_2),
.E(n_3),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_64),
.C(n_30),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_64),
.C(n_30),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_23),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.C1(n_9),
.C2(n_7),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_289),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_290),
.C(n_285),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_7),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_291),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_7),
.A3(n_12),
.B1(n_11),
.B2(n_9),
.C1(n_13),
.C2(n_6),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_11),
.Y(n_291)
);

AO21x1_ASAP7_75t_SL g299 ( 
.A1(n_292),
.A2(n_293),
.B(n_296),
.Y(n_299)
);

AOI31xp67_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_272),
.A3(n_278),
.B(n_271),
.Y(n_293)
);

AOI31xp67_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_270),
.A3(n_12),
.B(n_13),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_1),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_6),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_4),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_299),
.B(n_4),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_5),
.C(n_304),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_5),
.Y(n_308)
);


endmodule