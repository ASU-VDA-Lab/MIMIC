module real_jpeg_25620_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_28),
.B1(n_51),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_28),
.B1(n_56),
.B2(n_57),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_54),
.B(n_163),
.C(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_55),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_57),
.B(n_77),
.C(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_1),
.B(n_22),
.C(n_35),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_1),
.B(n_75),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_1),
.B(n_11),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_1),
.B(n_38),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_4),
.A2(n_43),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_6),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_6),
.A2(n_33),
.B1(n_37),
.B2(n_105),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_105),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_40),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_132),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_130),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_106),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_106),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_85),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_64),
.B2(n_65),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_20),
.A2(n_29),
.B1(n_45),
.B2(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_20),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_20),
.A2(n_45),
.B1(n_189),
.B2(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_27),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_21),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_21),
.B(n_27),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_21),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_22),
.B(n_230),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_28),
.A2(n_53),
.B(n_57),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_28),
.A2(n_37),
.B(n_79),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_29),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_30),
.A2(n_68),
.B(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_31),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_31),
.B(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_31),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_32)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_33),
.A2(n_37),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_33),
.B(n_207),
.Y(n_206)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_38),
.B(n_194),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_39),
.A2(n_70),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_41),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_41),
.B(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_59),
.B(n_60),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_49),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_49),
.B(n_61),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_51),
.Y(n_164)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_55),
.B(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_57),
.B1(n_77),
.B2(n_79),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_73),
.B(n_84),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_67),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_72),
.B(n_204),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_80),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_75),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_83),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_81),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_76),
.B(n_123),
.Y(n_156)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_80),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_81),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.C(n_100),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_87),
.B(n_93),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_88),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_89),
.B(n_219),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_91),
.A2(n_116),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_91),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_100),
.B1(n_101),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_95),
.B(n_154),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_97),
.B(n_147),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_107),
.B(n_110),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_112),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_124),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_113),
.A2(n_114),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_120),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_118),
.B(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_122),
.A2(n_124),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_122),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_124),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_269),
.B(n_273),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_182),
.B(n_255),
.C(n_268),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_170),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_135),
.B(n_170),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_151),
.B2(n_169),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_149),
.B2(n_150),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_138),
.B(n_150),
.C(n_169),
.Y(n_256)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_141),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_161),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_153),
.B(n_160),
.C(n_161),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.C(n_177),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_172),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_254),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_198),
.B(n_253),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_185),
.B(n_195),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_191),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_191),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_189),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_248),
.B(n_252),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_239),
.B(n_247),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_221),
.B(n_238),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_202),
.B(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_220),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_214),
.C(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_237),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_236),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_265),
.B2(n_266),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_266),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);


endmodule