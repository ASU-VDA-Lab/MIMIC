module fake_jpeg_9152_n_71 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_48;
wire n_35;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_14),
.B1(n_18),
.B2(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_12),
.C(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_42),
.B1(n_44),
.B2(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_1),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_2),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B(n_39),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_54),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_43),
.B1(n_38),
.B2(n_13),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_6),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_59),
.B(n_61),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_56),
.C(n_16),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_11),
.C(n_17),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_19),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_23),
.C(n_25),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_26),
.A3(n_27),
.B1(n_28),
.B2(n_30),
.C(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_57),
.Y(n_71)
);


endmodule