module fake_jpeg_32182_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_1),
.C(n_2),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_40),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_6),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_7),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_8),
.B(n_9),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_19),
.B(n_23),
.C(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_10),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_59),
.C(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_16),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_16),
.B1(n_24),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_21),
.B1(n_10),
.B2(n_11),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_11),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_67),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_73),
.B1(n_56),
.B2(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_31),
.C(n_30),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_31),
.B1(n_39),
.B2(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_46),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_89),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_88),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_97),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_60),
.C(n_67),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_77),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_75),
.B1(n_70),
.B2(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_72),
.B(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_57),
.B1(n_68),
.B2(n_43),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_103),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_89),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_107),
.B(n_96),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_91),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_78),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_78),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_94),
.B(n_90),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_101),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_86),
.C(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_108),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_103),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_86),
.B(n_49),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_114),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_121),
.B(n_49),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);


endmodule