module fake_netlist_5_2026_n_112 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_112);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_112;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_0),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_34),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_36),
.B(n_48),
.C(n_25),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_25),
.B(n_24),
.C(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_43),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_45),
.B(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_44),
.B1(n_47),
.B2(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

AO32x2_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_24),
.A3(n_50),
.B1(n_27),
.B2(n_45),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_57),
.B(n_50),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_50),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_51),
.B(n_52),
.C(n_42),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_52),
.B(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_R g74 ( 
.A(n_64),
.B(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_71),
.Y(n_76)
);

AO21x2_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_66),
.B(n_69),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_66),
.B1(n_37),
.B2(n_45),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_81),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_79),
.B(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_89),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_88),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_68),
.B(n_71),
.Y(n_98)
);

OAI221xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_74),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_77),
.B(n_78),
.Y(n_100)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_45),
.B1(n_83),
.B2(n_7),
.C(n_8),
.Y(n_101)
);

OAI211xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_85),
.B(n_87),
.C(n_8),
.Y(n_102)
);

OAI211xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_101),
.B(n_102),
.C(n_100),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_99),
.A2(n_94),
.B(n_6),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_85),
.B(n_9),
.C(n_2),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

OAI322xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_106),
.A3(n_105),
.B1(n_2),
.B2(n_73),
.C1(n_16),
.C2(n_17),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_73),
.B1(n_14),
.B2(n_77),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_56),
.B(n_77),
.C(n_107),
.Y(n_112)
);


endmodule