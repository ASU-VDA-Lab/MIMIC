module fake_jpeg_26987_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_29),
.B1(n_30),
.B2(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_47),
.B1(n_15),
.B2(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_29),
.B1(n_30),
.B2(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_29),
.B1(n_30),
.B2(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_17),
.B1(n_16),
.B2(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_26),
.B1(n_31),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_15),
.B1(n_28),
.B2(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_62),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_80),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_77),
.B1(n_24),
.B2(n_32),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_49),
.B1(n_19),
.B2(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_31),
.B1(n_17),
.B2(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_110),
.B1(n_83),
.B2(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_49),
.B1(n_35),
.B2(n_32),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_103),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_39),
.A3(n_37),
.B1(n_32),
.B2(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_69),
.B1(n_72),
.B2(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_51),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_49),
.B1(n_32),
.B2(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_108),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_48),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_59),
.B(n_37),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_79),
.B(n_1),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_39),
.B1(n_37),
.B2(n_48),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_61),
.B1(n_74),
.B2(n_71),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_122),
.B1(n_123),
.B2(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_77),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_66),
.B1(n_81),
.B2(n_75),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_131),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_37),
.B1(n_57),
.B2(n_43),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_96),
.B1(n_98),
.B2(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_108),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_85),
.B(n_57),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_134),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_68),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_124),
.B(n_119),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_68),
.B1(n_24),
.B2(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_68),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_109),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_93),
.B1(n_90),
.B2(n_99),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_132),
.C(n_119),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_164),
.C(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_97),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_141),
.B(n_155),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_159),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_110),
.B(n_100),
.C(n_89),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_154),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_100),
.B(n_107),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_166),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_102),
.C(n_9),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_11),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_96),
.B(n_98),
.C(n_99),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_126),
.C(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_104),
.B1(n_12),
.B2(n_11),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_124),
.B1(n_117),
.B2(n_133),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_143),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_180),
.B1(n_192),
.B2(n_167),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_129),
.B1(n_122),
.B2(n_135),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_189),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_130),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_184),
.B(n_146),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_121),
.C(n_104),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_195),
.C(n_147),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_0),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_152),
.Y(n_201)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_12),
.C(n_10),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_159),
.B(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_201),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_202),
.B1(n_172),
.B2(n_142),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_139),
.B1(n_166),
.B2(n_153),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_209),
.C(n_184),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_178),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_163),
.B(n_148),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_210),
.B(n_174),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_146),
.C(n_148),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_163),
.B(n_148),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_161),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_215),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_196),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_217),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_161),
.B1(n_151),
.B2(n_142),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_179),
.B1(n_180),
.B2(n_176),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_223),
.B1(n_232),
.B2(n_233),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_234),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_198),
.C(n_210),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_225),
.C(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_194),
.B1(n_181),
.B2(n_169),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_208),
.C(n_203),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_200),
.B(n_201),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_171),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_228),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_178),
.C(n_189),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_186),
.B1(n_182),
.B2(n_191),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_195),
.B1(n_193),
.B2(n_172),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_243),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_215),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_202),
.C(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_235),
.B1(n_226),
.B2(n_224),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_2),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_8),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_216),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_10),
.C(n_9),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_230),
.B1(n_228),
.B2(n_234),
.C(n_227),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_263),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_2),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_255)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_3),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_243),
.B(n_239),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_5),
.B(n_6),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_268),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_237),
.C(n_241),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_275),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_237),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_273),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_274),
.B(n_255),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_260),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_6),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_272),
.A2(n_259),
.B1(n_261),
.B2(n_260),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_259),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_282),
.C(n_5),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_267),
.B(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_288),
.C(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_5),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_279),
.C(n_278),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_285),
.B(n_283),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_291),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_295),
.A2(n_7),
.B1(n_290),
.B2(n_262),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_7),
.Y(n_297)
);


endmodule