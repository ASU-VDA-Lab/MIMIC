module fake_jpeg_19689_n_316 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_46),
.B1(n_35),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_20),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_18),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_57),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_34),
.B1(n_29),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_60),
.B1(n_68),
.B2(n_73),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_34),
.B1(n_29),
.B2(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_74),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_35),
.B1(n_31),
.B2(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_21),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_43),
.B1(n_49),
.B2(n_32),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_79),
.B1(n_101),
.B2(n_105),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_23),
.B1(n_17),
.B2(n_26),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_85),
.Y(n_147)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_57),
.B1(n_72),
.B2(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_86),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_87),
.Y(n_150)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_26),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_4),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_20),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_55),
.A2(n_19),
.B1(n_30),
.B2(n_25),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_19),
.B1(n_27),
.B2(n_30),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_110),
.B(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_32),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_1),
.B(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_114),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_57),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_25),
.B1(n_27),
.B2(n_20),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_69),
.B1(n_55),
.B2(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_84),
.B1(n_91),
.B2(n_85),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_69),
.B1(n_72),
.B2(n_75),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_117),
.A2(n_131),
.B1(n_143),
.B2(n_141),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_27),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_1),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_127),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_4),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_129),
.B(n_110),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_10),
.C(n_6),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_112),
.C(n_76),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_96),
.B(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_144),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_15),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_6),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_14),
.B(n_11),
.C(n_12),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_9),
.Y(n_167)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_165),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_176),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_93),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_87),
.B(n_81),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_138),
.B(n_129),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_77),
.B(n_107),
.C(n_111),
.D(n_112),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_163),
.B(n_128),
.C(n_160),
.D(n_159),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_76),
.C(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_102),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_102),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_90),
.C(n_82),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_123),
.C(n_150),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_124),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_90),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

OR2x4_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_82),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_126),
.B(n_142),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_80),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_101),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_134),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_139),
.C(n_127),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_166),
.B(n_145),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_204),
.B(n_206),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_148),
.B1(n_137),
.B2(n_136),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_212),
.B1(n_210),
.B2(n_199),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_188),
.B(n_196),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_154),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_120),
.Y(n_196)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_201),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_175),
.B(n_142),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_134),
.B1(n_146),
.B2(n_116),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_211),
.B1(n_178),
.B2(n_158),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_210),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_125),
.B1(n_145),
.B2(n_83),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_154),
.C(n_173),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_223),
.C(n_227),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_224),
.B1(n_206),
.B2(n_190),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_170),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_221),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_182),
.C(n_153),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_181),
.B1(n_175),
.B2(n_153),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_191),
.C(n_207),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_174),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_185),
.A2(n_160),
.B1(n_174),
.B2(n_152),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_160),
.B(n_175),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_234),
.B(n_193),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_209),
.B1(n_190),
.B2(n_193),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_184),
.B(n_158),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_211),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_207),
.C(n_203),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_233),
.C(n_223),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_228),
.B1(n_236),
.B2(n_234),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_246),
.A2(n_255),
.B1(n_235),
.B2(n_232),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_247),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_183),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_231),
.B(n_195),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_195),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_229),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_267),
.B(n_238),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_259),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_214),
.C(n_233),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_263),
.C(n_270),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_240),
.C(n_244),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_273),
.B1(n_248),
.B2(n_246),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_198),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_R g277 ( 
.A(n_269),
.B(n_268),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_194),
.C(n_192),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_166),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_272),
.C(n_250),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_137),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_217),
.B1(n_226),
.B2(n_192),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_269),
.B(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_282),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_248),
.B1(n_254),
.B2(n_247),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_238),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_242),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_252),
.B1(n_226),
.B2(n_125),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_130),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_263),
.C(n_258),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_265),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_272),
.B(n_259),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_280),
.B(n_275),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_283),
.B1(n_278),
.B2(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_197),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_300),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_302),
.B(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_284),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_276),
.B1(n_118),
.B2(n_14),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_304),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_299),
.B(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_294),
.B(n_289),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.C(n_12),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_308),
.B1(n_276),
.B2(n_13),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_312),
.Y(n_314)
);

XOR2x2_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_13),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_13),
.Y(n_316)
);


endmodule