module real_aes_8373_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_397;
wire n_275;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_0), .A2(n_71), .B1(n_491), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_1), .A2(n_168), .B1(n_696), .B2(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_2), .A2(n_254), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_3), .A2(n_197), .B1(n_356), .B2(n_359), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_4), .A2(n_228), .B1(n_323), .B2(n_330), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_5), .A2(n_99), .B1(n_367), .B2(n_595), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g835 ( .A1(n_6), .A2(n_31), .B1(n_115), .B2(n_410), .C1(n_414), .C2(n_695), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_7), .A2(n_33), .B1(n_367), .B2(n_643), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_8), .A2(n_118), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_9), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_10), .A2(n_124), .B1(n_378), .B2(n_379), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_11), .A2(n_207), .B1(n_523), .B2(n_526), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_12), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_13), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_14), .A2(n_35), .B1(n_361), .B2(n_560), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_15), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_16), .A2(n_221), .B1(n_340), .B2(n_491), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_17), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_18), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_19), .B(n_418), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_20), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_21), .A2(n_125), .B1(n_461), .B2(n_549), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_22), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_23), .A2(n_100), .B1(n_811), .B2(n_813), .C(n_814), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_24), .A2(n_44), .B1(n_711), .B2(n_830), .C(n_831), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_25), .A2(n_204), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_26), .A2(n_264), .B1(n_553), .B2(n_591), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_27), .Y(n_609) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_28), .A2(n_88), .B1(n_292), .B2(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g805 ( .A(n_28), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_29), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_30), .A2(n_236), .B1(n_448), .B2(n_560), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_32), .A2(n_73), .B1(n_530), .B2(n_821), .C(n_824), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_34), .A2(n_256), .B1(n_367), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_36), .A2(n_150), .B1(n_437), .B2(n_521), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_37), .A2(n_185), .B1(n_597), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_38), .A2(n_47), .B1(n_365), .B2(n_525), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_39), .A2(n_130), .B1(n_443), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_40), .A2(n_231), .B1(n_521), .B2(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_41), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_42), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_43), .A2(n_186), .B1(n_387), .B2(n_683), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_45), .A2(n_161), .B1(n_362), .B2(n_601), .Y(n_600) );
AO22x2_ASAP7_75t_L g295 ( .A1(n_46), .A2(n_91), .B1(n_292), .B2(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g806 ( .A(n_46), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_48), .A2(n_98), .B1(n_448), .B2(n_634), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_49), .A2(n_242), .B1(n_633), .B2(n_634), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_50), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_51), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_52), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_53), .B(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_54), .A2(n_203), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_55), .A2(n_237), .B1(n_356), .B2(n_643), .Y(n_642) );
AOI222xp33_ASAP7_75t_L g767 ( .A1(n_56), .A2(n_147), .B1(n_159), .B2(n_289), .C1(n_304), .C2(n_768), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_57), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_58), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_59), .A2(n_110), .B1(n_357), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_60), .A2(n_149), .B1(n_414), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_61), .A2(n_139), .B1(n_366), .B2(n_643), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_62), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_63), .A2(n_225), .B1(n_310), .B2(n_696), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_64), .A2(n_230), .B1(n_648), .B2(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_65), .A2(n_172), .B1(n_511), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_66), .A2(n_86), .B1(n_310), .B2(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_67), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_68), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_69), .A2(n_122), .B1(n_364), .B2(n_366), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_70), .A2(n_129), .B1(n_415), .B2(n_461), .Y(n_460) );
XNOR2x2_ASAP7_75t_L g747 ( .A(n_72), .B(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_74), .Y(n_845) );
OA22x2_ASAP7_75t_L g846 ( .A1(n_74), .A2(n_845), .B1(n_847), .B2(n_864), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_75), .B(n_665), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_76), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_77), .A2(n_95), .B1(n_648), .B2(n_649), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_78), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_79), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g694 ( .A1(n_80), .A2(n_156), .B1(n_166), .B2(n_410), .C1(n_695), .C2(n_696), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g303 ( .A1(n_81), .A2(n_219), .B1(n_304), .B2(n_310), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_82), .A2(n_83), .B1(n_485), .B2(n_529), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g322 ( .A1(n_84), .A2(n_135), .B1(n_323), .B2(n_330), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_85), .A2(n_148), .B1(n_316), .B2(n_455), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g742 ( .A1(n_87), .A2(n_90), .B1(n_121), .B2(n_289), .C1(n_455), .C2(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_89), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_92), .Y(n_612) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_93), .A2(n_253), .B1(n_478), .B2(n_511), .Y(n_782) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_94), .A2(n_215), .B1(n_736), .B2(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g277 ( .A(n_96), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_97), .A2(n_249), .B1(n_387), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_101), .A2(n_265), .B1(n_601), .B2(n_724), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_102), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_103), .A2(n_374), .B1(n_428), .B2(n_429), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_103), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_104), .Y(n_790) );
INVx1_ASAP7_75t_L g274 ( .A(n_105), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_106), .A2(n_173), .B1(n_379), .B2(n_485), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_107), .A2(n_238), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_108), .A2(n_127), .B1(n_311), .B2(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_109), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_111), .A2(n_232), .B1(n_437), .B2(n_439), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_112), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_113), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_114), .B(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_116), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g857 ( .A1(n_117), .A2(n_205), .B1(n_446), .B2(n_858), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_119), .A2(n_123), .B1(n_682), .B2(n_683), .Y(n_681) );
OA22x2_ASAP7_75t_L g466 ( .A1(n_120), .A2(n_467), .B1(n_468), .B2(n_493), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_120), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_126), .A2(n_137), .B1(n_589), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_128), .A2(n_157), .B1(n_643), .B2(n_717), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_131), .A2(n_250), .B1(n_347), .B2(n_383), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_132), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_133), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_134), .B(n_323), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_136), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_138), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g278 ( .A(n_140), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_141), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_142), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_143), .A2(n_171), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_144), .A2(n_268), .B1(n_304), .B2(n_418), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_145), .A2(n_152), .B1(n_437), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_146), .A2(n_151), .B1(n_719), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_153), .A2(n_266), .B1(n_346), .B2(n_351), .Y(n_859) );
AND2x6_ASAP7_75t_L g273 ( .A(n_154), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_154), .Y(n_799) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_155), .A2(n_218), .B1(n_292), .B2(n_296), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_158), .A2(n_184), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g335 ( .A1(n_160), .A2(n_224), .B1(n_336), .B2(n_340), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_162), .B(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_163), .A2(n_247), .B1(n_442), .B2(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_164), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g345 ( .A1(n_165), .A2(n_259), .B1(n_346), .B2(n_351), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_167), .A2(n_201), .B1(n_446), .B2(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g534 ( .A(n_169), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_170), .A2(n_222), .B1(n_315), .B2(n_319), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_174), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_175), .A2(n_183), .B1(n_304), .B2(n_316), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_176), .B(n_614), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_177), .A2(n_198), .B1(n_365), .B2(n_382), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_178), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_179), .A2(n_269), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_180), .A2(n_211), .B1(n_381), .B2(n_383), .Y(n_380) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_181), .A2(n_240), .B1(n_292), .B2(n_293), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_182), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_187), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_188), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_189), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_190), .A2(n_202), .B1(n_652), .B2(n_682), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_191), .Y(n_661) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_192), .A2(n_234), .B1(n_520), .B2(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_193), .Y(n_818) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_194), .A2(n_271), .B(n_279), .C(n_807), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_195), .A2(n_217), .B1(n_461), .B2(n_549), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_196), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_199), .A2(n_639), .B1(n_670), .B2(n_671), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_199), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_200), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_206), .Y(n_545) );
INVx1_ASAP7_75t_L g761 ( .A(n_208), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_209), .A2(n_246), .B1(n_520), .B2(n_521), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_210), .B(n_689), .Y(n_709) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_212), .A2(n_251), .B1(n_310), .B2(n_549), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_213), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_214), .B(n_781), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_216), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_218), .B(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_220), .Y(n_667) );
OA22x2_ASAP7_75t_L g283 ( .A1(n_223), .A2(n_284), .B1(n_285), .B2(n_369), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_223), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_226), .Y(n_412) );
INVx1_ASAP7_75t_L g433 ( .A(n_227), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_229), .B(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_233), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_235), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_239), .Y(n_850) );
INVx1_ASAP7_75t_L g802 ( .A(n_240), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_241), .A2(n_257), .B1(n_446), .B2(n_485), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_243), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_244), .A2(n_248), .B1(n_340), .B2(n_448), .Y(n_492) );
XNOR2x2_ASAP7_75t_L g727 ( .A(n_245), .B(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_252), .Y(n_562) );
INVx1_ASAP7_75t_L g292 ( .A(n_255), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_255), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_258), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_260), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_261), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_262), .Y(n_554) );
OA22x2_ASAP7_75t_L g537 ( .A1(n_263), .A2(n_538), .B1(n_539), .B2(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_263), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_267), .A2(n_809), .B1(n_836), .B2(n_837), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_267), .Y(n_836) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_274), .Y(n_798) );
OA21x2_ASAP7_75t_L g843 ( .A1(n_275), .A2(n_797), .B(n_844), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_575), .B1(n_792), .B2(n_793), .C(n_794), .Y(n_279) );
INVx1_ASAP7_75t_L g792 ( .A(n_280), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_430), .B1(n_573), .B2(n_574), .Y(n_280) );
INVx1_ASAP7_75t_L g573 ( .A(n_281), .Y(n_573) );
OAI22xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_283), .B1(n_370), .B2(n_371), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g369 ( .A(n_285), .Y(n_369) );
NAND3x1_ASAP7_75t_L g285 ( .A(n_286), .B(n_334), .C(n_354), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_313), .Y(n_286) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_302), .B(n_303), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_288), .A2(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx4_ASAP7_75t_L g411 ( .A(n_289), .Y(n_411) );
BUFx3_ASAP7_75t_L g458 ( .A(n_289), .Y(n_458) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_289), .Y(n_486) );
INVx2_ASAP7_75t_L g660 ( .A(n_289), .Y(n_660) );
AND2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_297), .Y(n_289) );
AND2x4_ASAP7_75t_L g319 ( .A(n_290), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g406 ( .A(n_290), .Y(n_406) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
AND2x2_ASAP7_75t_L g309 ( .A(n_291), .B(n_299), .Y(n_309) );
INVx2_ASAP7_75t_L g329 ( .A(n_291), .Y(n_329) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g296 ( .A(n_294), .Y(n_296) );
INVx2_ASAP7_75t_L g308 ( .A(n_295), .Y(n_308) );
INVx1_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
OR2x2_ASAP7_75t_L g328 ( .A(n_295), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_295), .B(n_329), .Y(n_333) );
AND2x6_ASAP7_75t_L g339 ( .A(n_297), .B(n_327), .Y(n_339) );
AND2x2_ASAP7_75t_L g358 ( .A(n_297), .B(n_344), .Y(n_358) );
AND2x4_ASAP7_75t_L g365 ( .A(n_297), .B(n_333), .Y(n_365) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
AND2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_301), .Y(n_326) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_299), .B(n_301), .Y(n_343) );
AND2x2_ASAP7_75t_L g350 ( .A(n_299), .B(n_321), .Y(n_350) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g307 ( .A(n_301), .Y(n_307) );
INVx1_ASAP7_75t_L g321 ( .A(n_301), .Y(n_321) );
BUFx4f_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_305), .Y(n_415) );
BUFx2_ASAP7_75t_L g488 ( .A(n_305), .Y(n_488) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_305), .Y(n_511) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_305), .Y(n_553) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g312 ( .A(n_307), .Y(n_312) );
AND2x2_ASAP7_75t_L g344 ( .A(n_308), .B(n_329), .Y(n_344) );
INVx1_ASAP7_75t_L g401 ( .A(n_308), .Y(n_401) );
AND2x4_ASAP7_75t_L g311 ( .A(n_309), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g316 ( .A(n_309), .B(n_317), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g400 ( .A(n_309), .B(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g418 ( .A(n_310), .Y(n_418) );
BUFx3_ASAP7_75t_L g665 ( .A(n_310), .Y(n_665) );
INVx2_ASAP7_75t_L g744 ( .A(n_310), .Y(n_744) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx12f_ASAP7_75t_L g461 ( .A(n_311), .Y(n_461) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_311), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_322), .Y(n_313) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g478 ( .A(n_316), .Y(n_478) );
BUFx3_ASAP7_75t_L g591 ( .A(n_316), .Y(n_591) );
INVx1_ASAP7_75t_L g737 ( .A(n_316), .Y(n_737) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x6_ASAP7_75t_L g353 ( .A(n_318), .B(n_343), .Y(n_353) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_319), .Y(n_455) );
BUFx2_ASAP7_75t_SL g549 ( .A(n_319), .Y(n_549) );
BUFx2_ASAP7_75t_SL g696 ( .A(n_319), .Y(n_696) );
BUFx3_ASAP7_75t_L g854 ( .A(n_319), .Y(n_854) );
INVx1_ASAP7_75t_L g407 ( .A(n_320), .Y(n_407) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g830 ( .A(n_323), .Y(n_830) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g689 ( .A(n_324), .Y(n_689) );
INVx2_ASAP7_75t_L g734 ( .A(n_324), .Y(n_734) );
INVx5_ASAP7_75t_L g764 ( .A(n_324), .Y(n_764) );
INVx4_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x6_ASAP7_75t_L g332 ( .A(n_326), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g362 ( .A(n_326), .B(n_344), .Y(n_362) );
INVx1_ASAP7_75t_L g423 ( .A(n_326), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_326), .B(n_333), .Y(n_427) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g422 ( .A(n_328), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g589 ( .A(n_332), .Y(n_589) );
BUFx4f_ASAP7_75t_L g711 ( .A(n_332), .Y(n_711) );
BUFx2_ASAP7_75t_L g779 ( .A(n_332), .Y(n_779) );
AND2x2_ASAP7_75t_L g349 ( .A(n_333), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_333), .B(n_350), .Y(n_817) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_345), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
INVx5_ASAP7_75t_SL g595 ( .A(n_338), .Y(n_595) );
INVx4_ASAP7_75t_L g716 ( .A(n_338), .Y(n_716) );
INVx2_ASAP7_75t_L g751 ( .A(n_338), .Y(n_751) );
INVx2_ASAP7_75t_SL g823 ( .A(n_338), .Y(n_823) );
INVx11_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx11_ASAP7_75t_L g440 ( .A(n_339), .Y(n_440) );
INVxp67_ASAP7_75t_L g396 ( .A(n_340), .Y(n_396) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g449 ( .A(n_341), .Y(n_449) );
BUFx2_ASAP7_75t_SL g521 ( .A(n_341), .Y(n_521) );
BUFx3_ASAP7_75t_L g597 ( .A(n_341), .Y(n_597) );
BUFx3_ASAP7_75t_L g719 ( .A(n_341), .Y(n_719) );
BUFx2_ASAP7_75t_SL g789 ( .A(n_341), .Y(n_789) );
BUFx3_ASAP7_75t_L g813 ( .A(n_341), .Y(n_813) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
AND2x2_ASAP7_75t_L g443 ( .A(n_342), .B(n_401), .Y(n_443) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g368 ( .A(n_344), .B(n_350), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_344), .B(n_350), .Y(n_392) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
INVx5_ASAP7_75t_L g442 ( .A(n_348), .Y(n_442) );
INVx4_ASAP7_75t_L g525 ( .A(n_348), .Y(n_525) );
BUFx3_ASAP7_75t_L g684 ( .A(n_348), .Y(n_684) );
INVx3_ASAP7_75t_L g722 ( .A(n_348), .Y(n_722) );
INVx8_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
BUFx2_ASAP7_75t_L g560 ( .A(n_352), .Y(n_560) );
BUFx2_ASAP7_75t_L g634 ( .A(n_352), .Y(n_634) );
BUFx4f_ASAP7_75t_SL g653 ( .A(n_352), .Y(n_653) );
INVx6_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_353), .A2(n_405), .B1(n_480), .B2(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g526 ( .A(n_353), .Y(n_526) );
INVx1_ASAP7_75t_SL g601 ( .A(n_353), .Y(n_601) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_363), .Y(n_354) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g378 ( .A(n_357), .Y(n_378) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_357), .Y(n_757) );
INVx3_ASAP7_75t_L g812 ( .A(n_357), .Y(n_812) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g438 ( .A(n_358), .Y(n_438) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_358), .Y(n_520) );
BUFx2_ASAP7_75t_SL g741 ( .A(n_358), .Y(n_741) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_360), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g645 ( .A(n_361), .Y(n_645) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g448 ( .A(n_362), .Y(n_448) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_362), .Y(n_532) );
BUFx3_ASAP7_75t_L g633 ( .A(n_362), .Y(n_633) );
INVx2_ASAP7_75t_L g725 ( .A(n_362), .Y(n_725) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx6_ASAP7_75t_L g388 ( .A(n_365), .Y(n_388) );
BUFx3_ASAP7_75t_L g446 ( .A(n_365), .Y(n_446) );
BUFx3_ASAP7_75t_L g827 ( .A(n_365), .Y(n_827) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g485 ( .A(n_368), .Y(n_485) );
BUFx3_ASAP7_75t_L g717 ( .A(n_368), .Y(n_717) );
BUFx3_ASAP7_75t_L g758 ( .A(n_368), .Y(n_758) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_375), .B(n_397), .Y(n_374) );
NOR3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_384), .C(n_393), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
INVx2_ASAP7_75t_L g567 ( .A(n_379), .Y(n_567) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g819 ( .A(n_383), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_389), .B2(n_390), .Y(n_384) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g648 ( .A(n_388), .Y(n_648) );
INVx2_ASAP7_75t_L g682 ( .A(n_388), .Y(n_682) );
INVx3_ASAP7_75t_L g752 ( .A(n_388), .Y(n_752) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g570 ( .A(n_391), .Y(n_570) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR3xp33_ASAP7_75t_SL g397 ( .A(n_398), .B(n_408), .C(n_419), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_402), .B2(n_403), .Y(n_398) );
INVx4_ASAP7_75t_L g515 ( .A(n_400), .Y(n_515) );
BUFx3_ASAP7_75t_L g555 ( .A(n_400), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_403), .A2(n_513), .B1(n_514), .B2(n_516), .Y(n_512) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g658 ( .A(n_404), .Y(n_658) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_405), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B1(n_413), .B2(n_416), .C(n_417), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx4_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g508 ( .A(n_411), .Y(n_508) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g623 ( .A(n_415), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_424), .B2(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g619 ( .A(n_421), .Y(n_619) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_422), .A2(n_451), .B1(n_452), .B2(n_453), .C(n_454), .Y(n_450) );
BUFx3_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
INVx2_ASAP7_75t_L g502 ( .A(n_422), .Y(n_502) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g474 ( .A(n_426), .Y(n_474) );
INVx1_ASAP7_75t_L g762 ( .A(n_426), .Y(n_762) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g452 ( .A(n_427), .Y(n_452) );
INVx1_ASAP7_75t_L g574 ( .A(n_430), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_462), .B2(n_572), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
XNOR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
NOR4xp75_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .C(n_450), .D(n_456), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_436), .B(n_441), .Y(n_435) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g491 ( .A(n_438), .Y(n_491) );
INVx4_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI21xp33_ASAP7_75t_SL g475 ( .A1(n_440), .A2(n_476), .B(n_477), .Y(n_475) );
INVx2_ASAP7_75t_SL g529 ( .A(n_440), .Y(n_529) );
INVx4_ASAP7_75t_L g643 ( .A(n_440), .Y(n_643) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_442), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx2_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
BUFx3_ASAP7_75t_L g669 ( .A(n_452), .Y(n_669) );
INVx1_ASAP7_75t_SL g615 ( .A(n_455), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_459), .B(n_460), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_457), .A2(n_547), .B(n_548), .Y(n_546) );
OAI21xp5_ASAP7_75t_SL g849 ( .A1(n_457), .A2(n_850), .B(n_851), .Y(n_849) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx4f_ASAP7_75t_SL g695 ( .A(n_461), .Y(n_695) );
INVx1_ASAP7_75t_L g572 ( .A(n_462), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_494), .B2(n_571), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g493 ( .A(n_468), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_482), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_475), .C(n_479), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_470) );
OA211x2_ASAP7_75t_L g686 ( .A1(n_474), .A2(n_687), .B(n_688), .C(n_690), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g650 ( .A(n_485), .Y(n_650) );
INVx2_ASAP7_75t_L g608 ( .A(n_486), .Y(n_608) );
INVx1_ASAP7_75t_L g662 ( .A(n_488), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g571 ( .A(n_494), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_535), .B2(n_536), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_534), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_517), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_506), .C(n_512), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_503), .B2(n_504), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_501), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_666) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g542 ( .A1(n_504), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_504), .A2(n_617), .B1(n_618), .B2(n_620), .Y(n_616) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
BUFx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_514), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
INVx3_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g833 ( .A(n_515), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_L g563 ( .A(n_520), .Y(n_563) );
INVx1_ASAP7_75t_SL g565 ( .A(n_521), .Y(n_565) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_525), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
INVx4_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g754 ( .A(n_531), .Y(n_754) );
INVx4_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_556), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .C(n_550), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_554), .B2(n_555), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_555), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .C(n_566), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_570), .A2(n_825), .B1(n_826), .B2(n_828), .Y(n_824) );
INVx1_ASAP7_75t_L g793 ( .A(n_575), .Y(n_793) );
XOR2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_746), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_578), .B1(n_674), .B2(n_675), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_637), .B1(n_672), .B2(n_673), .Y(n_578) );
INVx2_ASAP7_75t_SL g672 ( .A(n_579), .Y(n_672) );
AO22x2_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_603), .B1(n_604), .B2(n_636), .Y(n_579) );
INVx3_ASAP7_75t_L g636 ( .A(n_580), .Y(n_636) );
XOR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_602), .Y(n_580) );
NAND2x1_ASAP7_75t_SL g581 ( .A(n_582), .B(n_592), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .C(n_590), .Y(n_586) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_598), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
BUFx2_ASAP7_75t_L g863 ( .A(n_597), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_635), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_625), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_616), .C(n_621), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_610), .B2(n_612), .C(n_613), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_608), .A2(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx4f_ASAP7_75t_L g768 ( .A(n_611), .Y(n_768) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
BUFx2_ASAP7_75t_L g858 ( .A(n_633), .Y(n_858) );
INVx1_ASAP7_75t_L g673 ( .A(n_637), .Y(n_673) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g671 ( .A(n_639), .Y(n_671) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_640), .B(n_654), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_646), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_659), .C(n_666), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_658), .A2(n_832), .B1(n_833), .B2(n_834), .Y(n_831) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .C(n_664), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g774 ( .A1(n_660), .A2(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_698), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
XNOR2x2_ASAP7_75t_L g770 ( .A(n_678), .B(n_771), .Y(n_770) );
XOR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_697), .Y(n_678) );
NAND4xp75_ASAP7_75t_L g679 ( .A(n_680), .B(n_686), .C(n_691), .D(n_694), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_685), .Y(n_680) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_727), .B2(n_745), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
XOR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_726), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_704), .B(n_713), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .C(n_712), .Y(n_708) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_720), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g745 ( .A(n_727), .Y(n_745) );
NAND4xp75_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .C(n_738), .D(n_742), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
AND2x2_ASAP7_75t_SL g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g766 ( .A(n_737), .Y(n_766) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_769), .B1(n_770), .B2(n_791), .Y(n_746) );
INVx1_ASAP7_75t_L g791 ( .A(n_747), .Y(n_791) );
NAND4xp75_ASAP7_75t_L g748 ( .A(n_749), .B(n_755), .C(n_760), .D(n_767), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
OA211x2_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B(n_763), .C(n_765), .Y(n_760) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_764), .Y(n_781) );
INVx2_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
XOR2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_790), .Y(n_771) );
NAND3x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_783), .C(n_786), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .C(n_782), .Y(n_777) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .Y(n_795) );
OR2x2_ASAP7_75t_SL g866 ( .A(n_796), .B(n_801), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_798), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_798), .B(n_842), .Y(n_844) );
CKINVDCx16_ASAP7_75t_R g842 ( .A(n_799), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
OAI322xp33_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_838), .A3(n_839), .B1(n_843), .B2(n_845), .C1(n_846), .C2(n_865), .Y(n_807) );
INVx1_ASAP7_75t_L g837 ( .A(n_809), .Y(n_837) );
AND4x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_820), .C(n_829), .D(n_835), .Y(n_809) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_818), .B2(n_819), .Y(n_814) );
BUFx2_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_SL g864 ( .A(n_847), .Y(n_864) );
NAND3x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_856), .C(n_860), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_852), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
AND2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_859), .Y(n_856) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
endmodule