module fake_jpeg_25187_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx16f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_SL g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.C(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_9),
.B(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_9),
.B(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_12),
.B(n_6),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_16),
.B1(n_6),
.B2(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_6),
.B1(n_11),
.B2(n_8),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_13),
.C(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_7),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_11),
.B1(n_8),
.B2(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_3),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_26),
.C(n_13),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_7),
.Y(n_35)
);

OAI221xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_7),
.B1(n_1),
.B2(n_5),
.C(n_4),
.Y(n_36)
);


endmodule