module fake_jpeg_22913_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_13),
.B(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_37),
.Y(n_42)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_17),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_SL g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_54),
.B1(n_41),
.B2(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_59),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_76),
.Y(n_96)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_38),
.B1(n_41),
.B2(n_37),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_48),
.B1(n_53),
.B2(n_57),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_73),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_29),
.B1(n_30),
.B2(n_19),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_29),
.B1(n_28),
.B2(n_15),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_79),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_15),
.B(n_28),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_47),
.C(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_47),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_86),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_25),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_50),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_65),
.C(n_77),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_48),
.B1(n_39),
.B2(n_41),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_73),
.B1(n_70),
.B2(n_71),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_19),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_46),
.B1(n_20),
.B2(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_46),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_102),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_21),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_119),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_99),
.C(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_114),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_65),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_26),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_93),
.B1(n_80),
.B2(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_134),
.C(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_85),
.B(n_83),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_131),
.B(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_70),
.B1(n_23),
.B2(n_18),
.Y(n_154)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_84),
.C(n_97),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_25),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_87),
.B(n_30),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_92),
.C(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_109),
.B1(n_116),
.B2(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_150),
.B1(n_124),
.B2(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_134),
.C(n_123),
.Y(n_159)
);

OAI322xp33_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_112),
.A3(n_101),
.B1(n_113),
.B2(n_102),
.C1(n_107),
.C2(n_24),
.Y(n_147)
);

OAI322xp33_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_135),
.A3(n_128),
.B1(n_122),
.B2(n_10),
.C1(n_12),
.C2(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_151),
.B1(n_123),
.B2(n_131),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_2),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_82),
.B1(n_24),
.B2(n_23),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_71),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_141),
.B(n_145),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_158),
.B1(n_150),
.B2(n_143),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_163),
.C(n_164),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_156),
.CI(n_163),
.CON(n_172),
.SN(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_23),
.C(n_71),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_145),
.C(n_140),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_166),
.B(n_161),
.C(n_5),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_172),
.A2(n_177),
.B(n_178),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_142),
.C(n_139),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_12),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_2),
.C(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_186),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_173),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_3),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_173),
.C(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_179),
.C(n_8),
.Y(n_197)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_9),
.B(n_6),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_194),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_193),
.B(n_190),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_187),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_201),
.B(n_8),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_195),
.B(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.C(n_8),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_204),
.B(n_9),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_9),
.Y(n_206)
);


endmodule