module real_jpeg_16893_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_520),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_0),
.B(n_521),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_1),
.A2(n_325),
.B1(n_328),
.B2(n_331),
.Y(n_324)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_1),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_1),
.A2(n_331),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_1),
.A2(n_217),
.B1(n_331),
.B2(n_501),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_4),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_4),
.A2(n_86),
.B1(n_177),
.B2(n_182),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_4),
.A2(n_86),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_4),
.A2(n_86),
.B1(n_395),
.B2(n_438),
.Y(n_437)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_6),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_6),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_7),
.A2(n_105),
.B1(n_264),
.B2(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_7),
.A2(n_105),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_7),
.A2(n_105),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_8),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_8),
.Y(n_358)
);

BUFx8_ASAP7_75t_L g483 ( 
.A(n_8),
.Y(n_483)
);

BUFx5_ASAP7_75t_L g515 ( 
.A(n_8),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_9),
.A2(n_72),
.B1(n_73),
.B2(n_78),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_72),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_9),
.A2(n_72),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_9),
.A2(n_72),
.B1(n_338),
.B2(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_10),
.Y(n_279)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_10),
.Y(n_351)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_11),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_11),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_11),
.B(n_70),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_11),
.A2(n_43),
.B1(n_203),
.B2(n_208),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_224),
.A3(n_226),
.B1(n_227),
.B2(n_231),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_11),
.B(n_276),
.Y(n_275)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_11),
.A2(n_333),
.A3(n_337),
.B1(n_341),
.B2(n_345),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_11),
.A2(n_43),
.B1(n_362),
.B2(n_364),
.Y(n_361)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_12),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_13),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_14),
.A2(n_291),
.B1(n_297),
.B2(n_301),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_14),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_14),
.A2(n_301),
.B1(n_413),
.B2(n_415),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_14),
.A2(n_301),
.B1(n_473),
.B2(n_477),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_15),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_16),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_16),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_16),
.A2(n_250),
.B1(n_380),
.B2(n_382),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_16),
.A2(n_250),
.B1(n_442),
.B2(n_446),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_16),
.A2(n_250),
.B1(n_513),
.B2(n_514),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_17),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_490),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_456),
.B(n_488),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_384),
.B(n_453),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_310),
.B(n_383),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_255),
.B(n_309),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_169),
.B(n_254),
.Y(n_26)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_127),
.B(n_168),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_81),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_29),
.B(n_81),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_52),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_30),
.A2(n_52),
.B1(n_53),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_30),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.A3(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_33),
.Y(n_416)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_36),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_43),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_43),
.A2(n_91),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_43),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_43),
.B(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_49),
.A2(n_114),
.B1(n_115),
.B2(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_51),
.Y(n_330)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_111),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_70),
.B1(n_71),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_57),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_57),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_57),
.B(n_379),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_60),
.Y(n_183)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_66),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_66),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_66),
.A2(n_174),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_67),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_67),
.Y(n_253)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_67),
.Y(n_327)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_70),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_70),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_77),
.Y(n_230)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_80),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_107),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_82),
.B(n_108),
.C(n_119),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_91),
.B(n_96),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_131),
.B1(n_147),
.B2(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_91),
.B(n_246),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_91),
.A2(n_103),
.B(n_463),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_97),
.B(n_302),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_100),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_101),
.Y(n_245)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_103),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_119),
.Y(n_107)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_112),
.Y(n_428)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_114),
.A2(n_115),
.B1(n_216),
.B2(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_114),
.A2(n_115),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_120),
.B(n_441),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_120),
.A2(n_399),
.B1(n_499),
.B2(n_500),
.Y(n_498)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_125),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_142),
.B(n_167),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_140),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_140),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_135),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_135),
.A2(n_290),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_135),
.A2(n_242),
.B(n_324),
.Y(n_409)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_159),
.B(n_166),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_146),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_165),
.Y(n_166)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_162),
.A2(n_290),
.B(n_302),
.Y(n_289)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_170),
.B(n_171),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_222),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_184),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_173),
.B(n_184),
.C(n_222),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_174),
.A2(n_263),
.B(n_378),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_174),
.A2(n_378),
.B(n_426),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_183),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_202),
.B1(n_212),
.B2(n_221),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_185),
.A2(n_212),
.B1(n_221),
.B2(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_185),
.A2(n_221),
.B1(n_304),
.B2(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_185),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_185),
.A2(n_402),
.B(n_440),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_185),
.A2(n_221),
.B1(n_471),
.B2(n_472),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B1(n_195),
.B2(n_198),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_191),
.Y(n_374)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_193),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_193),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_205),
.Y(n_376)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_206),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_207),
.Y(n_344)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_208),
.Y(n_502)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_211),
.Y(n_477)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_221),
.B(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_240),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_240),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_235),
.Y(n_403)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_236),
.Y(n_445)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_236),
.Y(n_476)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_256),
.B(n_257),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_271),
.B1(n_272),
.B2(n_308),
.Y(n_257)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_271),
.C(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_262),
.B(n_504),
.Y(n_503)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_303),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_288),
.B2(n_289),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_303),
.C(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OR2x6_ASAP7_75t_L g354 ( 
.A(n_276),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_276),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_276),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_276),
.B(n_512),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B1(n_282),
.B2(n_285),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx2_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_313),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_352),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_316),
.B(n_318),
.C(n_352),
.Y(n_450)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_332),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_320),
.B(n_332),
.Y(n_406)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_351),
.A2(n_356),
.B1(n_357),
.B2(n_359),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_371),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_372),
.C(n_377),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_361),
.B1(n_367),
.B2(n_370),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_354),
.Y(n_392)
);

OAI22x1_ASAP7_75t_SL g436 ( 
.A1(n_354),
.A2(n_370),
.B1(n_394),
.B2(n_437),
.Y(n_436)
);

OAI21x1_ASAP7_75t_SL g478 ( 
.A1(n_354),
.A2(n_437),
.B(n_479),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_354),
.A2(n_510),
.B(n_511),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_360),
.Y(n_366)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_380),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_449),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_418),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_387),
.B(n_418),
.C(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_407),
.C(n_408),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_452),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_406),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_398),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_406),
.C(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_400),
.B(n_401),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_408),
.Y(n_452)
);

XOR2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_410),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_432),
.C(n_448),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_432),
.B1(n_433),
.B2(n_448),
.Y(n_421)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_424),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_436),
.C(n_439),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_439),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_459),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_468),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_468),
.C(n_485),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_461)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_462),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_SL g507 ( 
.A(n_462),
.B(n_466),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_462),
.A2(n_467),
.B1(n_509),
.B2(n_516),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2x1_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_484),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_478),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_472),
.Y(n_499)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_484),
.C(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_480),
.Y(n_510)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_519),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_493),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_506),
.B1(n_517),
.B2(n_518),
.Y(n_496)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

OAI21xp33_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_503),
.B(n_505),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_503),
.Y(n_505)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_509),
.Y(n_516)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx8_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);


endmodule