module fake_jpeg_19480_n_293 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_41),
.B1(n_33),
.B2(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_30),
.B1(n_17),
.B2(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_45),
.A2(n_54),
.B1(n_58),
.B2(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_89)
);

NAND2x1_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_31),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_17),
.B1(n_34),
.B2(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_34),
.B1(n_21),
.B2(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_22),
.B1(n_31),
.B2(n_19),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_27),
.B1(n_29),
.B2(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_23),
.B1(n_32),
.B2(n_20),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_42),
.B1(n_31),
.B2(n_35),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_19),
.B1(n_20),
.B2(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_20),
.B1(n_22),
.B2(n_31),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_71),
.B1(n_94),
.B2(n_47),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_91),
.B(n_92),
.Y(n_105)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_78),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_76),
.B1(n_63),
.B2(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_90),
.Y(n_98)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_42),
.C(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_81),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_40),
.C(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_40),
.CI(n_35),
.CON(n_83),
.SN(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_56),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_40),
.B(n_36),
.C(n_31),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_22),
.B1(n_18),
.B2(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_65),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_100),
.A2(n_101),
.B1(n_121),
.B2(n_47),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_112),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_62),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_24),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_123),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_89),
.B1(n_71),
.B2(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_61),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_54),
.B(n_28),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_1),
.B(n_2),
.Y(n_153)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_61),
.B1(n_47),
.B2(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_59),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_92),
.Y(n_127)
);

HAxp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_125),
.CON(n_163),
.SN(n_163)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_132),
.B1(n_137),
.B2(n_102),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_133),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_67),
.B1(n_93),
.B2(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_98),
.B(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_138),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_148),
.B1(n_125),
.B2(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_47),
.B1(n_95),
.B2(n_18),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_18),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_24),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_150),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_117),
.B(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

XOR2x2_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_24),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_4),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_99),
.B(n_118),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_104),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_154),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_28),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_118),
.C(n_100),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_166),
.C(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_124),
.B1(n_125),
.B2(n_105),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_165),
.B1(n_175),
.B2(n_127),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_167),
.B(n_168),
.Y(n_187)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_118),
.C(n_113),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_113),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_170),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_125),
.B(n_113),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_143),
.B(n_140),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_111),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_126),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_125),
.C(n_111),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_102),
.B1(n_110),
.B2(n_108),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_4),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_130),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_4),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_134),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_134),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_192),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_204),
.B(n_185),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_152),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_199),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_142),
.C(n_127),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_210),
.C(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_170),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_129),
.B1(n_142),
.B2(n_141),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_168),
.B1(n_163),
.B2(n_158),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_153),
.B(n_147),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_209),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_146),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_207),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_130),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_5),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_176),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_5),
.C(n_6),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_230),
.B(n_197),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_179),
.B1(n_171),
.B2(n_161),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

AOI22x1_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_167),
.B1(n_183),
.B2(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_161),
.B1(n_178),
.B2(n_180),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_194),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_164),
.C(n_156),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_207),
.C(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_156),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_195),
.CI(n_206),
.CON(n_232),
.SN(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_236),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_188),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_245),
.C(n_213),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_187),
.CI(n_203),
.CON(n_239),
.SN(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_216),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_204),
.B(n_197),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_255),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_245),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_R g251 ( 
.A(n_233),
.B(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_230),
.B1(n_219),
.B2(n_214),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_253),
.B1(n_257),
.B2(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_230),
.B1(n_217),
.B2(n_210),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_231),
.B(n_222),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_228),
.B1(n_189),
.B2(n_194),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_228),
.B1(n_7),
.B2(n_8),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_10),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_268),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_247),
.B(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_263),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_239),
.B(n_232),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_232),
.B(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_234),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_243),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_259),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_257),
.B1(n_253),
.B2(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_11),
.C(n_12),
.Y(n_278)
);

AOI21x1_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_265),
.B(n_264),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_281),
.B(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_268),
.B(n_14),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_13),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_285),
.B(n_13),
.Y(n_289)
);

NAND2x1p5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_13),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_287),
.B(n_288),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_277),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_289),
.A2(n_15),
.B(n_16),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_15),
.B(n_16),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_291),
.Y(n_293)
);


endmodule