module fake_jpeg_25404_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_14),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_34),
.B1(n_16),
.B2(n_21),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_62),
.B1(n_35),
.B2(n_41),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_50),
.B(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_17),
.B1(n_34),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_16),
.B1(n_34),
.B2(n_17),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_34),
.B1(n_16),
.B2(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_27),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_16),
.B1(n_50),
.B2(n_25),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_45),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_38),
.B(n_45),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_40),
.B1(n_35),
.B2(n_33),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_96),
.B1(n_22),
.B2(n_18),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_80),
.B1(n_91),
.B2(n_102),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_56),
.B1(n_24),
.B2(n_48),
.Y(n_127)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_41),
.B1(n_22),
.B2(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_95),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_61),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_44),
.C(n_42),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_45),
.Y(n_107)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_22),
.B1(n_18),
.B2(n_29),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_107),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_56),
.B1(n_53),
.B2(n_52),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_127),
.B1(n_75),
.B2(n_74),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_121),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_86),
.B(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_65),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_130),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_31),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_132),
.B(n_125),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_79),
.B1(n_97),
.B2(n_68),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_143),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_68),
.B1(n_69),
.B2(n_77),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_99),
.B(n_24),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_153),
.B(n_149),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_139),
.A2(n_145),
.B1(n_154),
.B2(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_105),
.B1(n_116),
.B2(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_75),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_146),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_85),
.B1(n_74),
.B2(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_101),
.B1(n_100),
.B2(n_82),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_48),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_88),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_86),
.B1(n_90),
.B2(n_42),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_155),
.B1(n_108),
.B2(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_119),
.B1(n_115),
.B2(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_106),
.B1(n_115),
.B2(n_104),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_104),
.A2(n_44),
.B1(n_42),
.B2(n_45),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_111),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_38),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_44),
.C(n_61),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_120),
.C(n_108),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_89),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_31),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_38),
.A3(n_28),
.B1(n_31),
.B2(n_61),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_180),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_184),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_13),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_178),
.B(n_181),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_139),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_173),
.A2(n_176),
.B(n_190),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_12),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_134),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_153),
.C(n_157),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_155),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_138),
.B(n_28),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_152),
.B1(n_136),
.B2(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_11),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_132),
.B(n_84),
.Y(n_182)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_150),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_196),
.B1(n_28),
.B2(n_20),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_117),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_214),
.B1(n_226),
.B2(n_165),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_172),
.C(n_197),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_174),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_195),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_137),
.B1(n_163),
.B2(n_162),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_204),
.B1(n_210),
.B2(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_147),
.B1(n_156),
.B2(n_117),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_205),
.A2(n_209),
.B(n_219),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_0),
.B(n_1),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_117),
.B1(n_125),
.B2(n_93),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_83),
.B1(n_38),
.B2(n_31),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_31),
.B1(n_28),
.B2(n_20),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_12),
.C(n_11),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_225),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_3),
.B(n_4),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_28),
.B(n_20),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_12),
.B1(n_9),
.B2(n_8),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_166),
.B1(n_183),
.B2(n_184),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_9),
.B1(n_8),
.B2(n_2),
.Y(n_226)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_230),
.A2(n_249),
.B1(n_210),
.B2(n_204),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_176),
.B(n_177),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_209),
.B(n_205),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_193),
.B1(n_164),
.B2(n_171),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_200),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_248),
.C(n_226),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_177),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_241),
.A2(n_242),
.B(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_183),
.B(n_170),
.C(n_172),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_215),
.B(n_221),
.Y(n_266)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_244),
.A2(n_246),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_8),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_0),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_198),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_1),
.C(n_2),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_212),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_255),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_202),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_261),
.B(n_266),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_233),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_264),
.C(n_269),
.Y(n_272)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_201),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_230),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_203),
.C(n_221),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_211),
.C(n_214),
.Y(n_269)
);

FAx1_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_236),
.CI(n_227),
.CON(n_274),
.SN(n_274)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_254),
.B(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_227),
.B1(n_243),
.B2(n_249),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_240),
.C(n_232),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_251),
.C(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_248),
.B(n_229),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_271),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_257),
.A3(n_262),
.B1(n_263),
.B2(n_219),
.C1(n_269),
.C2(n_232),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_297),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

OAI22x1_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_274),
.B1(n_285),
.B2(n_283),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_272),
.B(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_265),
.C(n_259),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_208),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_208),
.C(n_216),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_302),
.B(n_305),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_292),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_250),
.C2(n_307),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_285),
.B(n_274),
.Y(n_307)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_308),
.A3(n_310),
.B(n_300),
.Y(n_313)
);

OA21x2_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_271),
.B(n_275),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_289),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_315),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_5),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_287),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_287),
.C(n_288),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_319),
.B1(n_4),
.B2(n_5),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_324),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_319),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_322),
.B(n_323),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_325),
.B1(n_324),
.B2(n_321),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_6),
.B(n_7),
.Y(n_330)
);


endmodule