module real_jpeg_4805_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_137),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_1),
.A2(n_199),
.B1(n_227),
.B2(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_1),
.A2(n_199),
.B1(n_310),
.B2(n_315),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_1),
.A2(n_199),
.B1(n_216),
.B2(n_408),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_51),
.B1(n_122),
.B2(n_127),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_2),
.A2(n_51),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_4),
.A2(n_41),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_5),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_5),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_5),
.A2(n_78),
.B1(n_187),
.B2(n_191),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_78),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_6),
.A2(n_35),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_7),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_7),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_7),
.A2(n_149),
.B1(n_265),
.B2(n_279),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_7),
.A2(n_149),
.B1(n_310),
.B2(n_315),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_7),
.A2(n_149),
.B1(n_224),
.B2(n_367),
.Y(n_366)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_9),
.Y(n_174)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_9),
.Y(n_340)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_9),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_9),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_155),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_10),
.A2(n_52),
.B1(n_155),
.B2(n_298),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_10),
.A2(n_155),
.B1(n_319),
.B2(n_323),
.Y(n_318)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_11),
.Y(n_140)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_11),
.Y(n_264)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_13),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_13),
.A2(n_267),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_13),
.B(n_305),
.C(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_13),
.B(n_106),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_13),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_13),
.B(n_85),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_13),
.B(n_377),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_14),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_14),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_14),
.Y(n_152)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_14),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_16),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_16),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_16),
.A2(n_52),
.B1(n_116),
.B2(n_181),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_16),
.A2(n_116),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_16),
.A2(n_116),
.B1(n_383),
.B2(n_385),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_242),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_241),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_207),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_20),
.B(n_207),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_161),
.C(n_176),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_21),
.B(n_161),
.CI(n_176),
.CON(n_282),
.SN(n_282)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_86),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_22),
.B(n_87),
.C(n_130),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_23),
.B(n_46),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_37),
.B2(n_40),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_24),
.A2(n_40),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_24),
.A2(n_37),
.B1(n_270),
.B2(n_275),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_24),
.A2(n_309),
.B(n_317),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_24),
.A2(n_267),
.B(n_317),
.Y(n_341)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_25),
.A2(n_186),
.B1(n_193),
.B2(n_194),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_25),
.B(n_318),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_25),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_25),
.A2(n_271),
.B1(n_382),
.B2(n_414),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_30),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_30),
.Y(n_385)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_31),
.Y(n_193)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_33),
.Y(n_192)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_34),
.Y(n_314)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_38),
.B(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_45),
.Y(n_316)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_45),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_77),
.B2(n_85),
.Y(n_46)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_47),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_49),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_49),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_49),
.Y(n_295)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_50),
.Y(n_371)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_55),
.A2(n_77),
.B1(n_85),
.B2(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_55),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_55),
.A2(n_85),
.B1(n_164),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_55),
.B(n_297),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_59),
.Y(n_167)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_59),
.Y(n_228)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_59),
.Y(n_303)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_67),
.Y(n_329)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_68),
.A2(n_327),
.B(n_330),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_70),
.Y(n_305)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_74),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_74),
.Y(n_384)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_83),
.Y(n_109)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_85),
.B(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_130),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_111),
.B1(n_120),
.B2(n_121),
.Y(n_87)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_88),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_88),
.A2(n_120),
.B1(n_278),
.B2(n_407),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_106),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_98),
.B2(n_103),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_91),
.Y(n_392)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_92),
.Y(n_396)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_96),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_96),
.Y(n_378)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_105),
.Y(n_260)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g200 ( 
.A1(n_106),
.A2(n_201),
.B1(n_202),
.B2(n_206),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_106),
.A2(n_201),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_110),
.Y(n_294)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI32xp33_ASAP7_75t_L g389 ( 
.A1(n_117),
.A2(n_168),
.A3(n_376),
.B1(n_390),
.B2(n_393),
.Y(n_389)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_120),
.B(n_203),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_120),
.A2(n_407),
.B(n_410),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g374 ( 
.A1(n_123),
.A2(n_267),
.B(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_126),
.Y(n_265)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_126),
.Y(n_409)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_147),
.B(n_153),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_131),
.A2(n_141),
.B1(n_147),
.B2(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_132),
.B(n_154),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_132),
.A2(n_430),
.B(n_431),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_141),
.B(n_267),
.Y(n_412)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g256 ( 
.A1(n_145),
.A2(n_257),
.A3(n_261),
.B1(n_262),
.B2(n_266),
.Y(n_256)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_153),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_156),
.B(n_267),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_SL g430 ( 
.A1(n_156),
.A2(n_266),
.B(n_267),
.Y(n_430)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_160),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_171),
.B2(n_175),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_171),
.Y(n_232)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_175),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_195),
.C(n_200),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_177),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_185),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_178),
.B(n_185),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_179),
.A2(n_292),
.B(n_296),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_179),
.A2(n_183),
.B1(n_327),
.B2(n_366),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_179),
.A2(n_296),
.B(n_366),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_180),
.A2(n_183),
.B(n_330),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_186),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_197),
.A2(n_240),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_201),
.A2(n_277),
.B(n_281),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_201),
.A2(n_281),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_201),
.B(n_202),
.Y(n_410)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_230),
.B2(n_231),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_220),
.B(n_229),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_221),
.Y(n_229)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g393 ( 
.A(n_226),
.B(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_283),
.B(n_459),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_282),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_245),
.B(n_282),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.C(n_251),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_250),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_251),
.B(n_449),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_276),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_252),
.A2(n_253),
.B1(n_276),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_255),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_268),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_256),
.A2(n_268),
.B1(n_269),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_276),
.Y(n_444)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g462 ( 
.A(n_282),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_437),
.B(n_456),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_418),
.B(n_436),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_398),
.B(n_417),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_360),
.B(n_397),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_333),
.B(n_359),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_307),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_307),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_291),
.A2(n_300),
.B1(n_301),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_291),
.Y(n_357)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_324),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_325),
.C(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_331),
.B2(n_332),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_349),
.B(n_358),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_342),
.B(n_348),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_340),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_347),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B(n_346),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_344),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_346),
.A2(n_381),
.B(n_386),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_356),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_356),
.Y(n_358)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_362),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_379),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_372),
.B2(n_373),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_372),
.C(n_379),
.Y(n_399)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx5_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_389),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_389),
.Y(n_404)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_399),
.B(n_400),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_405),
.B2(n_416),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_404),
.C(n_416),
.Y(n_419)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_412),
.C(n_413),
.Y(n_424)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_419),
.B(n_420),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_427),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_421)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_422),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_424),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_425),
.C(n_427),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_432),
.B2(n_435),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_433),
.C(n_434),
.Y(n_447)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_432),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_451),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_440),
.A2(n_457),
.B(n_458),
.Y(n_456)
);

NOR2x1_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_448),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_448),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.C(n_447),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_445),
.A2(n_446),
.B1(n_447),
.B2(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_447),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_453),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);


endmodule