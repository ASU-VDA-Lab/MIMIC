module fake_jpeg_1381_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_37),
.B1(n_45),
.B2(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_46),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_37),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_40),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_38),
.B1(n_42),
.B2(n_41),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_47),
.B1(n_45),
.B2(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_77),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_43),
.B(n_50),
.C(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_0),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_40),
.C(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_61),
.B(n_68),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_32),
.B(n_30),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_95),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_67),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_79),
.B1(n_82),
.B2(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_81),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_106),
.C(n_5),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_0),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_3),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_17),
.C(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_4),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_92),
.B(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_90),
.B1(n_88),
.B2(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_5),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_29),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_120),
.C(n_27),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_125),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_20),
.C(n_25),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_9),
.B(n_10),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_109),
.B1(n_110),
.B2(n_11),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_120),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_136),
.B1(n_132),
.B2(n_130),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_119),
.B1(n_112),
.B2(n_117),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_133),
.B1(n_128),
.B2(n_15),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_124),
.B(n_115),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_136),
.B(n_14),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_140),
.B(n_142),
.Y(n_144)
);

AOI31xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_140),
.A3(n_22),
.B(n_21),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_23),
.C(n_24),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_12),
.B(n_14),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_15),
.Y(n_148)
);


endmodule