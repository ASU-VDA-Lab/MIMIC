module fake_jpeg_10147_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_240;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_53),
.B1(n_59),
.B2(n_20),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_62),
.B1(n_67),
.B2(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_64),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_34),
.B2(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_27),
.B1(n_17),
.B2(n_30),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_28),
.CON(n_63),
.SN(n_63)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_39),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_87),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_39),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_43),
.B1(n_39),
.B2(n_18),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_43),
.B1(n_36),
.B2(n_41),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_81),
.B(n_30),
.Y(n_98)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_49),
.A3(n_58),
.B1(n_54),
.B2(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_9),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_33),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_58),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_50),
.C(n_37),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_95),
.C(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_40),
.C(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_99),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_29),
.B(n_33),
.Y(n_125)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_101),
.B1(n_91),
.B2(n_74),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_43),
.B1(n_39),
.B2(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_40),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_46),
.B(n_44),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_48),
.B(n_39),
.C(n_58),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_115),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_118),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_41),
.C(n_49),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_44),
.B1(n_54),
.B2(n_35),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_15),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_108),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_143),
.C(n_144),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_128),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_82),
.B(n_77),
.C(n_70),
.D(n_84),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_137),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_131),
.B1(n_133),
.B2(n_142),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_92),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_140),
.B(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_33),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_91),
.B1(n_46),
.B2(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_45),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_106),
.B(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_45),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_29),
.A3(n_44),
.B1(n_33),
.B2(n_31),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_86),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_35),
.B1(n_60),
.B2(n_80),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_44),
.C(n_35),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_44),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_150),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_106),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_154),
.B(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_94),
.C(n_105),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_166),
.C(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_159),
.B(n_161),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_109),
.B1(n_107),
.B2(n_105),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_165),
.B1(n_96),
.B2(n_31),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_109),
.B1(n_102),
.B2(n_103),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_118),
.C(n_35),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_169),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_35),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_140),
.B1(n_128),
.B2(n_137),
.Y(n_170)
);

OAI22x1_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_29),
.B1(n_31),
.B2(n_25),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_60),
.C(n_102),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_25),
.C(n_22),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_127),
.B1(n_140),
.B2(n_130),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_173),
.A2(n_179),
.B1(n_1),
.B2(n_4),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_126),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_126),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_124),
.B1(n_135),
.B2(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_147),
.B1(n_170),
.B2(n_156),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_196),
.B1(n_164),
.B2(n_147),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_192),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_0),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_4),
.B(n_5),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_22),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_25),
.C(n_22),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_16),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_25),
.C(n_0),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_151),
.B1(n_160),
.B2(n_146),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_151),
.B1(n_146),
.B2(n_154),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_166),
.C(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_211),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_207),
.C(n_175),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_157),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_175),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_165),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_16),
.B1(n_2),
.B2(n_4),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_187),
.B(n_173),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_217),
.B(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_216),
.B1(n_187),
.B2(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_193),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_221),
.B(n_224),
.Y(n_234)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_227),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g222 ( 
.A(n_213),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_191),
.B(n_174),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_206),
.C(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_184),
.B(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_232),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_197),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_236),
.C(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_210),
.C(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_174),
.C(n_186),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_209),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_223),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_221),
.C(n_230),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_212),
.B1(n_208),
.B2(n_202),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_219),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_253),
.B(n_255),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_219),
.B(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_240),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_254),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_188),
.B(n_217),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_5),
.B(n_6),
.Y(n_255)
);

NAND2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_244),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_261),
.B(n_262),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_234),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_239),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_247),
.B(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_236),
.C(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_8),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_6),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_260),
.B(n_9),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_265),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_152),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_11),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_275),
.A2(n_273),
.B(n_13),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_13),
.Y(n_277)
);


endmodule