module real_jpeg_26558_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_341, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_341;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_0),
.A2(n_47),
.B1(n_58),
.B2(n_61),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_0),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_1),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_114),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_1),
.A2(n_58),
.B1(n_61),
.B2(n_114),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_114),
.Y(n_252)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_134),
.B(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_4),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_119),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_4),
.A2(n_58),
.B1(n_61),
.B2(n_119),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_25),
.B1(n_52),
.B2(n_53),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_25),
.B1(n_58),
.B2(n_61),
.Y(n_156)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_11),
.B(n_58),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_45),
.B1(n_58),
.B2(n_61),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_36),
.B1(n_58),
.B2(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_11),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_11),
.B(n_30),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_11),
.A2(n_30),
.B(n_160),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_117),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_11),
.B(n_78),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_11),
.A2(n_98),
.B1(n_99),
.B2(n_211),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_15),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_112),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_15),
.A2(n_58),
.B1(n_61),
.B2(n_112),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_339),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_83),
.B(n_337),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_21),
.A2(n_43),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_22),
.A2(n_32),
.B(n_82),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_22),
.A2(n_26),
.B(n_32),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_26),
.B(n_27),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_27),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_23),
.B(n_117),
.CON(n_116),
.SN(n_116)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_32),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_27),
.B(n_30),
.Y(n_131)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_29),
.A2(n_33),
.B1(n_116),
.B2(n_131),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_29),
.A2(n_52),
.A3(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_31),
.A2(n_44),
.B(n_48),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_32),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_48),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_38),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_75),
.C(n_80),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_39),
.A2(n_40),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.C(n_64),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_41),
.A2(n_42),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_43),
.A2(n_48),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_43),
.A2(n_48),
.B1(n_125),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_48),
.B(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_49),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_49),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_49),
.A2(n_64),
.B1(n_305),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_62),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_62),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_50),
.A2(n_57),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_50),
.A2(n_168),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_50),
.A2(n_57),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_50),
.A2(n_57),
.B1(n_167),
.B2(n_186),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_50),
.A2(n_57),
.B1(n_93),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_50),
.A2(n_107),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_53),
.B(n_67),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_53),
.A2(n_56),
.B(n_117),
.C(n_188),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_57),
.B(n_117),
.Y(n_209)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_99),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_61),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_63),
.B(n_108),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_64),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_77),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_73),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_66),
.A2(n_73),
.B1(n_111),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_66),
.A2(n_73),
.B1(n_143),
.B2(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_66),
.B(n_72),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_66),
.A2(n_73),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_71),
.A2(n_78),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_77),
.A2(n_79),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_77),
.A2(n_255),
.B(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_80),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_330),
.B(n_336),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_300),
.A3(n_322),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_281),
.B(n_299),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_259),
.B(n_280),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_148),
.B(n_235),
.C(n_258),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_135),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_89),
.B(n_135),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_120),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_91),
.B(n_104),
.C(n_120),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_92),
.B(n_97),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_94),
.B(n_178),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_98),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_98),
.A2(n_203),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_98),
.A2(n_212),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_103),
.Y(n_102)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_99),
.B(n_117),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_102),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_122),
.B(n_127),
.C(n_129),
.Y(n_256)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_132),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_136),
.A2(n_137),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_141),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_234),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_227),
.B(n_233),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_179),
.B(n_226),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_169),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_152),
.B(n_169),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.C(n_165),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_153),
.A2(n_154),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_198),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_176),
.C(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_220),
.B(n_225),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_199),
.B(n_219),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_182),
.B(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_196),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_207),
.B(n_218),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_205),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_213),
.B(n_217),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_237),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_256),
.B2(n_257),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_247),
.C(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_261),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_279),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_273),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_275),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_275),
.A2(n_293),
.B(n_296),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_297),
.B2(n_298),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_292),
.C(n_298),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B(n_291),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_302),
.C(n_312),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_302),
.B1(n_303),
.B2(n_327),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_291),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_320),
.C(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_313),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule