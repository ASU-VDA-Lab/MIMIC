module fake_jpeg_20232_n_150 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_34),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_8),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_81),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_48),
.B1(n_74),
.B2(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_73),
.B1(n_56),
.B2(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_58),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_67),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_51),
.B1(n_70),
.B2(n_68),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_105),
.B1(n_0),
.B2(n_1),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_81),
.B1(n_78),
.B2(n_82),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_75),
.B1(n_59),
.B2(n_54),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_76),
.B1(n_80),
.B2(n_49),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_17),
.B1(n_46),
.B2(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_63),
.B1(n_74),
.B2(n_69),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_60),
.B1(n_83),
.B2(n_62),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_72),
.B1(n_59),
.B2(n_53),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_66),
.B1(n_64),
.B2(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_118),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_11),
.B1(n_27),
.B2(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_123),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_0),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_20),
.B1(n_43),
.B2(n_31),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_14),
.B1(n_30),
.B2(n_29),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_111),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_132),
.Y(n_135)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_9),
.B(n_23),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_116),
.B1(n_118),
.B2(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_138),
.B1(n_124),
.B2(n_131),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_135),
.B(n_139),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_138),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_128),
.Y(n_144)
);

OAI21x1_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_133),
.B(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_128),
.C(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_13),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

OAI21x1_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_47),
.B(n_6),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_7),
.Y(n_150)
);


endmodule