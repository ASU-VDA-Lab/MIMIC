module fake_jpeg_29392_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_18),
.A2(n_15),
.B1(n_8),
.B2(n_11),
.Y(n_22)
);

OAI32xp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_10),
.A3(n_14),
.B1(n_11),
.B2(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_19),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_17),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.C(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_10),
.Y(n_32)
);

OAI22x1_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_9),
.B1(n_14),
.B2(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_24),
.B(n_37),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_44),
.B1(n_15),
.B2(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_34),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_37),
.B(n_5),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_41),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_45),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_15),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_4),
.Y(n_56)
);


endmodule