module fake_jpeg_487_n_200 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_200);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_69),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_69),
.B1(n_62),
.B2(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_62),
.B1(n_68),
.B2(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_73),
.B1(n_71),
.B2(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_66),
.C(n_59),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_59),
.Y(n_119)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_65),
.B1(n_51),
.B2(n_54),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_72),
.B(n_58),
.Y(n_116)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_64),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_71),
.B1(n_60),
.B2(n_61),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_109),
.B1(n_72),
.B2(n_53),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_78),
.B1(n_75),
.B2(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_81),
.B1(n_80),
.B2(n_78),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_116),
.B1(n_125),
.B2(n_126),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_94),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_49),
.B(n_70),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_93),
.B(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_23),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_78),
.B1(n_75),
.B2(n_51),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_75),
.B1(n_64),
.B2(n_50),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_28),
.B1(n_44),
.B2(n_43),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_138),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_29),
.B(n_40),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_96),
.C(n_98),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_137),
.C(n_140),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_24),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_26),
.B1(n_47),
.B2(n_46),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_149),
.B1(n_150),
.B2(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_19),
.C(n_45),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_146),
.B(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_0),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_2),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_148),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_4),
.B(n_5),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_5),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_22),
.C(n_42),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_12),
.C(n_14),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_6),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_35),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_110),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_166),
.B1(n_168),
.B2(n_14),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_9),
.B(n_11),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_30),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_167),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_12),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_153),
.B1(n_152),
.B2(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_172),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_48),
.A3(n_27),
.B1(n_31),
.B2(n_39),
.C(n_36),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_173),
.B1(n_164),
.B2(n_162),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_182),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_163),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_185),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_160),
.C(n_158),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_186),
.C(n_176),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_154),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_159),
.C(n_167),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_189),
.C(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_179),
.C(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_175),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_33),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_191),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_188),
.B(n_194),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.C(n_17),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_198),
.A2(n_16),
.B(n_18),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_18),
.Y(n_200)
);


endmodule