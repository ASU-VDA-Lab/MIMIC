module fake_jpeg_29883_n_358 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_0),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_8),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_31),
.B1(n_24),
.B2(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_69),
.B1(n_78),
.B2(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_25),
.B1(n_18),
.B2(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_30),
.B1(n_29),
.B2(n_20),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_32),
.C(n_31),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_77),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_40),
.B(n_47),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_20),
.B(n_26),
.C(n_50),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_25),
.B1(n_35),
.B2(n_23),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_72),
.B1(n_53),
.B2(n_41),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_24),
.B1(n_34),
.B2(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_25),
.B1(n_35),
.B2(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_38),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_18),
.B(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_24),
.B1(n_34),
.B2(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_79),
.B(n_96),
.Y(n_130)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_90),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_67),
.Y(n_82)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_53),
.B1(n_49),
.B2(n_41),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_107),
.B1(n_76),
.B2(n_67),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_99),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_85),
.Y(n_135)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_33),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_35),
.B1(n_23),
.B2(n_29),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_106),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_67),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_22),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_63),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_45),
.B1(n_44),
.B2(n_26),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_65),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_51),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_50),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_62),
.B(n_9),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_30),
.C(n_56),
.Y(n_133)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_144),
.B1(n_113),
.B2(n_92),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_58),
.B1(n_76),
.B2(n_73),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_124),
.B1(n_128),
.B2(n_107),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_86),
.B(n_79),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_97),
.B(n_111),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_76),
.B1(n_73),
.B2(n_56),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_102),
.B1(n_95),
.B2(n_88),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_86),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_80),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_56),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_0),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_48),
.B1(n_9),
.B2(n_10),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_147),
.B(n_158),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_149),
.B(n_151),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_101),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_164),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_96),
.B(n_80),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_153),
.A2(n_125),
.B(n_127),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_96),
.B(n_81),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_175),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_93),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_155),
.B(n_156),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_110),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_109),
.B(n_105),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_134),
.B(n_137),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_82),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_166),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_123),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_114),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_117),
.B1(n_118),
.B2(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_87),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_91),
.B1(n_112),
.B2(n_99),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_91),
.B1(n_99),
.B2(n_48),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_134),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_87),
.B(n_48),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_176),
.B(n_121),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_128),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_131),
.B(n_148),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_178),
.A2(n_187),
.B(n_189),
.C(n_197),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_139),
.C(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_186),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_207),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_131),
.B(n_116),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_139),
.B(n_135),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_135),
.B(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_194),
.B(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_118),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_202),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_165),
.B(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_205),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_133),
.C(n_119),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_167),
.B(n_121),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_125),
.B(n_116),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_210),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_120),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_124),
.C(n_132),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g209 ( 
.A1(n_151),
.A2(n_132),
.B1(n_141),
.B2(n_127),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_170),
.B1(n_174),
.B2(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_232),
.B1(n_235),
.B2(n_183),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_190),
.A2(n_169),
.B1(n_161),
.B2(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_186),
.B1(n_196),
.B2(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_191),
.B(n_172),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_226),
.B(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_157),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_176),
.B1(n_161),
.B2(n_152),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_125),
.B1(n_138),
.B2(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_10),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

OA21x2_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_138),
.B(n_8),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_208),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_1),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_189),
.B(n_180),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_266),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_179),
.C(n_204),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_263),
.C(n_228),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_256),
.B1(n_217),
.B2(n_234),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_197),
.B(n_193),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_183),
.B1(n_187),
.B2(n_206),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_255),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_178),
.B(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_261),
.Y(n_269)
);

OAI22x1_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_178),
.B1(n_209),
.B2(n_194),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_215),
.A2(n_195),
.B1(n_178),
.B2(n_199),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_232),
.B1(n_234),
.B2(n_213),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_202),
.C(n_201),
.Y(n_263)
);

XOR2x2_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_209),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_219),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_214),
.A2(n_195),
.B(n_138),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_280),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_276),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_277),
.B(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_218),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_229),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_229),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_254),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_282),
.B(n_251),
.CI(n_11),
.CON(n_301),
.SN(n_301)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_234),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_258),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_221),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_259),
.B1(n_264),
.B2(n_248),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_211),
.Y(n_288)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_264),
.C(n_253),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_287),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_266),
.C(n_242),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_265),
.B1(n_241),
.B2(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_250),
.B(n_257),
.Y(n_295)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_249),
.B1(n_252),
.B2(n_247),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_252),
.B1(n_258),
.B2(n_244),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_301),
.Y(n_314)
);

NOR2x1p5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_257),
.Y(n_298)
);

NOR2x1p5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_5),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_251),
.C(n_11),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_304),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_7),
.C(n_16),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_313),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_267),
.B(n_269),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_278),
.B(n_283),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_292),
.B(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_7),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_14),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_6),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_11),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_321),
.Y(n_329)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_299),
.C(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_327),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_324),
.B(n_333),
.Y(n_342)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_299),
.C(n_293),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_301),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_332),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_312),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_309),
.B(n_304),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_334),
.B(n_335),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_314),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_339),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_298),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g346 ( 
.A1(n_338),
.A2(n_328),
.A3(n_14),
.B1(n_5),
.B2(n_15),
.C1(n_17),
.C2(n_3),
.Y(n_346)
);

BUFx12_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_311),
.B(n_325),
.C(n_333),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_343),
.A2(n_1),
.B(n_2),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_348),
.B(n_349),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_15),
.C(n_17),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_347),
.B(n_334),
.C(n_342),
.Y(n_351)
);

OAI21x1_ASAP7_75t_SL g348 ( 
.A1(n_339),
.A2(n_15),
.B(n_17),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_1),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_350),
.A2(n_2),
.A3(n_3),
.B1(n_341),
.B2(n_342),
.C1(n_344),
.C2(n_345),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_354),
.Y(n_356)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_353),
.Y(n_355)
);

OA21x2_ASAP7_75t_SL g354 ( 
.A1(n_347),
.A2(n_2),
.B(n_3),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_352),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_355),
.Y(n_358)
);


endmodule