module fake_netlist_6_2554_n_3965 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_865, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_839, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_777, n_407, n_450, n_103, n_808, n_867, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_860, n_481, n_788, n_819, n_821, n_325, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_864, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_817, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_846, n_501, n_841, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3965);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_865;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_839;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_821;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_864;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_846;
input n_501;
input n_841;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3965;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_2576;
wire n_1234;
wire n_1458;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_3773;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_2260;
wire n_3222;
wire n_1387;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_2557;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1009;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_1285;
wire n_3946;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1143;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_2739;
wire n_2480;
wire n_1300;
wire n_3023;
wire n_1541;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_2212;
wire n_3929;
wire n_3494;
wire n_3048;
wire n_3063;
wire n_2418;
wire n_2864;
wire n_2729;
wire n_1163;
wire n_1455;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_2873;
wire n_1820;
wire n_1345;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_1054;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_3943;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_3728;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1162;
wire n_1530;
wire n_3798;
wire n_939;
wire n_3488;
wire n_2811;
wire n_1543;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_3857;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1605;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_3927;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_2714;
wire n_3092;
wire n_2245;
wire n_3055;
wire n_1289;
wire n_3492;
wire n_3895;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_3861;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_1801;
wire n_2347;
wire n_1886;
wire n_928;
wire n_2092;
wire n_1214;
wire n_1654;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_2963;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_3873;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_2943;
wire n_1294;
wire n_1420;
wire n_3780;
wire n_3696;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_3337;
wire n_1465;
wire n_3450;
wire n_3431;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1627;
wire n_1295;
wire n_1164;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_1128;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_2535;
wire n_1026;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_2693;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_2767;
wire n_3793;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_1139;
wire n_3922;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3426;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_3580;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_2134;
wire n_1176;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_2958;
wire n_1577;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_947;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_1299;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3893;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_2127;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_3201;
wire n_1284;
wire n_3633;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_2354;
wire n_1398;
wire n_2682;
wire n_884;
wire n_1048;
wire n_1201;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_2581;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_3641;
wire n_1837;
wire n_964;
wire n_2218;
wire n_1314;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_2416;
wire n_1427;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3909;
wire n_3944;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_3364;
wire n_2929;
wire n_1597;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_1533;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_1745;
wire n_914;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_1459;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_2720;
wire n_1520;
wire n_3126;
wire n_2159;
wire n_906;
wire n_2289;
wire n_2315;
wire n_1733;
wire n_1077;
wire n_2863;
wire n_1390;
wire n_3299;
wire n_1419;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_3917;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_3870;
wire n_1696;
wire n_2829;
wire n_2181;
wire n_1594;
wire n_1995;
wire n_3751;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_3886;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_1037;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_2716;
wire n_3249;
wire n_1320;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_3137;
wire n_3382;
wire n_1535;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_3819;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2373;
wire n_2120;
wire n_2050;
wire n_1472;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_2376;
wire n_1405;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_2670;
wire n_1332;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_2258;
wire n_1485;
wire n_1544;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1475;
wire n_1235;
wire n_1318;
wire n_1229;
wire n_2759;
wire n_3457;
wire n_2945;
wire n_3061;
wire n_3517;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3613;
wire n_3483;
wire n_2128;
wire n_1650;
wire n_1045;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_2398;
wire n_1725;
wire n_1928;
wire n_1559;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3818;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2885;
wire n_3776;
wire n_3711;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_3511;
wire n_2054;
wire n_876;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_1023;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1378;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_2584;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_3473;
wire n_895;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_2465;
wire n_1112;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1737;
wire n_1464;
wire n_2430;
wire n_3486;
wire n_1414;
wire n_3584;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_2743;
wire n_3962;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_990;
wire n_1821;
wire n_1500;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_904;
wire n_1253;
wire n_2242;
wire n_1266;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_2609;
wire n_1161;
wire n_2802;
wire n_1085;
wire n_3796;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1156;
wire n_1362;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_2033;
wire n_3086;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2071;
wire n_1144;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_2805;
wire n_1301;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_3925;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_2221;
wire n_1170;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_3274;
wire n_2899;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g875 ( 
.A(n_224),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_543),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_657),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_492),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_645),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_360),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_220),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_701),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_851),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_613),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_410),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_353),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_850),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_861),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_815),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_780),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_733),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_782),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_602),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_758),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_355),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_271),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_88),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_859),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_673),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_246),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_582),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_43),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_61),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_14),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_322),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_136),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_830),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_256),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_668),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_314),
.Y(n_910)
);

BUFx8_ASAP7_75t_SL g911 ( 
.A(n_677),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_609),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_203),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_502),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_681),
.Y(n_915)
);

BUFx10_ASAP7_75t_L g916 ( 
.A(n_420),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_273),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_120),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_17),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_574),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_573),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_647),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_98),
.Y(n_923)
);

BUFx10_ASAP7_75t_L g924 ( 
.A(n_710),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_258),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_779),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_215),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_565),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_128),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_365),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_869),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_687),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_694),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_307),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_649),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_233),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_686),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_312),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_12),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_707),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_391),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_106),
.Y(n_942)
);

CKINVDCx14_ASAP7_75t_R g943 ( 
.A(n_565),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_808),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_647),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_762),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_271),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_97),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_482),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_21),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_521),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_12),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_784),
.Y(n_953)
);

BUFx10_ASAP7_75t_L g954 ( 
.A(n_603),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_500),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_161),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_235),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_44),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_652),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_515),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_728),
.Y(n_961)
);

BUFx10_ASAP7_75t_L g962 ( 
.A(n_826),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_590),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_644),
.Y(n_964)
);

BUFx10_ASAP7_75t_L g965 ( 
.A(n_333),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_638),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_817),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_839),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_99),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_643),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_658),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_637),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_860),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_790),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_730),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_79),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_117),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_213),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_601),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_278),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_470),
.Y(n_981)
);

BUFx5_ASAP7_75t_L g982 ( 
.A(n_695),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_679),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_203),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_181),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_121),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_64),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_375),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_381),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_863),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_770),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_757),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_571),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_158),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_585),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_594),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_279),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_765),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_759),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_446),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_834),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_675),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_185),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_814),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_47),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_618),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_366),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_816),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_781),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_349),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_270),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_490),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_242),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_777),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_843),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_368),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_666),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_354),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_601),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_396),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_853),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_590),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_418),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_587),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_676),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_147),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_735),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_804),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_403),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_572),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_498),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_862),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_767),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_403),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_446),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_665),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_364),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_136),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_600),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_120),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_865),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_452),
.Y(n_1042)
);

INVxp67_ASAP7_75t_SL g1043 ( 
.A(n_631),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_579),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_46),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_455),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_416),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_477),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_828),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_150),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_766),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_651),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_871),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_696),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_327),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_584),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_362),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_604),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_56),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_569),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_365),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_252),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_304),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_751),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_764),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_708),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_592),
.Y(n_1067)
);

BUFx5_ASAP7_75t_L g1068 ( 
.A(n_477),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_752),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_106),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_745),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_400),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_835),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_713),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_597),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_322),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_709),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_470),
.Y(n_1078)
);

BUFx10_ASAP7_75t_L g1079 ( 
.A(n_545),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_441),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_612),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_249),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_704),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_389),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_584),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_640),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_645),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_768),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_632),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_39),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_129),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_670),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_753),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_87),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_812),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_818),
.Y(n_1096)
);

BUFx10_ASAP7_75t_L g1097 ( 
.A(n_786),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_452),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_375),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_778),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_473),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_114),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_793),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_426),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_606),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_488),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_107),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_534),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_721),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_60),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_29),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_392),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_726),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_621),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_130),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_289),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_566),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_212),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_272),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_275),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_743),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_663),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_41),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_212),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_577),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_556),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_190),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_772),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_719),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_678),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_115),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_855),
.Y(n_1133)
);

BUFx5_ASAP7_75t_L g1134 ( 
.A(n_304),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_605),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_625),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_342),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_671),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_700),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_827),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_874),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_272),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_791),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_639),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_545),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_842),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_168),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_390),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_336),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_298),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_632),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_650),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_724),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_761),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_542),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_371),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_4),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_648),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_792),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_124),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_626),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_363),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_160),
.Y(n_1163)
);

BUFx2_ASAP7_75t_SL g1164 ( 
.A(n_661),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_284),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_369),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_831),
.Y(n_1167)
);

CKINVDCx16_ASAP7_75t_R g1168 ( 
.A(n_544),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_824),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_356),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_685),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_180),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_313),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_168),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_691),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_396),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_669),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_688),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_567),
.Y(n_1179)
);

CKINVDCx16_ASAP7_75t_R g1180 ( 
.A(n_663),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_674),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_127),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_420),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_586),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_539),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_866),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_594),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_787),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_837),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_562),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_187),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_233),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_518),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_598),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_819),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_849),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_794),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_825),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_123),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_552),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_241),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_467),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_608),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_513),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_612),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_327),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_697),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_157),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_339),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_275),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_539),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_18),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_146),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_583),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_254),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_736),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_711),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_660),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_744),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_376),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_162),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_616),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_802),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_180),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_723),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_654),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_7),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_737),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_395),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_846),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_455),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_226),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_672),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_384),
.Y(n_1234)
);

BUFx10_ASAP7_75t_L g1235 ( 
.A(n_591),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_185),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_216),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_18),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_245),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_771),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_279),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_306),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_561),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_821),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_11),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_178),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_684),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_702),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_750),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_178),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_642),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_811),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_252),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_288),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_368),
.Y(n_1255)
);

BUFx10_ASAP7_75t_L g1256 ( 
.A(n_399),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_49),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_580),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_130),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_472),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_407),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_800),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_563),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_659),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_836),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_3),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_615),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_346),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_98),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_774),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_313),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_623),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_262),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_183),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_256),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_172),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_205),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_62),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_240),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_689),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_661),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_806),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_444),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_514),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_595),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_731),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_575),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_799),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_610),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_509),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_641),
.Y(n_1291)
);

CKINVDCx16_ASAP7_75t_R g1292 ( 
.A(n_653),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_421),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_653),
.Y(n_1294)
);

CKINVDCx16_ASAP7_75t_R g1295 ( 
.A(n_116),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_746),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_712),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_867),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_785),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_123),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_186),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_596),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_589),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_720),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_228),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_845),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_847),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_175),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_586),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_393),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_492),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_463),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_311),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_167),
.Y(n_1314)
);

BUFx8_ASAP7_75t_SL g1315 ( 
.A(n_14),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_49),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_630),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_303),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_748),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_53),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_625),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_237),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_292),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_562),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_154),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_628),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_635),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_634),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_833),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_108),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_664),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_656),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_324),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_381),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_742),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_775),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_35),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_540),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_810),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_182),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_487),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_665),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_844),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_113),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_353),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_426),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_258),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_656),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_109),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_485),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_56),
.Y(n_1351)
);

BUFx8_ASAP7_75t_SL g1352 ( 
.A(n_348),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_100),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_795),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_706),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_773),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_128),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_749),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_754),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_522),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_196),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_78),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_521),
.Y(n_1363)
);

BUFx10_ASAP7_75t_L g1364 ( 
.A(n_614),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_129),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_832),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_153),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_738),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_789),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_46),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_870),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_690),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_505),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_511),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_221),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_698),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_312),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_643),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_763),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_538),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_646),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_523),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_822),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_829),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_809),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_617),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_137),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_415),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_237),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_440),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_854),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_717),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_722),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_542),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_424),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_803),
.Y(n_1396)
);

CKINVDCx16_ASAP7_75t_R g1397 ( 
.A(n_619),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_577),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_421),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_349),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_872),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_86),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_174),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_715),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_624),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_121),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_6),
.Y(n_1407)
);

BUFx5_ASAP7_75t_L g1408 ( 
.A(n_118),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_308),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_868),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_611),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_483),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_602),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_311),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_138),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_422),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_32),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_504),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_618),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_841),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_165),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_359),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_740),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_42),
.Y(n_1424)
);

INVxp33_ASAP7_75t_SL g1425 ( 
.A(n_568),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_116),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_55),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_838),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_633),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_219),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_622),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_428),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_338),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_354),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_629),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_35),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_411),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_436),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_658),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_807),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_23),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_613),
.Y(n_1442)
);

BUFx10_ASAP7_75t_L g1443 ( 
.A(n_693),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_747),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_44),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_682),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_156),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_788),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_718),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_729),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_649),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_627),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_650),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_848),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_639),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_351),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_607),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_397),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_769),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_756),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_437),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_274),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_798),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_801),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_576),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_570),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_541),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_755),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_140),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_640),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_655),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_620),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_38),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_371),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_588),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_504),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_216),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_760),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_303),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_524),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_692),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_352),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_820),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_451),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_456),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_560),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_362),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_182),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_165),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_143),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_783),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_84),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_593),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_840),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_572),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_578),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_122),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_703),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_489),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_503),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_714),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_633),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_631),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_331),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_300),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_621),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_417),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_416),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_141),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_705),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_716),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_858),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_805),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_725),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_727),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_615),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_291),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_227),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_338),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_797),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_660),
.Y(n_1522)
);

CKINVDCx14_ASAP7_75t_R g1523 ( 
.A(n_95),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_302),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_525),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_133),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_662),
.Y(n_1527)
);

CKINVDCx14_ASAP7_75t_R g1528 ( 
.A(n_104),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_581),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_823),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_206),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_582),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_501),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_253),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_440),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_680),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_240),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_267),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_535),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_597),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_207),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_219),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_132),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_290),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_564),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_638),
.Y(n_1546)
);

BUFx10_ASAP7_75t_L g1547 ( 
.A(n_557),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_599),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_683),
.Y(n_1549)
);

CKINVDCx11_ASAP7_75t_R g1550 ( 
.A(n_520),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_796),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_324),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_10),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_852),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_532),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_307),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_78),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_51),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_277),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_459),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_6),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_856),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_813),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_864),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_741),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_432),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_776),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_732),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_84),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_449),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_288),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_739),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_21),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_119),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_857),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_82),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_192),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_873),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_636),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_286),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_247),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_734),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_443),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_555),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_8),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_382),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_377),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_220),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_183),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_591),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_347),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_435),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_16),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_337),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_201),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_667),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_664),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_699),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1068),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1068),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1315),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1068),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1068),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1068),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1068),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1229),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1068),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1550),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1134),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1329),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1315),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1134),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1134),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1550),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1134),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1134),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1134),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1408),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1408),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1408),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1408),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1408),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1408),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1408),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1352),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_897),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1358),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_881),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_937),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1352),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_955),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_995),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_881),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_995),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_882),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_974),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_944),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1011),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1011),
.Y(n_1639)
);

CKINVDCx16_ASAP7_75t_R g1640 ( 
.A(n_1156),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1237),
.Y(n_1641)
);

INVxp33_ASAP7_75t_SL g1642 ( 
.A(n_1442),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1017),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1017),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1022),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_998),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1460),
.Y(n_1647)
);

CKINVDCx16_ASAP7_75t_R g1648 ( 
.A(n_1168),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1070),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1130),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1070),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1101),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1101),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1109),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1578),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1265),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1209),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1180),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_932),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1209),
.Y(n_1660)
);

INVxp33_ASAP7_75t_SL g1661 ( 
.A(n_1531),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_883),
.Y(n_1662)
);

INVxp33_ASAP7_75t_L g1663 ( 
.A(n_1566),
.Y(n_1663)
);

CKINVDCx16_ASAP7_75t_R g1664 ( 
.A(n_1292),
.Y(n_1664)
);

INVxp33_ASAP7_75t_SL g1665 ( 
.A(n_1573),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1122),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_891),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_898),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1375),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1375),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1412),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1513),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1412),
.Y(n_1673)
);

INVxp67_ASAP7_75t_SL g1674 ( 
.A(n_1516),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1508),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_974),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1508),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1590),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_1371),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1592),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1592),
.Y(n_1681)
);

INVxp33_ASAP7_75t_SL g1682 ( 
.A(n_879),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1594),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_881),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_907),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1594),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_881),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_885),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_885),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_885),
.Y(n_1690)
);

INVxp67_ASAP7_75t_SL g1691 ( 
.A(n_1001),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1024),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1024),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1295),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1024),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1024),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_915),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1040),
.Y(n_1698)
);

CKINVDCx14_ASAP7_75t_R g1699 ( 
.A(n_943),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1040),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1040),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1001),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_916),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1336),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1040),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_1336),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1063),
.Y(n_1707)
);

CKINVDCx14_ASAP7_75t_R g1708 ( 
.A(n_943),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_911),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1063),
.Y(n_1710)
);

INVxp33_ASAP7_75t_L g1711 ( 
.A(n_875),
.Y(n_1711)
);

CKINVDCx20_ASAP7_75t_R g1712 ( 
.A(n_911),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1063),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1142),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_926),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1028),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1142),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1142),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1142),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1312),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1312),
.Y(n_1721)
);

CKINVDCx16_ASAP7_75t_R g1722 ( 
.A(n_1397),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1312),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1312),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1386),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_946),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1386),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1386),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1356),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_953),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1386),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1430),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1430),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1430),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1356),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1430),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_877),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_878),
.Y(n_1738)
);

CKINVDCx20_ASAP7_75t_R g1739 ( 
.A(n_1523),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_SL g1740 ( 
.A(n_947),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1587),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1468),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_947),
.Y(n_1743)
);

CKINVDCx16_ASAP7_75t_R g1744 ( 
.A(n_1523),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1468),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1588),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_982),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_961),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_968),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1549),
.Y(n_1750)
);

CKINVDCx16_ASAP7_75t_R g1751 ( 
.A(n_1528),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1586),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_975),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1596),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1549),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_884),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_983),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_902),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_903),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_932),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_887),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1581),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1528),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1583),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_904),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_990),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_910),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_991),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_999),
.Y(n_1769)
);

BUFx12f_ASAP7_75t_L g1770 ( 
.A(n_1625),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1628),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1633),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1684),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1658),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1635),
.B(n_1228),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1689),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1662),
.B(n_1297),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1699),
.B(n_924),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1599),
.A2(n_1602),
.B(n_1600),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1659),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1682),
.B(n_1425),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1667),
.B(n_889),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1668),
.B(n_889),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1661),
.A2(n_1020),
.B1(n_1147),
.B2(n_1012),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1739),
.A2(n_1333),
.B1(n_918),
.B2(n_952),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1672),
.B(n_1195),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1698),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1708),
.B(n_924),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1659),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1674),
.B(n_1676),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1744),
.B(n_924),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1701),
.Y(n_1792)
);

OAI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1603),
.A2(n_1092),
.B(n_992),
.Y(n_1793)
);

BUFx12f_ASAP7_75t_L g1794 ( 
.A(n_1608),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1636),
.Y(n_1795)
);

CKINVDCx11_ASAP7_75t_R g1796 ( 
.A(n_1709),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1687),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1751),
.B(n_962),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1685),
.B(n_1092),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1688),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1690),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1659),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1692),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1697),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1693),
.Y(n_1805)
);

INVx6_ASAP7_75t_L g1806 ( 
.A(n_1640),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1695),
.Y(n_1807)
);

BUFx8_ASAP7_75t_L g1808 ( 
.A(n_1740),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1696),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1700),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1694),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1760),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1705),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1691),
.B(n_1702),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1716),
.B(n_1735),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1665),
.A2(n_1485),
.B1(n_1043),
.B2(n_886),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1760),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1729),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1715),
.B(n_1726),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1707),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1730),
.B(n_1196),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1710),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1713),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1745),
.B(n_1750),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1742),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1714),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1642),
.A2(n_895),
.B1(n_900),
.B2(n_893),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1717),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_SL g1829 ( 
.A(n_1763),
.B(n_962),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1626),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1760),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1648),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1718),
.Y(n_1833)
);

CKINVDCx11_ASAP7_75t_R g1834 ( 
.A(n_1712),
.Y(n_1834)
);

OA21x2_ASAP7_75t_L g1835 ( 
.A1(n_1604),
.A2(n_890),
.B(n_888),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1605),
.A2(n_1198),
.B(n_1196),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1719),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1720),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1721),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1723),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1724),
.B(n_892),
.Y(n_1841)
);

INVx5_ASAP7_75t_L g1842 ( 
.A(n_1664),
.Y(n_1842)
);

INVx5_ASAP7_75t_L g1843 ( 
.A(n_1722),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1725),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1727),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1607),
.A2(n_1449),
.B(n_1270),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1728),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1731),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1748),
.B(n_1270),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1732),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1609),
.A2(n_899),
.B(n_894),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1733),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1734),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1752),
.B(n_962),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1736),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1749),
.B(n_1449),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1610),
.A2(n_920),
.B1(n_925),
.B2(n_921),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1753),
.B(n_1298),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1737),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1738),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1741),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1746),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1612),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1754),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1755),
.B(n_1304),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1764),
.B(n_1761),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1757),
.B(n_1568),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1663),
.A2(n_929),
.B1(n_935),
.B2(n_927),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1627),
.A2(n_936),
.B1(n_939),
.B2(n_938),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1647),
.B(n_1655),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1613),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1767),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1766),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1615),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1756),
.Y(n_1875)
);

BUFx12f_ASAP7_75t_L g1876 ( 
.A(n_1614),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_L g1877 ( 
.A(n_1616),
.B(n_909),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1617),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1758),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1759),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1762),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1618),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_SL g1883 ( 
.A(n_1601),
.B(n_967),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1765),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1619),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1620),
.Y(n_1886)
);

CKINVDCx14_ASAP7_75t_R g1887 ( 
.A(n_1629),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1621),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1606),
.B(n_1641),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1622),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1768),
.B(n_1568),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1623),
.Y(n_1892)
);

INVx4_ASAP7_75t_L g1893 ( 
.A(n_1769),
.Y(n_1893)
);

NOR2x1_ASAP7_75t_L g1894 ( 
.A(n_1624),
.B(n_931),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1631),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1632),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1747),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1634),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1703),
.A2(n_942),
.B1(n_949),
.B2(n_945),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1638),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1639),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1643),
.B(n_933),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1644),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1645),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1649),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1651),
.B(n_940),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1711),
.B(n_967),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1652),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1653),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1743),
.B(n_1307),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1654),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1657),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1611),
.Y(n_1913)
);

INVx5_ASAP7_75t_L g1914 ( 
.A(n_1740),
.Y(n_1914)
);

INVx4_ASAP7_75t_L g1915 ( 
.A(n_1630),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1660),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1669),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1670),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1671),
.B(n_973),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1673),
.B(n_1675),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1677),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1678),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1680),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1681),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1683),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1686),
.Y(n_1926)
);

INVx4_ASAP7_75t_L g1927 ( 
.A(n_1637),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1646),
.Y(n_1928)
);

AOI22x1_ASAP7_75t_SL g1929 ( 
.A1(n_1706),
.A2(n_1042),
.B1(n_1135),
.B2(n_908),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1650),
.Y(n_1930)
);

CKINVDCx16_ASAP7_75t_R g1931 ( 
.A(n_1656),
.Y(n_1931)
);

BUFx12f_ASAP7_75t_L g1932 ( 
.A(n_1679),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1666),
.B(n_1354),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1628),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1682),
.B(n_1530),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1628),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1661),
.A2(n_958),
.B1(n_959),
.B2(n_956),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1659),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1628),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1661),
.A2(n_963),
.B1(n_964),
.B2(n_960),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1666),
.B(n_1582),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1628),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1658),
.B(n_901),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1661),
.A2(n_969),
.B1(n_970),
.B2(n_966),
.Y(n_1944)
);

AND2x6_ASAP7_75t_L g1945 ( 
.A(n_1626),
.B(n_906),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1699),
.B(n_967),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1636),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1752),
.Y(n_1948)
);

BUFx12f_ASAP7_75t_L g1949 ( 
.A(n_1625),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1628),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1661),
.A2(n_972),
.B1(n_977),
.B2(n_976),
.Y(n_1951)
);

OA21x2_ASAP7_75t_L g1952 ( 
.A1(n_1599),
.A2(n_1004),
.B(n_1002),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1659),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1739),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1628),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1628),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1659),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1628),
.Y(n_1958)
);

OA21x2_ASAP7_75t_L g1959 ( 
.A1(n_1599),
.A2(n_1049),
.B(n_1033),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1628),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1628),
.Y(n_1961)
);

BUFx8_ASAP7_75t_L g1962 ( 
.A(n_1740),
.Y(n_1962)
);

CKINVDCx11_ASAP7_75t_R g1963 ( 
.A(n_1709),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1659),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1628),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1599),
.A2(n_1054),
.B(n_1053),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1661),
.A2(n_978),
.B1(n_984),
.B2(n_981),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1628),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1628),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1636),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1666),
.B(n_1444),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1628),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1628),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1635),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1659),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1682),
.B(n_1065),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1628),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1628),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1628),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1659),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1635),
.B(n_1069),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1628),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1636),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1682),
.B(n_1073),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1635),
.B(n_1077),
.Y(n_1985)
);

AOI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1661),
.A2(n_985),
.B1(n_988),
.B2(n_987),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1661),
.A2(n_993),
.B1(n_997),
.B2(n_994),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1635),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1628),
.Y(n_1989)
);

BUFx12f_ASAP7_75t_L g1990 ( 
.A(n_1625),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1659),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1628),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1635),
.B(n_1093),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1628),
.Y(n_1994)
);

OAI21x1_ASAP7_75t_L g1995 ( 
.A1(n_1599),
.A2(n_1096),
.B(n_1095),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1666),
.B(n_1143),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1744),
.B(n_1097),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1628),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1628),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1659),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1659),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1635),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1628),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1628),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_L g2005 ( 
.A1(n_1599),
.A2(n_1171),
.B(n_1146),
.Y(n_2005)
);

BUFx2_ASAP7_75t_L g2006 ( 
.A(n_1739),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1628),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1628),
.Y(n_2008)
);

BUFx12f_ASAP7_75t_L g2009 ( 
.A(n_1625),
.Y(n_2009)
);

BUFx3_ASAP7_75t_L g2010 ( 
.A(n_1636),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1659),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1658),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1635),
.B(n_1188),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1628),
.Y(n_2014)
);

AND2x6_ASAP7_75t_L g2015 ( 
.A(n_1626),
.B(n_950),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1658),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1636),
.Y(n_2017)
);

INVx5_ASAP7_75t_L g2018 ( 
.A(n_1659),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1628),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1699),
.B(n_1097),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1628),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1628),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1628),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1628),
.Y(n_2024)
);

NAND2x1p5_ASAP7_75t_L g2025 ( 
.A(n_1636),
.B(n_932),
.Y(n_2025)
);

CKINVDCx16_ASAP7_75t_R g2026 ( 
.A(n_1744),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1699),
.B(n_1097),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1661),
.A2(n_1019),
.B1(n_1031),
.B2(n_1030),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1666),
.B(n_1189),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1699),
.B(n_1114),
.Y(n_2030)
);

INVx6_ASAP7_75t_L g2031 ( 
.A(n_1640),
.Y(n_2031)
);

INVx6_ASAP7_75t_L g2032 ( 
.A(n_1640),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1659),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1628),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1628),
.Y(n_2035)
);

OA21x2_ASAP7_75t_L g2036 ( 
.A1(n_1599),
.A2(n_1244),
.B(n_1219),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1666),
.B(n_1247),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1699),
.B(n_1114),
.Y(n_2038)
);

BUFx3_ASAP7_75t_L g2039 ( 
.A(n_1636),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1599),
.A2(n_1335),
.B(n_1252),
.Y(n_2040)
);

INVx4_ASAP7_75t_L g2041 ( 
.A(n_1635),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1635),
.B(n_1355),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1666),
.B(n_1359),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1666),
.B(n_1372),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1636),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1628),
.Y(n_2046)
);

AND2x6_ASAP7_75t_L g2047 ( 
.A(n_1626),
.B(n_1007),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1658),
.Y(n_2048)
);

AOI22x1_ASAP7_75t_SL g2049 ( 
.A1(n_1704),
.A2(n_1199),
.B1(n_1203),
.B2(n_1179),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1628),
.Y(n_2050)
);

CKINVDCx11_ASAP7_75t_R g2051 ( 
.A(n_1709),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1628),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1661),
.A2(n_1038),
.B1(n_1039),
.B2(n_1034),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1628),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1699),
.B(n_1114),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1628),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1628),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1658),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1659),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1628),
.Y(n_2060)
);

OAI21x1_ASAP7_75t_L g2061 ( 
.A1(n_1599),
.A2(n_1384),
.B(n_1383),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1628),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1661),
.A2(n_1052),
.B1(n_1057),
.B2(n_1044),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1659),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1628),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1628),
.Y(n_2066)
);

OA21x2_ASAP7_75t_L g2067 ( 
.A1(n_1599),
.A2(n_1423),
.B(n_1401),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_R g2068 ( 
.A(n_1887),
.B(n_1008),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_1780),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_R g2070 ( 
.A(n_1954),
.B(n_2006),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1804),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1858),
.B(n_1045),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1873),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1814),
.B(n_1009),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_R g2075 ( 
.A(n_1974),
.B(n_1988),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_2002),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1839),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1839),
.Y(n_2078)
);

CKINVDCx20_ASAP7_75t_R g2079 ( 
.A(n_1931),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1898),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1932),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1796),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1901),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1872),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_R g2085 ( 
.A(n_2026),
.B(n_1014),
.Y(n_2085)
);

NAND2x1_ASAP7_75t_L g2086 ( 
.A(n_1779),
.B(n_932),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1795),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1834),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_R g2089 ( 
.A(n_1963),
.B(n_1015),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_2051),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1850),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1815),
.B(n_1021),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1903),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1850),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1908),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1930),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1930),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1770),
.Y(n_2098)
);

NOR2xp67_ASAP7_75t_L g2099 ( 
.A(n_1842),
.B(n_1025),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_1818),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1852),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1935),
.B(n_1080),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1771),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1825),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1949),
.Y(n_2105)
);

CKINVDCx20_ASAP7_75t_R g2106 ( 
.A(n_1927),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1990),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_2009),
.Y(n_2108)
);

CKINVDCx20_ASAP7_75t_R g2109 ( 
.A(n_1806),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1912),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_R g2111 ( 
.A(n_1794),
.B(n_1027),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1893),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1917),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1832),
.Y(n_2114)
);

CKINVDCx16_ASAP7_75t_R g2115 ( 
.A(n_1829),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_2041),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_2031),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_2032),
.Y(n_2118)
);

BUFx10_ASAP7_75t_L g2119 ( 
.A(n_1781),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1876),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1859),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_1780),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1861),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1808),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1962),
.Y(n_2125)
);

NAND2xp33_ASAP7_75t_SL g2126 ( 
.A(n_1791),
.B(n_1218),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1862),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1819),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1773),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1843),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1843),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_2010),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1950),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1947),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_2039),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_1928),
.Y(n_2136)
);

INVxp67_ASAP7_75t_L g2137 ( 
.A(n_1907),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_R g2138 ( 
.A(n_1948),
.B(n_1032),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1879),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1914),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1881),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1884),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_R g2143 ( 
.A(n_1913),
.B(n_1059),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1914),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1885),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1970),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1983),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_2017),
.Y(n_2148)
);

CKINVDCx20_ASAP7_75t_R g2149 ( 
.A(n_1774),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_2045),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_R g2151 ( 
.A(n_1883),
.B(n_1041),
.Y(n_2151)
);

CKINVDCx20_ASAP7_75t_R g2152 ( 
.A(n_1811),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1886),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1775),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1777),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_1830),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1956),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1960),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_R g2159 ( 
.A(n_1782),
.B(n_1051),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1785),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_R g2161 ( 
.A(n_1783),
.B(n_1064),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1824),
.B(n_1066),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1976),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1984),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1799),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1920),
.B(n_905),
.Y(n_2166)
);

CKINVDCx20_ASAP7_75t_R g2167 ( 
.A(n_2016),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1890),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1979),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1821),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_1816),
.A2(n_1067),
.B1(n_1242),
.B2(n_1173),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1895),
.Y(n_2172)
);

CKINVDCx20_ASAP7_75t_R g2173 ( 
.A(n_2048),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1849),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_2058),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1895),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1900),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1900),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1866),
.B(n_947),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1909),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1909),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1856),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1867),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1891),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1981),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1985),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1993),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1865),
.B(n_1071),
.Y(n_2188)
);

CKINVDCx20_ASAP7_75t_R g2189 ( 
.A(n_2012),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_2013),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_2042),
.Y(n_2191)
);

CKINVDCx20_ASAP7_75t_R g2192 ( 
.A(n_1915),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_1786),
.A2(n_1349),
.B1(n_1398),
.B2(n_1303),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1940),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1994),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1790),
.B(n_1116),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1971),
.B(n_1074),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1870),
.B(n_1127),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1929),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_R g2200 ( 
.A(n_1778),
.B(n_1083),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_2049),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1789),
.Y(n_2202)
);

CKINVDCx20_ASAP7_75t_R g2203 ( 
.A(n_1997),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1937),
.Y(n_2204)
);

CKINVDCx16_ASAP7_75t_R g2205 ( 
.A(n_1798),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1944),
.Y(n_2206)
);

INVxp33_ASAP7_75t_L g2207 ( 
.A(n_1943),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_1789),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1916),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1951),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1967),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1916),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1998),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1926),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1986),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1987),
.Y(n_2216)
);

INVx1_ASAP7_75t_SL g2217 ( 
.A(n_1910),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_2028),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_2053),
.Y(n_2219)
);

AND2x6_ASAP7_75t_L g2220 ( 
.A(n_1788),
.B(n_1100),
.Y(n_2220)
);

BUFx10_ASAP7_75t_L g2221 ( 
.A(n_1889),
.Y(n_2221)
);

BUFx10_ASAP7_75t_L g2222 ( 
.A(n_1933),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_1802),
.Y(n_2223)
);

CKINVDCx5p33_ASAP7_75t_R g2224 ( 
.A(n_2063),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_1941),
.B(n_1854),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_1827),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1926),
.Y(n_2227)
);

CKINVDCx16_ASAP7_75t_R g2228 ( 
.A(n_1946),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1868),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1857),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_1869),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1905),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_1899),
.Y(n_2233)
);

CKINVDCx20_ASAP7_75t_R g2234 ( 
.A(n_2020),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1896),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1918),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1996),
.Y(n_2237)
);

NOR2xp67_ASAP7_75t_L g2238 ( 
.A(n_1904),
.B(n_1911),
.Y(n_2238)
);

CKINVDCx20_ASAP7_75t_R g2239 ( 
.A(n_2027),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_SL g2240 ( 
.A(n_1945),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_2029),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_2037),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_2043),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_2044),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1923),
.Y(n_2245)
);

CKINVDCx20_ASAP7_75t_R g2246 ( 
.A(n_2030),
.Y(n_2246)
);

CKINVDCx20_ASAP7_75t_R g2247 ( 
.A(n_2038),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2055),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1784),
.Y(n_2249)
);

AOI21x1_ASAP7_75t_L g2250 ( 
.A1(n_1863),
.A2(n_1440),
.B(n_1428),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1925),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2008),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_1860),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2014),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_1945),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_2015),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_2015),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1871),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_2047),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_2047),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1864),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1874),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_1864),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1875),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1875),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2019),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1878),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1882),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1880),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_1880),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2022),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2023),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1921),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_1922),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1888),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1924),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_2034),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1892),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_1902),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_1877),
.A2(n_1429),
.B1(n_1518),
.B2(n_1400),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_2046),
.Y(n_2281)
);

AOI21x1_ASAP7_75t_L g2282 ( 
.A1(n_1897),
.A2(n_1459),
.B(n_1450),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1833),
.B(n_954),
.Y(n_2283)
);

CKINVDCx20_ASAP7_75t_R g2284 ( 
.A(n_1906),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1831),
.Y(n_2285)
);

AOI21x1_ASAP7_75t_L g2286 ( 
.A1(n_1894),
.A2(n_1478),
.B(n_1464),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1797),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1919),
.Y(n_2288)
);

CKINVDCx20_ASAP7_75t_R g2289 ( 
.A(n_1835),
.Y(n_2289)
);

CKINVDCx20_ASAP7_75t_R g2290 ( 
.A(n_1851),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2056),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1812),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_1812),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2057),
.B(n_1088),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1800),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1817),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_R g2297 ( 
.A(n_1837),
.B(n_1103),
.Y(n_2297)
);

CKINVDCx16_ASAP7_75t_R g2298 ( 
.A(n_1841),
.Y(n_2298)
);

CKINVDCx20_ASAP7_75t_R g2299 ( 
.A(n_1952),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1803),
.Y(n_2300)
);

CKINVDCx20_ASAP7_75t_R g2301 ( 
.A(n_1959),
.Y(n_2301)
);

CKINVDCx20_ASAP7_75t_R g2302 ( 
.A(n_2036),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1817),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_1938),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1938),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_R g2306 ( 
.A(n_1807),
.B(n_1110),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_1953),
.Y(n_2307)
);

BUFx8_ASAP7_75t_L g2308 ( 
.A(n_1809),
.Y(n_2308)
);

CKINVDCx20_ASAP7_75t_R g2309 ( 
.A(n_2067),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2060),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_1953),
.Y(n_2311)
);

BUFx10_ASAP7_75t_L g2312 ( 
.A(n_1813),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1957),
.Y(n_2313)
);

CKINVDCx20_ASAP7_75t_R g2314 ( 
.A(n_1820),
.Y(n_2314)
);

OR2x6_ASAP7_75t_L g2315 ( 
.A(n_2025),
.B(n_1164),
.Y(n_2315)
);

BUFx10_ASAP7_75t_L g2316 ( 
.A(n_1822),
.Y(n_2316)
);

CKINVDCx20_ASAP7_75t_R g2317 ( 
.A(n_1823),
.Y(n_2317)
);

AOI22xp33_ASAP7_75t_SL g2318 ( 
.A1(n_1838),
.A2(n_1250),
.B1(n_1258),
.B2(n_1232),
.Y(n_2318)
);

CKINVDCx20_ASAP7_75t_R g2319 ( 
.A(n_1840),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_1964),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_1964),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_1975),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1844),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1975),
.B(n_1343),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1847),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_1980),
.Y(n_2326)
);

CKINVDCx5p33_ASAP7_75t_R g2327 ( 
.A(n_1980),
.Y(n_2327)
);

INVx8_ASAP7_75t_L g2328 ( 
.A(n_1991),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1853),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1991),
.Y(n_2330)
);

INVx4_ASAP7_75t_L g2331 ( 
.A(n_2261),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_2109),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2121),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2123),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2217),
.B(n_954),
.Y(n_2335)
);

OR2x2_ASAP7_75t_SL g2336 ( 
.A(n_2115),
.B(n_876),
.Y(n_2336)
);

BUFx3_ASAP7_75t_L g2337 ( 
.A(n_2117),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2127),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2185),
.B(n_1855),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_2084),
.Y(n_2340)
);

NAND3xp33_ASAP7_75t_L g2341 ( 
.A(n_2102),
.B(n_1061),
.C(n_1060),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2202),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2179),
.B(n_954),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_2207),
.B(n_2175),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2186),
.B(n_1129),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2187),
.A2(n_1483),
.B1(n_1494),
.B2(n_1481),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2139),
.Y(n_2347)
);

INVx5_ASAP7_75t_L g2348 ( 
.A(n_2221),
.Y(n_2348)
);

INVx3_ASAP7_75t_L g2349 ( 
.A(n_2156),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2114),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2141),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_2289),
.A2(n_1514),
.B1(n_1551),
.B2(n_1521),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2103),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_2118),
.Y(n_2354)
);

BUFx10_ASAP7_75t_L g2355 ( 
.A(n_2082),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2129),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2202),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2142),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_2075),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2202),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2133),
.Y(n_2361)
);

NOR2x1p5_ASAP7_75t_L g2362 ( 
.A(n_2124),
.B(n_1072),
.Y(n_2362)
);

INVx5_ASAP7_75t_L g2363 ( 
.A(n_2221),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2223),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2096),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2157),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2163),
.B(n_1075),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2190),
.B(n_1131),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_2164),
.B(n_1076),
.Y(n_2369)
);

NAND3xp33_ASAP7_75t_L g2370 ( 
.A(n_2072),
.B(n_2225),
.C(n_2137),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2080),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2158),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2083),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_2191),
.B(n_1078),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2279),
.B(n_2288),
.Y(n_2375)
);

INVxp67_ASAP7_75t_SL g2376 ( 
.A(n_2253),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2169),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_2223),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2222),
.B(n_2283),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2150),
.B(n_1772),
.Y(n_2380)
);

BUFx3_ASAP7_75t_L g2381 ( 
.A(n_2097),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2093),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_2149),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2165),
.B(n_1081),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2143),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2095),
.Y(n_2386)
);

AND2x6_ASAP7_75t_L g2387 ( 
.A(n_2198),
.B(n_2196),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2170),
.B(n_1082),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2110),
.Y(n_2389)
);

INVx2_ASAP7_75t_SL g2390 ( 
.A(n_2222),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2113),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2195),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2172),
.B(n_1776),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2174),
.B(n_2182),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2183),
.B(n_2184),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_2176),
.B(n_1787),
.Y(n_2396)
);

BUFx10_ASAP7_75t_L g2397 ( 
.A(n_2088),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2213),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2177),
.B(n_1792),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2154),
.B(n_1801),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2263),
.B(n_965),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2264),
.Y(n_2402)
);

BUFx6f_ASAP7_75t_L g2403 ( 
.A(n_2328),
.Y(n_2403)
);

INVx1_ASAP7_75t_SL g2404 ( 
.A(n_2152),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2265),
.B(n_965),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2155),
.B(n_1084),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2287),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2290),
.A2(n_1554),
.B1(n_1572),
.B2(n_1567),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2295),
.Y(n_2409)
);

INVx4_ASAP7_75t_L g2410 ( 
.A(n_2269),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2300),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2252),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2323),
.Y(n_2413)
);

BUFx4f_ASAP7_75t_L g2414 ( 
.A(n_2255),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2128),
.B(n_1086),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2254),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_R g2417 ( 
.A(n_2071),
.B(n_1133),
.Y(n_2417)
);

AND2x6_ASAP7_75t_L g2418 ( 
.A(n_2166),
.B(n_1100),
.Y(n_2418)
);

INVx3_ASAP7_75t_L g2419 ( 
.A(n_2270),
.Y(n_2419)
);

AND2x6_ASAP7_75t_L g2420 ( 
.A(n_2166),
.B(n_1100),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2328),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_2330),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2178),
.B(n_1934),
.Y(n_2423)
);

OR2x6_ASAP7_75t_L g2424 ( 
.A(n_2315),
.B(n_1220),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2258),
.B(n_1805),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2262),
.B(n_1810),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2229),
.B(n_1089),
.Y(n_2427)
);

INVx1_ASAP7_75t_SL g2428 ( 
.A(n_2167),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2205),
.B(n_965),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2325),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2228),
.B(n_1079),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2329),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2266),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2271),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2173),
.Y(n_2435)
);

BUFx10_ASAP7_75t_L g2436 ( 
.A(n_2090),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2272),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2248),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_L g2439 ( 
.A(n_2284),
.B(n_1090),
.Y(n_2439)
);

AND2x2_ASAP7_75t_SL g2440 ( 
.A(n_2298),
.B(n_876),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2299),
.A2(n_2301),
.B1(n_2309),
.B2(n_2302),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2267),
.B(n_1826),
.Y(n_2442)
);

INVx1_ASAP7_75t_SL g2443 ( 
.A(n_2189),
.Y(n_2443)
);

INVx1_ASAP7_75t_SL g2444 ( 
.A(n_2314),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2193),
.B(n_1482),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2188),
.B(n_1091),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2281),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2292),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2291),
.Y(n_2449)
);

HB1xp67_ASAP7_75t_L g2450 ( 
.A(n_2235),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2273),
.B(n_1138),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2310),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2274),
.B(n_1140),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2276),
.B(n_1079),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2268),
.B(n_1828),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2230),
.B(n_1094),
.Y(n_2456)
);

NAND3xp33_ASAP7_75t_L g2457 ( 
.A(n_2280),
.B(n_1104),
.C(n_1102),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2226),
.A2(n_1141),
.B1(n_1154),
.B2(n_1153),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2232),
.Y(n_2459)
);

OAI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2197),
.A2(n_1598),
.B1(n_1575),
.B2(n_1167),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2275),
.Y(n_2461)
);

BUFx3_ASAP7_75t_L g2462 ( 
.A(n_2293),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2119),
.B(n_1079),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2278),
.Y(n_2464)
);

CKINVDCx8_ASAP7_75t_R g2465 ( 
.A(n_2073),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2159),
.B(n_1845),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2317),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2161),
.B(n_1848),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2236),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2119),
.B(n_1099),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2180),
.B(n_1936),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2069),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_2076),
.Y(n_2473)
);

XOR2xp5_ASAP7_75t_L g2474 ( 
.A(n_2079),
.B(n_2106),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2245),
.Y(n_2475)
);

INVx1_ASAP7_75t_SL g2476 ( 
.A(n_2319),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2251),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2277),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2328),
.Y(n_2479)
);

AND2x4_ASAP7_75t_L g2480 ( 
.A(n_2181),
.B(n_1939),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2285),
.Y(n_2481)
);

AND2x2_ASAP7_75t_SL g2482 ( 
.A(n_2087),
.B(n_880),
.Y(n_2482)
);

OR2x2_ASAP7_75t_L g2483 ( 
.A(n_2126),
.B(n_1574),
.Y(n_2483)
);

AND2x6_ASAP7_75t_L g2484 ( 
.A(n_2074),
.B(n_1100),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2209),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2220),
.B(n_1942),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2077),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_2296),
.Y(n_2488)
);

INVx6_ASAP7_75t_L g2489 ( 
.A(n_2308),
.Y(n_2489)
);

AND2x6_ASAP7_75t_L g2490 ( 
.A(n_2092),
.B(n_1139),
.Y(n_2490)
);

BUFx4f_ASAP7_75t_L g2491 ( 
.A(n_2315),
.Y(n_2491)
);

OR2x2_ASAP7_75t_L g2492 ( 
.A(n_2162),
.B(n_1106),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2212),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2112),
.B(n_1159),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2220),
.B(n_1955),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2214),
.B(n_2227),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2122),
.Y(n_2497)
);

OR2x2_ASAP7_75t_L g2498 ( 
.A(n_2100),
.B(n_1107),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2078),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2146),
.B(n_2147),
.Y(n_2500)
);

AOI22xp33_ASAP7_75t_L g2501 ( 
.A1(n_2086),
.A2(n_982),
.B1(n_1836),
.B2(n_1793),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2122),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2303),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2148),
.B(n_1099),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2208),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2091),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2304),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2094),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2101),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2104),
.Y(n_2510)
);

INVx5_ASAP7_75t_L g2511 ( 
.A(n_2315),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2145),
.Y(n_2512)
);

INVx2_ASAP7_75t_SL g2513 ( 
.A(n_2312),
.Y(n_2513)
);

XNOR2xp5_ASAP7_75t_L g2514 ( 
.A(n_2081),
.B(n_1268),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2231),
.B(n_1108),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2134),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2220),
.B(n_1958),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2256),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2116),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2204),
.B(n_1111),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2294),
.B(n_1961),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2153),
.Y(n_2522)
);

AND2x4_ASAP7_75t_L g2523 ( 
.A(n_2238),
.B(n_1965),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2168),
.B(n_1968),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2151),
.B(n_1169),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2312),
.Y(n_2526)
);

INVx4_ASAP7_75t_L g2527 ( 
.A(n_2305),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2307),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2282),
.Y(n_2529)
);

AOI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2206),
.A2(n_1175),
.B1(n_1178),
.B2(n_1177),
.Y(n_2530)
);

BUFx4_ASAP7_75t_L g2531 ( 
.A(n_2125),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2311),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2316),
.Y(n_2533)
);

NAND2xp33_ASAP7_75t_L g2534 ( 
.A(n_2194),
.B(n_982),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_2237),
.B(n_1181),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2316),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2250),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2241),
.B(n_1186),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2257),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2286),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_2313),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2403),
.B(n_2320),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2403),
.B(n_2321),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2333),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2353),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2334),
.Y(n_2546)
);

INVx2_ASAP7_75t_SL g2547 ( 
.A(n_2344),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2356),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2338),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2361),
.Y(n_2550)
);

BUFx8_ASAP7_75t_L g2551 ( 
.A(n_2383),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2446),
.B(n_2200),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2352),
.A2(n_2408),
.B1(n_2441),
.B2(n_2395),
.Y(n_2553)
);

NAND2x1p5_ASAP7_75t_L g2554 ( 
.A(n_2421),
.B(n_2000),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2394),
.B(n_2210),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2366),
.Y(n_2556)
);

OAI221xp5_ASAP7_75t_L g2557 ( 
.A1(n_2346),
.A2(n_2318),
.B1(n_2211),
.B2(n_2218),
.C(n_2216),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2350),
.Y(n_2558)
);

BUFx2_ASAP7_75t_L g2559 ( 
.A(n_2340),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_L g2560 ( 
.A1(n_2534),
.A2(n_2219),
.B1(n_2224),
.B2(n_2215),
.Y(n_2560)
);

OR2x6_ASAP7_75t_SL g2561 ( 
.A(n_2519),
.B(n_2160),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2347),
.Y(n_2562)
);

INVxp67_ASAP7_75t_L g2563 ( 
.A(n_2335),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2387),
.B(n_2242),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2351),
.Y(n_2565)
);

NAND2x1p5_ASAP7_75t_L g2566 ( 
.A(n_2421),
.B(n_2001),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2387),
.B(n_2243),
.Y(n_2567)
);

AOI22xp33_ASAP7_75t_L g2568 ( 
.A1(n_2358),
.A2(n_2171),
.B1(n_2233),
.B2(n_2249),
.Y(n_2568)
);

INVx4_ASAP7_75t_L g2569 ( 
.A(n_2479),
.Y(n_2569)
);

OAI221xp5_ASAP7_75t_L g2570 ( 
.A1(n_2427),
.A2(n_2341),
.B1(n_2370),
.B2(n_2483),
.C(n_2458),
.Y(n_2570)
);

INVxp67_ASAP7_75t_L g2571 ( 
.A(n_2343),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_2479),
.B(n_2322),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2387),
.B(n_2244),
.Y(n_2573)
);

AND2x6_ASAP7_75t_L g2574 ( 
.A(n_2379),
.B(n_1139),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2371),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2373),
.Y(n_2576)
);

AO22x2_ASAP7_75t_L g2577 ( 
.A1(n_2445),
.A2(n_2375),
.B1(n_2476),
.B2(n_2444),
.Y(n_2577)
);

CKINVDCx16_ASAP7_75t_R g2578 ( 
.A(n_2365),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2374),
.B(n_2138),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2372),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2377),
.Y(n_2581)
);

OAI21xp33_ASAP7_75t_L g2582 ( 
.A1(n_2367),
.A2(n_2260),
.B(n_2259),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2482),
.B(n_2132),
.Y(n_2583)
);

AND2x2_ASAP7_75t_SL g2584 ( 
.A(n_2467),
.B(n_2240),
.Y(n_2584)
);

BUFx8_ASAP7_75t_L g2585 ( 
.A(n_2488),
.Y(n_2585)
);

AOI211xp5_ASAP7_75t_L g2586 ( 
.A1(n_2456),
.A2(n_2089),
.B(n_2324),
.C(n_2085),
.Y(n_2586)
);

CKINVDCx20_ASAP7_75t_R g2587 ( 
.A(n_2465),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2384),
.B(n_2388),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2382),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2369),
.B(n_2385),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2386),
.Y(n_2591)
);

AND2x4_ASAP7_75t_L g2592 ( 
.A(n_2381),
.B(n_2326),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2438),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2392),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2389),
.Y(n_2595)
);

AO22x2_ASAP7_75t_L g2596 ( 
.A1(n_2404),
.A2(n_928),
.B1(n_1029),
.B2(n_896),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2415),
.A2(n_2203),
.B1(n_2239),
.B2(n_2234),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2391),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2407),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2336),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2409),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_SL g2602 ( 
.A1(n_2515),
.A2(n_2247),
.B1(n_2246),
.B2(n_2136),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2411),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2413),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2400),
.B(n_2099),
.Y(n_2605)
);

INVxp67_ASAP7_75t_L g2606 ( 
.A(n_2401),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2520),
.A2(n_2070),
.B1(n_2135),
.B2(n_2192),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2398),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2430),
.A2(n_982),
.B1(n_1282),
.B2(n_1139),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2412),
.Y(n_2610)
);

NAND2x1_ASAP7_75t_L g2611 ( 
.A(n_2537),
.B(n_1969),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2432),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2433),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2449),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2492),
.A2(n_1310),
.B1(n_1317),
.B2(n_1274),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2425),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2426),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2339),
.B(n_2297),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2406),
.B(n_2306),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2443),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2442),
.Y(n_2621)
);

NAND2x1p5_ASAP7_75t_L g2622 ( 
.A(n_2402),
.B(n_2419),
.Y(n_2622)
);

NAND2x1p5_ASAP7_75t_L g2623 ( 
.A(n_2331),
.B(n_2410),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2521),
.B(n_2327),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_2405),
.Y(n_2625)
);

NAND2x1p5_ASAP7_75t_L g2626 ( 
.A(n_2507),
.B(n_2001),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2455),
.Y(n_2627)
);

AND2x6_ASAP7_75t_L g2628 ( 
.A(n_2540),
.B(n_1139),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2459),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2469),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2439),
.B(n_2130),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2473),
.Y(n_2632)
);

NAND2x1p5_ASAP7_75t_L g2633 ( 
.A(n_2488),
.B(n_2011),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2440),
.B(n_2068),
.Y(n_2634)
);

NAND3x1_ASAP7_75t_L g2635 ( 
.A(n_2530),
.B(n_2201),
.C(n_2199),
.Y(n_2635)
);

INVxp67_ASAP7_75t_L g2636 ( 
.A(n_2454),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2416),
.Y(n_2637)
);

NAND2x1p5_ASAP7_75t_L g2638 ( 
.A(n_2503),
.B(n_2011),
.Y(n_2638)
);

INVxp67_ASAP7_75t_L g2639 ( 
.A(n_2504),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2434),
.Y(n_2640)
);

OAI221xp5_ASAP7_75t_L g2641 ( 
.A1(n_2457),
.A2(n_914),
.B1(n_917),
.B2(n_913),
.C(n_912),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2437),
.Y(n_2642)
);

BUFx8_ASAP7_75t_L g2643 ( 
.A(n_2503),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2448),
.B(n_2120),
.Y(n_2644)
);

BUFx8_ASAP7_75t_L g2645 ( 
.A(n_2528),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2447),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2452),
.B(n_1972),
.Y(n_2647)
);

INVxp67_ASAP7_75t_L g2648 ( 
.A(n_2498),
.Y(n_2648)
);

NAND2xp33_ASAP7_75t_L g2649 ( 
.A(n_2484),
.B(n_2131),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2462),
.B(n_2098),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2463),
.B(n_2111),
.Y(n_2651)
);

BUFx6f_ASAP7_75t_L g2652 ( 
.A(n_2342),
.Y(n_2652)
);

AOI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2460),
.A2(n_1197),
.B1(n_1216),
.B2(n_1207),
.Y(n_2653)
);

BUFx3_ASAP7_75t_L g2654 ( 
.A(n_2528),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2345),
.B(n_1322),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2524),
.Y(n_2656)
);

AO22x2_ASAP7_75t_L g2657 ( 
.A1(n_2428),
.A2(n_1037),
.B1(n_1058),
.B2(n_1029),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2368),
.B(n_1348),
.Y(n_2658)
);

CKINVDCx20_ASAP7_75t_R g2659 ( 
.A(n_2359),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_2417),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2461),
.Y(n_2661)
);

BUFx8_ASAP7_75t_L g2662 ( 
.A(n_2532),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2464),
.Y(n_2663)
);

BUFx8_ASAP7_75t_L g2664 ( 
.A(n_2532),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2470),
.B(n_1421),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2475),
.Y(n_2666)
);

HB1xp67_ASAP7_75t_L g2667 ( 
.A(n_2541),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2477),
.A2(n_1217),
.B1(n_1225),
.B2(n_1223),
.Y(n_2668)
);

BUFx4f_ASAP7_75t_L g2669 ( 
.A(n_2541),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2481),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2487),
.Y(n_2671)
);

INVxp67_ASAP7_75t_L g2672 ( 
.A(n_2429),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2435),
.B(n_2105),
.Y(n_2673)
);

AO22x2_ASAP7_75t_L g2674 ( 
.A1(n_2474),
.A2(n_1058),
.B1(n_1124),
.B2(n_1037),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2513),
.B(n_1457),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2466),
.B(n_1973),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2511),
.B(n_2107),
.Y(n_2677)
);

CKINVDCx20_ASAP7_75t_R g2678 ( 
.A(n_2332),
.Y(n_2678)
);

BUFx6f_ASAP7_75t_SL g2679 ( 
.A(n_2355),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2500),
.B(n_2376),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2485),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2493),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2484),
.A2(n_982),
.B1(n_1282),
.B2(n_1474),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2468),
.B(n_2478),
.Y(n_2684)
);

AO22x2_ASAP7_75t_L g2685 ( 
.A1(n_2526),
.A2(n_2536),
.B1(n_2533),
.B2(n_2431),
.Y(n_2685)
);

A2O1A1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2491),
.A2(n_1846),
.B(n_1995),
.C(n_1966),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2499),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2522),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2342),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2393),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2484),
.B(n_1977),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2396),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2490),
.B(n_1978),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2399),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2423),
.Y(n_2695)
);

INVxp67_ASAP7_75t_L g2696 ( 
.A(n_2450),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2471),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2510),
.A2(n_1492),
.B1(n_1499),
.B2(n_1476),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2349),
.B(n_2108),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2480),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2490),
.B(n_1982),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2506),
.Y(n_2702)
);

BUFx2_ASAP7_75t_L g2703 ( 
.A(n_2337),
.Y(n_2703)
);

BUFx2_ASAP7_75t_L g2704 ( 
.A(n_2354),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2516),
.B(n_1522),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2490),
.A2(n_982),
.B1(n_1282),
.B2(n_1525),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2508),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2512),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2529),
.A2(n_982),
.B1(n_1282),
.B2(n_1542),
.Y(n_2709)
);

CKINVDCx20_ASAP7_75t_R g2710 ( 
.A(n_2397),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2509),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2497),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2422),
.Y(n_2713)
);

NAND3xp33_ASAP7_75t_L g2714 ( 
.A(n_2451),
.B(n_2308),
.C(n_2144),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2502),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2545),
.Y(n_2716)
);

BUFx2_ASAP7_75t_SL g2717 ( 
.A(n_2654),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_R g2718 ( 
.A(n_2569),
.B(n_2489),
.Y(n_2718)
);

AOI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2605),
.A2(n_2525),
.B(n_2501),
.Y(n_2719)
);

OAI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2709),
.A2(n_2040),
.B(n_2005),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2588),
.B(n_2494),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2590),
.B(n_2453),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2544),
.Y(n_2723)
);

AO21x1_ASAP7_75t_L g2724 ( 
.A1(n_2553),
.A2(n_2495),
.B(n_2486),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_2555),
.B(n_2579),
.Y(n_2725)
);

BUFx2_ASAP7_75t_L g2726 ( 
.A(n_2559),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2558),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2656),
.B(n_2380),
.Y(n_2728)
);

OAI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2560),
.A2(n_2414),
.B1(n_2390),
.B2(n_2518),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2616),
.B(n_2523),
.Y(n_2730)
);

A2O1A1Ixp33_ASAP7_75t_L g2731 ( 
.A1(n_2655),
.A2(n_2505),
.B(n_2496),
.C(n_2535),
.Y(n_2731)
);

BUFx12f_ASAP7_75t_L g2732 ( 
.A(n_2585),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2618),
.A2(n_2517),
.B(n_2538),
.Y(n_2733)
);

OAI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2617),
.A2(n_2061),
.B(n_2472),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2570),
.A2(n_2539),
.B1(n_2420),
.B2(n_2418),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2546),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2549),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2552),
.A2(n_2684),
.B(n_2621),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_SL g2739 ( 
.A(n_2619),
.B(n_2527),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2627),
.A2(n_2364),
.B(n_2360),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2624),
.B(n_2418),
.Y(n_2741)
);

AND2x2_ASAP7_75t_SL g2742 ( 
.A(n_2669),
.B(n_2364),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2548),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_2680),
.B(n_2348),
.Y(n_2744)
);

AOI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2676),
.A2(n_2378),
.B(n_2357),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2665),
.B(n_2348),
.Y(n_2746)
);

O2A1O1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2571),
.A2(n_2424),
.B(n_922),
.C(n_923),
.Y(n_2747)
);

O2A1O1Ixp33_ASAP7_75t_SL g2748 ( 
.A1(n_2686),
.A2(n_930),
.B(n_934),
.C(n_919),
.Y(n_2748)
);

NOR2x1_ASAP7_75t_L g2749 ( 
.A(n_2587),
.B(n_2362),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2607),
.B(n_2363),
.Y(n_2750)
);

INVxp67_ASAP7_75t_L g2751 ( 
.A(n_2593),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_2563),
.B(n_2436),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2611),
.A2(n_2018),
.B(n_2033),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2562),
.B(n_2420),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2565),
.Y(n_2755)
);

AO31x2_ASAP7_75t_L g2756 ( 
.A1(n_2691),
.A2(n_1204),
.A3(n_1253),
.B(n_1170),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2651),
.B(n_2514),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2550),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_SL g2759 ( 
.A(n_2632),
.B(n_2660),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2556),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2575),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2658),
.A2(n_2420),
.B1(n_1233),
.B2(n_1240),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2576),
.B(n_1989),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2648),
.B(n_1099),
.Y(n_2764)
);

O2A1O1Ixp33_ASAP7_75t_L g2765 ( 
.A1(n_2634),
.A2(n_948),
.B(n_951),
.C(n_941),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2589),
.B(n_1992),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2659),
.Y(n_2767)
);

AO21x1_ASAP7_75t_L g2768 ( 
.A1(n_2693),
.A2(n_971),
.B(n_957),
.Y(n_2768)
);

OAI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2557),
.A2(n_1569),
.B1(n_1570),
.B2(n_1561),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2591),
.B(n_2595),
.Y(n_2770)
);

BUFx2_ASAP7_75t_L g2771 ( 
.A(n_2643),
.Y(n_2771)
);

A2O1A1Ixp33_ASAP7_75t_L g2772 ( 
.A1(n_2598),
.A2(n_2601),
.B(n_2603),
.C(n_2599),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2615),
.B(n_2140),
.Y(n_2773)
);

INVx3_ASAP7_75t_SL g2774 ( 
.A(n_2578),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2604),
.B(n_1999),
.Y(n_2775)
);

O2A1O1Ixp33_ASAP7_75t_L g2776 ( 
.A1(n_2641),
.A2(n_980),
.B(n_986),
.C(n_979),
.Y(n_2776)
);

OAI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2612),
.A2(n_2066),
.B(n_2065),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2568),
.A2(n_1248),
.B1(n_1249),
.B2(n_1230),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2620),
.B(n_2003),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2580),
.A2(n_2064),
.B(n_2059),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2652),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2629),
.B(n_2004),
.Y(n_2782)
);

AOI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2581),
.A2(n_2064),
.B(n_1262),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2630),
.A2(n_996),
.B(n_1000),
.C(n_989),
.Y(n_2784)
);

AOI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2712),
.A2(n_2021),
.B(n_2007),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2594),
.Y(n_2786)
);

A2O1A1Ixp33_ASAP7_75t_L g2787 ( 
.A1(n_2670),
.A2(n_1005),
.B(n_1006),
.C(n_1003),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2661),
.B(n_2024),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2663),
.B(n_2035),
.Y(n_2789)
);

O2A1O1Ixp33_ASAP7_75t_L g2790 ( 
.A1(n_2606),
.A2(n_1013),
.B(n_1016),
.C(n_1010),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2608),
.Y(n_2791)
);

INVx11_ASAP7_75t_L g2792 ( 
.A(n_2645),
.Y(n_2792)
);

NAND3xp33_ASAP7_75t_L g2793 ( 
.A(n_2705),
.B(n_1118),
.C(n_1117),
.Y(n_2793)
);

OR2x6_ASAP7_75t_L g2794 ( 
.A(n_2592),
.B(n_2531),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2666),
.B(n_2613),
.Y(n_2795)
);

BUFx6f_ASAP7_75t_L g2796 ( 
.A(n_2652),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2610),
.A2(n_1286),
.B(n_1280),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2636),
.A2(n_1296),
.B1(n_1299),
.B2(n_1288),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2547),
.B(n_1119),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_SL g2800 ( 
.A(n_2644),
.B(n_1343),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2681),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2678),
.Y(n_2802)
);

AO21x1_ASAP7_75t_L g2803 ( 
.A1(n_2701),
.A2(n_1023),
.B(n_1018),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2614),
.B(n_2050),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_2667),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2642),
.Y(n_2806)
);

A2O1A1Ixp33_ASAP7_75t_L g2807 ( 
.A1(n_2625),
.A2(n_1035),
.B(n_1036),
.C(n_1026),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2682),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2637),
.B(n_2052),
.Y(n_2809)
);

AOI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2639),
.A2(n_1319),
.B1(n_1339),
.B2(n_1306),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2631),
.B(n_1121),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2672),
.B(n_1184),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2640),
.B(n_2054),
.Y(n_2813)
);

BUFx4f_ASAP7_75t_L g2814 ( 
.A(n_2542),
.Y(n_2814)
);

CKINVDCx16_ASAP7_75t_R g2815 ( 
.A(n_2679),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2688),
.Y(n_2816)
);

INVx2_ASAP7_75t_SL g2817 ( 
.A(n_2543),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2715),
.A2(n_2564),
.B1(n_2573),
.B2(n_2567),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2582),
.B(n_1123),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2600),
.B(n_1184),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2675),
.B(n_1125),
.Y(n_2821)
);

AOI21x1_ASAP7_75t_L g2822 ( 
.A1(n_2647),
.A2(n_2062),
.B(n_1047),
.Y(n_2822)
);

AOI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2646),
.A2(n_1368),
.B(n_1366),
.Y(n_2823)
);

OAI321xp33_ASAP7_75t_L g2824 ( 
.A1(n_2698),
.A2(n_2683),
.A3(n_2706),
.B1(n_2586),
.B2(n_2583),
.C(n_2597),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2572),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2708),
.B(n_1369),
.Y(n_2826)
);

OAI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2702),
.A2(n_1379),
.B1(n_1385),
.B2(n_1376),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2707),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2671),
.A2(n_1392),
.B(n_1391),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2687),
.A2(n_1396),
.B(n_1393),
.Y(n_2830)
);

INVx2_ASAP7_75t_SL g2831 ( 
.A(n_2662),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2602),
.B(n_1404),
.Y(n_2832)
);

OAI21x1_ASAP7_75t_L g2833 ( 
.A1(n_2711),
.A2(n_1271),
.B(n_1253),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2690),
.A2(n_1420),
.B(n_1410),
.Y(n_2834)
);

O2A1O1Ixp5_ASAP7_75t_L g2835 ( 
.A1(n_2713),
.A2(n_1275),
.B(n_1283),
.C(n_1271),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2697),
.A2(n_2694),
.B(n_2692),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2695),
.A2(n_2700),
.B(n_2649),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2689),
.A2(n_1448),
.B(n_1446),
.Y(n_2838)
);

AO21x1_ASAP7_75t_L g2839 ( 
.A1(n_2653),
.A2(n_1048),
.B(n_1046),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2574),
.B(n_1454),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2574),
.B(n_1463),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2554),
.Y(n_2842)
);

NOR2x1_ASAP7_75t_R g2843 ( 
.A(n_2732),
.B(n_2650),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2725),
.B(n_2722),
.Y(n_2844)
);

NOR3xp33_ASAP7_75t_SL g2845 ( 
.A(n_2769),
.B(n_2714),
.C(n_2677),
.Y(n_2845)
);

AOI221x1_ASAP7_75t_L g2846 ( 
.A1(n_2818),
.A2(n_2577),
.B1(n_2821),
.B2(n_2738),
.C(n_2811),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2723),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2736),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2719),
.A2(n_2622),
.B(n_2623),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2737),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2721),
.B(n_2584),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2742),
.B(n_2696),
.Y(n_2852)
);

CKINVDCx16_ASAP7_75t_R g2853 ( 
.A(n_2759),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2728),
.B(n_2577),
.Y(n_2854)
);

A2O1A1Ixp33_ASAP7_75t_L g2855 ( 
.A1(n_2824),
.A2(n_2668),
.B(n_2699),
.C(n_2609),
.Y(n_2855)
);

INVx2_ASAP7_75t_SL g2856 ( 
.A(n_2814),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2802),
.B(n_2703),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2755),
.Y(n_2858)
);

AND2x4_ASAP7_75t_L g2859 ( 
.A(n_2817),
.B(n_2704),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2746),
.B(n_2664),
.Y(n_2860)
);

AO21x1_ASAP7_75t_L g2861 ( 
.A1(n_2733),
.A2(n_2626),
.B(n_1055),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2730),
.B(n_2596),
.Y(n_2862)
);

AOI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_2720),
.A2(n_2685),
.B(n_2566),
.Y(n_2863)
);

OR2x2_ASAP7_75t_L g2864 ( 
.A(n_2726),
.B(n_2673),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2757),
.B(n_2674),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2773),
.A2(n_2710),
.B1(n_2635),
.B2(n_2685),
.Y(n_2866)
);

AOI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2734),
.A2(n_2638),
.B(n_2633),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2761),
.Y(n_2868)
);

BUFx2_ASAP7_75t_L g2869 ( 
.A(n_2727),
.Y(n_2869)
);

OAI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2770),
.A2(n_2657),
.B1(n_2561),
.B2(n_2674),
.Y(n_2870)
);

OR2x6_ASAP7_75t_SL g2871 ( 
.A(n_2767),
.B(n_1144),
.Y(n_2871)
);

A2O1A1Ixp33_ASAP7_75t_L g2872 ( 
.A1(n_2819),
.A2(n_1056),
.B(n_1062),
.C(n_1050),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2801),
.B(n_2628),
.Y(n_2873)
);

OAI21xp33_ASAP7_75t_L g2874 ( 
.A1(n_2800),
.A2(n_1148),
.B(n_1145),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2748),
.A2(n_2628),
.B(n_1498),
.Y(n_2875)
);

AOI22xp5_ASAP7_75t_L g2876 ( 
.A1(n_2750),
.A2(n_2551),
.B1(n_1501),
.B2(n_1511),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2808),
.B(n_2628),
.Y(n_2877)
);

OR2x6_ASAP7_75t_L g2878 ( 
.A(n_2717),
.B(n_1580),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2731),
.A2(n_1512),
.B(n_1491),
.Y(n_2879)
);

AOI21x1_ASAP7_75t_L g2880 ( 
.A1(n_2724),
.A2(n_1087),
.B(n_1085),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2741),
.A2(n_1536),
.B(n_1515),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2816),
.B(n_1562),
.Y(n_2882)
);

A2O1A1Ixp33_ASAP7_75t_L g2883 ( 
.A1(n_2793),
.A2(n_1105),
.B(n_1112),
.C(n_1098),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2751),
.B(n_1149),
.Y(n_2884)
);

O2A1O1Ixp33_ASAP7_75t_L g2885 ( 
.A1(n_2807),
.A2(n_1115),
.B(n_1120),
.C(n_1113),
.Y(n_2885)
);

NOR2xp33_ASAP7_75t_L g2886 ( 
.A(n_2832),
.B(n_1150),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2799),
.B(n_1151),
.Y(n_2887)
);

BUFx4f_ASAP7_75t_L g2888 ( 
.A(n_2774),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2828),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2825),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2729),
.B(n_1443),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2739),
.A2(n_1565),
.B(n_1563),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2764),
.B(n_1184),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2795),
.B(n_1564),
.Y(n_2894)
);

NAND2xp33_ASAP7_75t_L g2895 ( 
.A(n_2772),
.B(n_1152),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2744),
.B(n_1155),
.Y(n_2896)
);

OR2x2_ASAP7_75t_L g2897 ( 
.A(n_2805),
.B(n_1158),
.Y(n_2897)
);

A2O1A1Ixp33_ASAP7_75t_SL g2898 ( 
.A1(n_2735),
.A2(n_1128),
.B(n_1132),
.C(n_1126),
.Y(n_2898)
);

BUFx6f_ASAP7_75t_L g2899 ( 
.A(n_2781),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2716),
.Y(n_2900)
);

OAI21xp33_ASAP7_75t_L g2901 ( 
.A1(n_2820),
.A2(n_1162),
.B(n_1161),
.Y(n_2901)
);

BUFx8_ASAP7_75t_SL g2902 ( 
.A(n_2771),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_2779),
.B(n_1235),
.Y(n_2903)
);

NOR3xp33_ASAP7_75t_SL g2904 ( 
.A(n_2752),
.B(n_1176),
.C(n_1174),
.Y(n_2904)
);

INVx4_ASAP7_75t_L g2905 ( 
.A(n_2781),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2743),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2745),
.A2(n_1137),
.B(n_1136),
.Y(n_2907)
);

A2O1A1Ixp33_ASAP7_75t_L g2908 ( 
.A1(n_2837),
.A2(n_1160),
.B(n_1163),
.C(n_1157),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2758),
.B(n_1165),
.Y(n_2909)
);

A2O1A1Ixp33_ASAP7_75t_L g2910 ( 
.A1(n_2836),
.A2(n_1172),
.B(n_1185),
.C(n_1166),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2760),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2786),
.B(n_1187),
.Y(n_2912)
);

INVx1_ASAP7_75t_SL g2913 ( 
.A(n_2796),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2791),
.B(n_1194),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2806),
.B(n_1201),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2740),
.A2(n_1206),
.B(n_1205),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2763),
.B(n_1210),
.Y(n_2917)
);

A2O1A1Ixp33_ASAP7_75t_L g2918 ( 
.A1(n_2747),
.A2(n_1214),
.B(n_1215),
.C(n_1212),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2756),
.Y(n_2919)
);

BUFx3_ASAP7_75t_L g2920 ( 
.A(n_2794),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2826),
.A2(n_2834),
.B(n_2754),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2756),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2809),
.Y(n_2923)
);

NOR2x1_ASAP7_75t_L g2924 ( 
.A(n_2749),
.B(n_1226),
.Y(n_2924)
);

OAI21xp33_ASAP7_75t_L g2925 ( 
.A1(n_2778),
.A2(n_1183),
.B(n_1182),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2766),
.B(n_1238),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2833),
.A2(n_1241),
.B(n_1239),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2813),
.Y(n_2928)
);

AOI33xp33_ASAP7_75t_L g2929 ( 
.A1(n_2812),
.A2(n_1255),
.A3(n_1245),
.B1(n_1257),
.B2(n_1246),
.B3(n_1243),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2762),
.A2(n_1191),
.B1(n_1192),
.B2(n_1190),
.Y(n_2930)
);

OAI22xp5_ASAP7_75t_L g2931 ( 
.A1(n_2842),
.A2(n_1200),
.B1(n_1202),
.B2(n_1193),
.Y(n_2931)
);

OAI21xp33_ASAP7_75t_L g2932 ( 
.A1(n_2798),
.A2(n_1211),
.B(n_1208),
.Y(n_2932)
);

O2A1O1Ixp33_ASAP7_75t_L g2933 ( 
.A1(n_2765),
.A2(n_1263),
.B(n_1272),
.C(n_1264),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2756),
.Y(n_2934)
);

OAI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2810),
.A2(n_1221),
.B1(n_1222),
.B2(n_1213),
.Y(n_2935)
);

INVxp67_ASAP7_75t_L g2936 ( 
.A(n_2718),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2839),
.A2(n_1227),
.B1(n_1231),
.B2(n_1224),
.Y(n_2937)
);

AOI21xp33_ASAP7_75t_L g2938 ( 
.A1(n_2790),
.A2(n_1236),
.B(n_1234),
.Y(n_2938)
);

O2A1O1Ixp33_ASAP7_75t_L g2939 ( 
.A1(n_2784),
.A2(n_1300),
.B(n_1311),
.C(n_1293),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2775),
.B(n_1314),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2782),
.Y(n_2941)
);

A2O1A1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2776),
.A2(n_1330),
.B(n_1338),
.C(n_1327),
.Y(n_2942)
);

AOI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2797),
.A2(n_1342),
.B(n_1340),
.Y(n_2943)
);

OR2x2_ASAP7_75t_SL g2944 ( 
.A(n_2815),
.B(n_1287),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_SL g2945 ( 
.A1(n_2831),
.A2(n_1316),
.B1(n_1364),
.B2(n_1256),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2788),
.Y(n_2946)
);

INVx3_ASAP7_75t_SL g2947 ( 
.A(n_2792),
.Y(n_2947)
);

INVx3_ASAP7_75t_L g2948 ( 
.A(n_2785),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2838),
.B(n_1256),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2789),
.Y(n_2950)
);

O2A1O1Ixp33_ASAP7_75t_L g2951 ( 
.A1(n_2787),
.A2(n_1353),
.B(n_1365),
.C(n_1351),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2804),
.B(n_1367),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2777),
.B(n_1370),
.Y(n_2953)
);

OAI21x1_ASAP7_75t_L g2954 ( 
.A1(n_2835),
.A2(n_1305),
.B(n_1287),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2768),
.Y(n_2955)
);

INVx5_ASAP7_75t_SL g2956 ( 
.A(n_2878),
.Y(n_2956)
);

AOI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2887),
.A2(n_2827),
.B1(n_2841),
.B2(n_2840),
.Y(n_2957)
);

INVx1_ASAP7_75t_SL g2958 ( 
.A(n_2864),
.Y(n_2958)
);

CKINVDCx20_ASAP7_75t_R g2959 ( 
.A(n_2853),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2844),
.A2(n_2803),
.B1(n_2823),
.B2(n_2783),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_2902),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2859),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_2888),
.Y(n_2963)
);

INVx4_ASAP7_75t_L g2964 ( 
.A(n_2947),
.Y(n_2964)
);

INVx5_ASAP7_75t_SL g2965 ( 
.A(n_2878),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2859),
.Y(n_2966)
);

BUFx4f_ASAP7_75t_L g2967 ( 
.A(n_2899),
.Y(n_2967)
);

BUFx12f_ASAP7_75t_L g2968 ( 
.A(n_2856),
.Y(n_2968)
);

CKINVDCx20_ASAP7_75t_R g2969 ( 
.A(n_2857),
.Y(n_2969)
);

NAND2x1p5_ASAP7_75t_L g2970 ( 
.A(n_2905),
.B(n_2822),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2850),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2847),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2848),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2858),
.Y(n_2974)
);

BUFx3_ASAP7_75t_L g2975 ( 
.A(n_2869),
.Y(n_2975)
);

INVx6_ASAP7_75t_L g2976 ( 
.A(n_2899),
.Y(n_2976)
);

INVx2_ASAP7_75t_SL g2977 ( 
.A(n_2890),
.Y(n_2977)
);

BUFx4f_ASAP7_75t_SL g2978 ( 
.A(n_2913),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2905),
.Y(n_2979)
);

BUFx12f_ASAP7_75t_L g2980 ( 
.A(n_2944),
.Y(n_2980)
);

BUFx8_ASAP7_75t_L g2981 ( 
.A(n_2899),
.Y(n_2981)
);

BUFx6f_ASAP7_75t_L g2982 ( 
.A(n_2920),
.Y(n_2982)
);

INVx5_ASAP7_75t_L g2983 ( 
.A(n_2865),
.Y(n_2983)
);

INVx2_ASAP7_75t_SL g2984 ( 
.A(n_2860),
.Y(n_2984)
);

NAND2x1p5_ASAP7_75t_L g2985 ( 
.A(n_2852),
.B(n_2780),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2868),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2897),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2889),
.Y(n_2988)
);

INVx2_ASAP7_75t_SL g2989 ( 
.A(n_2924),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2900),
.Y(n_2990)
);

INVx6_ASAP7_75t_SL g2991 ( 
.A(n_2843),
.Y(n_2991)
);

INVx6_ASAP7_75t_SL g2992 ( 
.A(n_2953),
.Y(n_2992)
);

BUFx3_ASAP7_75t_L g2993 ( 
.A(n_2906),
.Y(n_2993)
);

INVx5_ASAP7_75t_L g2994 ( 
.A(n_2893),
.Y(n_2994)
);

NAND2x1p5_ASAP7_75t_L g2995 ( 
.A(n_2950),
.B(n_2753),
.Y(n_2995)
);

INVx5_ASAP7_75t_SL g2996 ( 
.A(n_2953),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2911),
.Y(n_2997)
);

BUFx12f_ASAP7_75t_L g2998 ( 
.A(n_2955),
.Y(n_2998)
);

INVx6_ASAP7_75t_L g2999 ( 
.A(n_2936),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2909),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2912),
.Y(n_3001)
);

INVx8_ASAP7_75t_L g3002 ( 
.A(n_2948),
.Y(n_3002)
);

BUFx3_ASAP7_75t_L g3003 ( 
.A(n_2871),
.Y(n_3003)
);

BUFx12f_ASAP7_75t_L g3004 ( 
.A(n_2904),
.Y(n_3004)
);

INVx1_ASAP7_75t_SL g3005 ( 
.A(n_2854),
.Y(n_3005)
);

BUFx24_ASAP7_75t_L g3006 ( 
.A(n_2845),
.Y(n_3006)
);

INVx3_ASAP7_75t_L g3007 ( 
.A(n_2941),
.Y(n_3007)
);

INVx6_ASAP7_75t_L g3008 ( 
.A(n_2884),
.Y(n_3008)
);

INVx4_ASAP7_75t_L g3009 ( 
.A(n_2923),
.Y(n_3009)
);

BUFx3_ASAP7_75t_L g3010 ( 
.A(n_2896),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2914),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2915),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2866),
.Y(n_3013)
);

INVx4_ASAP7_75t_L g3014 ( 
.A(n_2928),
.Y(n_3014)
);

BUFx12f_ASAP7_75t_L g3015 ( 
.A(n_2929),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2946),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2851),
.B(n_2829),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2862),
.Y(n_3018)
);

INVx5_ASAP7_75t_L g3019 ( 
.A(n_2948),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2886),
.A2(n_2830),
.B1(n_1251),
.B2(n_1254),
.Y(n_3020)
);

INVx1_ASAP7_75t_SL g3021 ( 
.A(n_2882),
.Y(n_3021)
);

INVx4_ASAP7_75t_L g3022 ( 
.A(n_2919),
.Y(n_3022)
);

BUFx3_ASAP7_75t_L g3023 ( 
.A(n_2876),
.Y(n_3023)
);

INVx1_ASAP7_75t_SL g3024 ( 
.A(n_2903),
.Y(n_3024)
);

BUFx3_ASAP7_75t_L g3025 ( 
.A(n_2873),
.Y(n_3025)
);

NAND2x1p5_ASAP7_75t_L g3026 ( 
.A(n_2849),
.B(n_1378),
.Y(n_3026)
);

CKINVDCx8_ASAP7_75t_R g3027 ( 
.A(n_2870),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2877),
.Y(n_3028)
);

AO21x2_ASAP7_75t_L g3029 ( 
.A1(n_2880),
.A2(n_1389),
.B(n_1380),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2908),
.Y(n_3030)
);

INVx3_ASAP7_75t_L g3031 ( 
.A(n_2922),
.Y(n_3031)
);

BUFx4f_ASAP7_75t_L g3032 ( 
.A(n_2934),
.Y(n_3032)
);

BUFx5_ASAP7_75t_L g3033 ( 
.A(n_2861),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_2917),
.Y(n_3034)
);

INVx1_ASAP7_75t_SL g3035 ( 
.A(n_2926),
.Y(n_3035)
);

INVx1_ASAP7_75t_SL g3036 ( 
.A(n_2940),
.Y(n_3036)
);

INVx5_ASAP7_75t_SL g3037 ( 
.A(n_2910),
.Y(n_3037)
);

BUFx2_ASAP7_75t_L g3038 ( 
.A(n_2952),
.Y(n_3038)
);

INVx1_ASAP7_75t_SL g3039 ( 
.A(n_2894),
.Y(n_3039)
);

HB1xp67_ASAP7_75t_L g3040 ( 
.A(n_2846),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2907),
.Y(n_3041)
);

INVx3_ASAP7_75t_L g3042 ( 
.A(n_2954),
.Y(n_3042)
);

BUFx6f_ASAP7_75t_L g3043 ( 
.A(n_2949),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2891),
.Y(n_3044)
);

BUFx3_ASAP7_75t_L g3045 ( 
.A(n_2931),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_3015),
.A2(n_2925),
.B1(n_2938),
.B2(n_2874),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2971),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2972),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2958),
.B(n_2872),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2973),
.Y(n_3050)
);

NAND2x1p5_ASAP7_75t_L g3051 ( 
.A(n_3009),
.B(n_2867),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_2975),
.B(n_2916),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2974),
.Y(n_3053)
);

OAI21x1_ASAP7_75t_L g3054 ( 
.A1(n_3042),
.A2(n_2921),
.B(n_2863),
.Y(n_3054)
);

CKINVDCx11_ASAP7_75t_R g3055 ( 
.A(n_2959),
.Y(n_3055)
);

AO21x2_ASAP7_75t_L g3056 ( 
.A1(n_3029),
.A2(n_2927),
.B(n_2875),
.Y(n_3056)
);

OAI21x1_ASAP7_75t_L g3057 ( 
.A1(n_3041),
.A2(n_2943),
.B(n_2879),
.Y(n_3057)
);

OAI21x1_ASAP7_75t_L g3058 ( 
.A1(n_3026),
.A2(n_3031),
.B(n_2970),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_3032),
.A2(n_2895),
.B(n_2855),
.Y(n_3059)
);

AO31x2_ASAP7_75t_L g3060 ( 
.A1(n_3022),
.A2(n_2942),
.A3(n_2883),
.B(n_2918),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2978),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_3007),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2990),
.Y(n_3063)
);

CKINVDCx6p67_ASAP7_75t_R g3064 ( 
.A(n_2994),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_3005),
.B(n_2898),
.Y(n_3065)
);

BUFx3_ASAP7_75t_L g3066 ( 
.A(n_2999),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_2964),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_3018),
.B(n_2937),
.Y(n_3068)
);

OAI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_3017),
.A2(n_2881),
.B(n_2892),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2997),
.Y(n_3070)
);

OAI22xp5_ASAP7_75t_L g3071 ( 
.A1(n_3013),
.A2(n_2945),
.B1(n_2930),
.B2(n_2932),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2986),
.Y(n_3072)
);

AOI21xp5_ASAP7_75t_L g3073 ( 
.A1(n_3040),
.A2(n_2933),
.B(n_2901),
.Y(n_3073)
);

OAI21xp33_ASAP7_75t_SL g3074 ( 
.A1(n_2957),
.A2(n_2935),
.B(n_1407),
.Y(n_3074)
);

OR2x6_ASAP7_75t_L g3075 ( 
.A(n_2984),
.B(n_2885),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2988),
.Y(n_3076)
);

OAI21x1_ASAP7_75t_L g3077 ( 
.A1(n_2995),
.A2(n_2951),
.B(n_2939),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2983),
.B(n_1406),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3016),
.Y(n_3079)
);

AOI22x1_ASAP7_75t_L g3080 ( 
.A1(n_3014),
.A2(n_1260),
.B1(n_1261),
.B2(n_1259),
.Y(n_3080)
);

BUFx6f_ASAP7_75t_L g3081 ( 
.A(n_2967),
.Y(n_3081)
);

A2O1A1Ixp33_ASAP7_75t_L g3082 ( 
.A1(n_3045),
.A2(n_3020),
.B(n_3023),
.C(n_3034),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2993),
.Y(n_3083)
);

OA21x2_ASAP7_75t_L g3084 ( 
.A1(n_3044),
.A2(n_2960),
.B(n_3030),
.Y(n_3084)
);

INVx1_ASAP7_75t_SL g3085 ( 
.A(n_3008),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3019),
.Y(n_3086)
);

INVx5_ASAP7_75t_SL g3087 ( 
.A(n_2982),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_3019),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_3000),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_3025),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3028),
.Y(n_3091)
);

OAI21x1_ASAP7_75t_L g3092 ( 
.A1(n_2985),
.A2(n_1597),
.B(n_1309),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3002),
.Y(n_3093)
);

OAI21x1_ASAP7_75t_L g3094 ( 
.A1(n_3001),
.A2(n_1313),
.B(n_1305),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_3038),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3039),
.B(n_3035),
.Y(n_3096)
);

AND2x6_ASAP7_75t_L g3097 ( 
.A(n_3037),
.B(n_1313),
.Y(n_3097)
);

OAI21x1_ASAP7_75t_L g3098 ( 
.A1(n_2979),
.A2(n_1580),
.B(n_1344),
.Y(n_3098)
);

HB1xp67_ASAP7_75t_L g3099 ( 
.A(n_3011),
.Y(n_3099)
);

OAI21x1_ASAP7_75t_L g3100 ( 
.A1(n_3033),
.A2(n_1344),
.B(n_1332),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2998),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3043),
.Y(n_3102)
);

OAI21x1_ASAP7_75t_L g3103 ( 
.A1(n_3033),
.A2(n_2966),
.B(n_2962),
.Y(n_3103)
);

CKINVDCx5p33_ASAP7_75t_R g3104 ( 
.A(n_2961),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_3033),
.A2(n_1373),
.B(n_1332),
.Y(n_3105)
);

OAI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_3027),
.A2(n_1414),
.B1(n_1418),
.B2(n_1390),
.Y(n_3106)
);

OAI21x1_ASAP7_75t_L g3107 ( 
.A1(n_3006),
.A2(n_1418),
.B(n_1414),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_3043),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_3048),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3050),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_3053),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3079),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3072),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_3076),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3063),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3070),
.Y(n_3116)
);

AOI21x1_ASAP7_75t_L g3117 ( 
.A1(n_3073),
.A2(n_2989),
.B(n_1416),
.Y(n_3117)
);

BUFx3_ASAP7_75t_L g3118 ( 
.A(n_3066),
.Y(n_3118)
);

OAI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_3071),
.A2(n_3010),
.B1(n_2994),
.B2(n_2992),
.Y(n_3119)
);

HB1xp67_ASAP7_75t_L g3120 ( 
.A(n_3095),
.Y(n_3120)
);

OAI21x1_ASAP7_75t_L g3121 ( 
.A1(n_3054),
.A2(n_1445),
.B(n_1424),
.Y(n_3121)
);

HB1xp67_ASAP7_75t_L g3122 ( 
.A(n_3090),
.Y(n_3122)
);

INVx5_ASAP7_75t_SL g3123 ( 
.A(n_3081),
.Y(n_3123)
);

OA21x2_ASAP7_75t_L g3124 ( 
.A1(n_3057),
.A2(n_1432),
.B(n_1411),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_3089),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_3099),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_3047),
.Y(n_3127)
);

BUFx2_ASAP7_75t_L g3128 ( 
.A(n_3051),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_3068),
.A2(n_3004),
.B1(n_3012),
.B2(n_3003),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_3083),
.B(n_2982),
.Y(n_3130)
);

BUFx2_ASAP7_75t_L g3131 ( 
.A(n_3103),
.Y(n_3131)
);

INVx2_ASAP7_75t_SL g3132 ( 
.A(n_3064),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_SL g3133 ( 
.A1(n_3059),
.A2(n_2996),
.B1(n_2969),
.B2(n_3024),
.Y(n_3133)
);

BUFx2_ASAP7_75t_SL g3134 ( 
.A(n_3061),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3091),
.Y(n_3135)
);

NAND2x1p5_ASAP7_75t_L g3136 ( 
.A(n_3086),
.B(n_3036),
.Y(n_3136)
);

INVx2_ASAP7_75t_SL g3137 ( 
.A(n_3067),
.Y(n_3137)
);

INVx2_ASAP7_75t_SL g3138 ( 
.A(n_3102),
.Y(n_3138)
);

BUFx3_ASAP7_75t_L g3139 ( 
.A(n_3081),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_3062),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3084),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3088),
.Y(n_3142)
);

INVx3_ASAP7_75t_L g3143 ( 
.A(n_3085),
.Y(n_3143)
);

INVx1_ASAP7_75t_SL g3144 ( 
.A(n_3096),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3065),
.Y(n_3145)
);

BUFx3_ASAP7_75t_L g3146 ( 
.A(n_3108),
.Y(n_3146)
);

CKINVDCx20_ASAP7_75t_R g3147 ( 
.A(n_3055),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3078),
.Y(n_3148)
);

AND2x4_ASAP7_75t_L g3149 ( 
.A(n_3101),
.B(n_2963),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_3046),
.A2(n_2987),
.B1(n_3021),
.B2(n_2980),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_3058),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_3094),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3049),
.Y(n_3153)
);

HB1xp67_ASAP7_75t_SL g3154 ( 
.A(n_3104),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3100),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_3093),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_3105),
.Y(n_3157)
);

AND2x4_ASAP7_75t_SL g3158 ( 
.A(n_3147),
.B(n_3143),
.Y(n_3158)
);

INVx2_ASAP7_75t_SL g3159 ( 
.A(n_3156),
.Y(n_3159)
);

INVx6_ASAP7_75t_L g3160 ( 
.A(n_3156),
.Y(n_3160)
);

BUFx3_ASAP7_75t_L g3161 ( 
.A(n_3118),
.Y(n_3161)
);

CKINVDCx5p33_ASAP7_75t_R g3162 ( 
.A(n_3154),
.Y(n_3162)
);

CKINVDCx5p33_ASAP7_75t_R g3163 ( 
.A(n_3134),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_3119),
.A2(n_3082),
.B(n_3074),
.Y(n_3164)
);

NOR3xp33_ASAP7_75t_SL g3165 ( 
.A(n_3145),
.B(n_3106),
.C(n_3069),
.Y(n_3165)
);

OAI22xp5_ASAP7_75t_L g3166 ( 
.A1(n_3133),
.A2(n_3075),
.B1(n_3052),
.B2(n_2965),
.Y(n_3166)
);

CKINVDCx5p33_ASAP7_75t_R g3167 ( 
.A(n_3139),
.Y(n_3167)
);

OR2x6_ASAP7_75t_L g3168 ( 
.A(n_3128),
.B(n_3107),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_R g3169 ( 
.A(n_3132),
.B(n_2981),
.Y(n_3169)
);

O2A1O1Ixp33_ASAP7_75t_L g3170 ( 
.A1(n_3153),
.A2(n_3075),
.B(n_1445),
.C(n_1490),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_3130),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3109),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_3149),
.Y(n_3173)
);

NOR2x1p5_ASAP7_75t_L g3174 ( 
.A(n_3148),
.B(n_2968),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3110),
.Y(n_3175)
);

NAND2xp33_ASAP7_75t_R g3176 ( 
.A(n_3149),
.B(n_0),
.Y(n_3176)
);

HB1xp67_ASAP7_75t_L g3177 ( 
.A(n_3122),
.Y(n_3177)
);

AOI22xp33_ASAP7_75t_L g3178 ( 
.A1(n_3128),
.A2(n_3097),
.B1(n_3080),
.B2(n_3077),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_3129),
.A2(n_3150),
.B1(n_3136),
.B2(n_3144),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_3126),
.B(n_3097),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_3120),
.B(n_3087),
.Y(n_3181)
);

INVxp67_ASAP7_75t_L g3182 ( 
.A(n_3142),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3111),
.Y(n_3183)
);

NAND2xp33_ASAP7_75t_SL g3184 ( 
.A(n_3137),
.B(n_2977),
.Y(n_3184)
);

BUFx6f_ASAP7_75t_L g3185 ( 
.A(n_3146),
.Y(n_3185)
);

CKINVDCx5p33_ASAP7_75t_R g3186 ( 
.A(n_3138),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3112),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_3140),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_3114),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3113),
.B(n_2956),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3115),
.B(n_3092),
.Y(n_3191)
);

OAI22xp33_ASAP7_75t_L g3192 ( 
.A1(n_3117),
.A2(n_2991),
.B1(n_1490),
.B2(n_1504),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3116),
.Y(n_3193)
);

BUFx2_ASAP7_75t_L g3194 ( 
.A(n_3131),
.Y(n_3194)
);

CKINVDCx5p33_ASAP7_75t_R g3195 ( 
.A(n_3127),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_3135),
.B(n_3098),
.Y(n_3196)
);

CKINVDCx5p33_ASAP7_75t_R g3197 ( 
.A(n_3125),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_3141),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_3131),
.B(n_1435),
.Y(n_3199)
);

CKINVDCx16_ASAP7_75t_R g3200 ( 
.A(n_3123),
.Y(n_3200)
);

NAND2xp33_ASAP7_75t_SL g3201 ( 
.A(n_3123),
.B(n_1424),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3151),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3152),
.Y(n_3203)
);

BUFx2_ASAP7_75t_SL g3204 ( 
.A(n_3155),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_3157),
.B(n_3124),
.Y(n_3205)
);

INVx3_ASAP7_75t_L g3206 ( 
.A(n_3121),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3109),
.Y(n_3207)
);

OAI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_3133),
.A2(n_2976),
.B1(n_1556),
.B2(n_1504),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3144),
.B(n_1437),
.Y(n_3209)
);

AO31x2_ASAP7_75t_L g3210 ( 
.A1(n_3131),
.A2(n_1556),
.A3(n_1451),
.B(n_1452),
.Y(n_3210)
);

INVx2_ASAP7_75t_SL g3211 ( 
.A(n_3158),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3198),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3202),
.Y(n_3213)
);

AND2x4_ASAP7_75t_L g3214 ( 
.A(n_3177),
.B(n_3056),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_3172),
.Y(n_3215)
);

OR2x2_ASAP7_75t_L g3216 ( 
.A(n_3194),
.B(n_3060),
.Y(n_3216)
);

CKINVDCx20_ASAP7_75t_R g3217 ( 
.A(n_3162),
.Y(n_3217)
);

AO21x2_ASAP7_75t_L g3218 ( 
.A1(n_3199),
.A2(n_1455),
.B(n_1438),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3175),
.Y(n_3219)
);

INVx3_ASAP7_75t_L g3220 ( 
.A(n_3185),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_3183),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_3187),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_3207),
.Y(n_3223)
);

CKINVDCx5p33_ASAP7_75t_R g3224 ( 
.A(n_3163),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3193),
.Y(n_3225)
);

INVx3_ASAP7_75t_L g3226 ( 
.A(n_3185),
.Y(n_3226)
);

OR2x2_ASAP7_75t_L g3227 ( 
.A(n_3182),
.B(n_1467),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3189),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3197),
.Y(n_3229)
);

INVxp67_ASAP7_75t_SL g3230 ( 
.A(n_3180),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3203),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_SL g3232 ( 
.A1(n_3164),
.A2(n_3166),
.B1(n_3179),
.B2(n_3208),
.Y(n_3232)
);

OAI33xp33_ASAP7_75t_L g3233 ( 
.A1(n_3209),
.A2(n_1486),
.A3(n_1475),
.B1(n_1496),
.B2(n_1477),
.B3(n_1469),
.Y(n_3233)
);

OR2x2_ASAP7_75t_L g3234 ( 
.A(n_3195),
.B(n_1497),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3181),
.B(n_1505),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3196),
.Y(n_3236)
);

AOI221xp5_ASAP7_75t_L g3237 ( 
.A1(n_3170),
.A2(n_3165),
.B1(n_1532),
.B2(n_1541),
.C(n_1524),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_3174),
.B(n_3173),
.Y(n_3238)
);

OR2x2_ASAP7_75t_L g3239 ( 
.A(n_3204),
.B(n_3210),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3188),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3191),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3213),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3213),
.Y(n_3243)
);

AOI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3232),
.A2(n_3176),
.B1(n_3178),
.B2(n_3192),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3219),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3219),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3231),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3230),
.B(n_3171),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3236),
.B(n_3210),
.Y(n_3249)
);

BUFx3_ASAP7_75t_L g3250 ( 
.A(n_3217),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3212),
.Y(n_3251)
);

A2O1A1Ixp33_ASAP7_75t_L g3252 ( 
.A1(n_3237),
.A2(n_3201),
.B(n_3184),
.C(n_1560),
.Y(n_3252)
);

BUFx2_ASAP7_75t_L g3253 ( 
.A(n_3238),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3241),
.Y(n_3254)
);

NAND3xp33_ASAP7_75t_L g3255 ( 
.A(n_3214),
.B(n_3168),
.C(n_3205),
.Y(n_3255)
);

INVxp67_ASAP7_75t_SL g3256 ( 
.A(n_3239),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3233),
.A2(n_3190),
.B(n_3159),
.Y(n_3257)
);

NOR4xp25_ASAP7_75t_L g3258 ( 
.A(n_3234),
.B(n_3200),
.C(n_3206),
.D(n_1364),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3215),
.Y(n_3259)
);

OAI221xp5_ASAP7_75t_L g3260 ( 
.A1(n_3227),
.A2(n_3186),
.B1(n_3161),
.B2(n_3160),
.C(n_1269),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3221),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3222),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_SL g3263 ( 
.A(n_3238),
.B(n_3167),
.Y(n_3263)
);

OAI211xp5_ASAP7_75t_L g3264 ( 
.A1(n_3216),
.A2(n_1267),
.B(n_1273),
.C(n_1266),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3223),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_3220),
.B(n_3160),
.Y(n_3266)
);

OR2x2_ASAP7_75t_L g3267 ( 
.A(n_3228),
.B(n_2),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3225),
.Y(n_3268)
);

OR2x2_ASAP7_75t_L g3269 ( 
.A(n_3226),
.B(n_2),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3235),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3253),
.B(n_3211),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3248),
.B(n_3229),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_3258),
.B(n_3224),
.Y(n_3273)
);

NOR3xp33_ASAP7_75t_SL g3274 ( 
.A(n_3264),
.B(n_1277),
.C(n_1276),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3270),
.B(n_3218),
.Y(n_3275)
);

INVx2_ASAP7_75t_SL g3276 ( 
.A(n_3266),
.Y(n_3276)
);

BUFx2_ASAP7_75t_L g3277 ( 
.A(n_3256),
.Y(n_3277)
);

INVxp67_ASAP7_75t_SL g3278 ( 
.A(n_3249),
.Y(n_3278)
);

INVxp67_ASAP7_75t_L g3279 ( 
.A(n_3267),
.Y(n_3279)
);

NOR2xp67_ASAP7_75t_L g3280 ( 
.A(n_3255),
.B(n_3240),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3251),
.B(n_3169),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_3261),
.B(n_3262),
.Y(n_3282)
);

INVx1_ASAP7_75t_SL g3283 ( 
.A(n_3250),
.Y(n_3283)
);

BUFx3_ASAP7_75t_L g3284 ( 
.A(n_3269),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_3259),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3243),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3260),
.A2(n_1547),
.B1(n_1316),
.B2(n_1279),
.Y(n_3287)
);

OR2x2_ASAP7_75t_L g3288 ( 
.A(n_3265),
.B(n_3),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3268),
.B(n_1278),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_3263),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3245),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3254),
.B(n_4),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3246),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3247),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3257),
.B(n_1281),
.Y(n_3295)
);

OR2x2_ASAP7_75t_L g3296 ( 
.A(n_3252),
.B(n_5),
.Y(n_3296)
);

AOI221xp5_ASAP7_75t_L g3297 ( 
.A1(n_3258),
.A2(n_1289),
.B1(n_1290),
.B2(n_1285),
.C(n_1284),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3242),
.Y(n_3298)
);

NAND4xp75_ASAP7_75t_L g3299 ( 
.A(n_3244),
.B(n_1547),
.C(n_9),
.D(n_7),
.Y(n_3299)
);

OAI211xp5_ASAP7_75t_L g3300 ( 
.A1(n_3244),
.A2(n_1294),
.B(n_1301),
.C(n_1291),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3242),
.Y(n_3301)
);

AND2x4_ASAP7_75t_L g3302 ( 
.A(n_3276),
.B(n_8),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_3271),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3290),
.B(n_9),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3279),
.B(n_10),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3280),
.B(n_3284),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_3277),
.B(n_11),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3281),
.B(n_13),
.Y(n_3308)
);

INVx2_ASAP7_75t_SL g3309 ( 
.A(n_3272),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3285),
.B(n_13),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3278),
.B(n_15),
.Y(n_3311)
);

INVx1_ASAP7_75t_SL g3312 ( 
.A(n_3283),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3298),
.Y(n_3313)
);

BUFx2_ASAP7_75t_L g3314 ( 
.A(n_3275),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_3293),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3292),
.B(n_1302),
.Y(n_3316)
);

NOR3xp33_ASAP7_75t_L g3317 ( 
.A(n_3300),
.B(n_1318),
.C(n_1308),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3294),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_3273),
.B(n_1571),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3282),
.Y(n_3320)
);

BUFx2_ASAP7_75t_L g3321 ( 
.A(n_3288),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3289),
.B(n_1320),
.Y(n_3322)
);

AND2x2_ASAP7_75t_SL g3323 ( 
.A(n_3297),
.B(n_3296),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3286),
.B(n_16),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3301),
.Y(n_3325)
);

OR2x2_ASAP7_75t_L g3326 ( 
.A(n_3291),
.B(n_17),
.Y(n_3326)
);

AND3x1_ASAP7_75t_L g3327 ( 
.A(n_3274),
.B(n_1547),
.C(n_19),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3295),
.B(n_19),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3299),
.B(n_20),
.Y(n_3329)
);

CKINVDCx5p33_ASAP7_75t_R g3330 ( 
.A(n_3287),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3312),
.B(n_1321),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3303),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_3306),
.B(n_20),
.Y(n_3333)
);

INVx1_ASAP7_75t_SL g3334 ( 
.A(n_3307),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3309),
.B(n_22),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3321),
.B(n_22),
.Y(n_3336)
);

HB1xp67_ASAP7_75t_L g3337 ( 
.A(n_3315),
.Y(n_3337)
);

BUFx2_ASAP7_75t_L g3338 ( 
.A(n_3302),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_3330),
.B(n_1323),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3302),
.Y(n_3340)
);

INVx1_ASAP7_75t_SL g3341 ( 
.A(n_3304),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3311),
.B(n_1324),
.Y(n_3342)
);

INVxp67_ASAP7_75t_SL g3343 ( 
.A(n_3315),
.Y(n_3343)
);

INVxp67_ASAP7_75t_SL g3344 ( 
.A(n_3326),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3323),
.B(n_1325),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3308),
.B(n_23),
.Y(n_3346)
);

CKINVDCx16_ASAP7_75t_R g3347 ( 
.A(n_3329),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3318),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3320),
.B(n_24),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3328),
.B(n_3324),
.Y(n_3350)
);

NAND2x1p5_ASAP7_75t_L g3351 ( 
.A(n_3327),
.B(n_25),
.Y(n_3351)
);

HB1xp67_ASAP7_75t_L g3352 ( 
.A(n_3313),
.Y(n_3352)
);

INVx1_ASAP7_75t_SL g3353 ( 
.A(n_3305),
.Y(n_3353)
);

AND3x2_ASAP7_75t_L g3354 ( 
.A(n_3319),
.B(n_25),
.C(n_26),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3314),
.B(n_26),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3310),
.B(n_27),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3325),
.B(n_27),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3316),
.Y(n_3358)
);

NOR2xp33_ASAP7_75t_L g3359 ( 
.A(n_3322),
.B(n_1326),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3317),
.B(n_28),
.Y(n_3360)
);

OR2x2_ASAP7_75t_L g3361 ( 
.A(n_3321),
.B(n_28),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_3312),
.B(n_1328),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3312),
.B(n_1331),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3306),
.B(n_29),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3338),
.B(n_30),
.Y(n_3365)
);

OR2x2_ASAP7_75t_L g3366 ( 
.A(n_3334),
.B(n_30),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3333),
.Y(n_3367)
);

BUFx2_ASAP7_75t_L g3368 ( 
.A(n_3343),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3340),
.B(n_1334),
.Y(n_3369)
);

NOR2xp67_ASAP7_75t_L g3370 ( 
.A(n_3337),
.B(n_31),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3341),
.B(n_1337),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_3351),
.B(n_1341),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3353),
.B(n_1345),
.Y(n_3373)
);

OAI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3350),
.A2(n_1347),
.B1(n_1350),
.B2(n_1346),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3333),
.Y(n_3375)
);

BUFx2_ASAP7_75t_L g3376 ( 
.A(n_3344),
.Y(n_3376)
);

AO21x2_ASAP7_75t_L g3377 ( 
.A1(n_3345),
.A2(n_32),
.B(n_33),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3364),
.B(n_33),
.Y(n_3378)
);

OR2x2_ASAP7_75t_L g3379 ( 
.A(n_3332),
.B(n_34),
.Y(n_3379)
);

AO21x2_ASAP7_75t_L g3380 ( 
.A1(n_3355),
.A2(n_3336),
.B(n_3361),
.Y(n_3380)
);

INVx3_ASAP7_75t_SL g3381 ( 
.A(n_3346),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_3335),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3354),
.B(n_1357),
.Y(n_3383)
);

BUFx6f_ASAP7_75t_L g3384 ( 
.A(n_3349),
.Y(n_3384)
);

HB1xp67_ASAP7_75t_L g3385 ( 
.A(n_3352),
.Y(n_3385)
);

NOR3xp33_ASAP7_75t_L g3386 ( 
.A(n_3358),
.B(n_1361),
.C(n_1360),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_3358),
.A2(n_1363),
.B1(n_1374),
.B2(n_1362),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3356),
.B(n_34),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3357),
.Y(n_3389)
);

INVx5_ASAP7_75t_L g3390 ( 
.A(n_3360),
.Y(n_3390)
);

INVx1_ASAP7_75t_SL g3391 ( 
.A(n_3331),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3362),
.B(n_1377),
.Y(n_3392)
);

AND2x4_ASAP7_75t_SL g3393 ( 
.A(n_3339),
.B(n_36),
.Y(n_3393)
);

HB1xp67_ASAP7_75t_L g3394 ( 
.A(n_3348),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3359),
.A2(n_1382),
.B1(n_1387),
.B2(n_1381),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3363),
.B(n_37),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3342),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_3338),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3338),
.B(n_37),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3338),
.B(n_38),
.Y(n_3400)
);

HB1xp67_ASAP7_75t_L g3401 ( 
.A(n_3338),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3338),
.B(n_39),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3338),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3347),
.B(n_1388),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3338),
.Y(n_3405)
);

OR2x2_ASAP7_75t_L g3406 ( 
.A(n_3334),
.B(n_40),
.Y(n_3406)
);

INVx1_ASAP7_75t_SL g3407 ( 
.A(n_3338),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3347),
.B(n_1394),
.Y(n_3408)
);

INVx1_ASAP7_75t_SL g3409 ( 
.A(n_3338),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3401),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3398),
.Y(n_3411)
);

OAI31xp33_ASAP7_75t_L g3412 ( 
.A1(n_3376),
.A2(n_45),
.A3(n_42),
.B(n_43),
.Y(n_3412)
);

AND2x2_ASAP7_75t_SL g3413 ( 
.A(n_3368),
.B(n_45),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3385),
.Y(n_3414)
);

NOR2x1_ASAP7_75t_L g3415 ( 
.A(n_3370),
.B(n_3377),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3403),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3381),
.B(n_1395),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3407),
.B(n_3409),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3390),
.B(n_1399),
.Y(n_3419)
);

OR2x2_ASAP7_75t_L g3420 ( 
.A(n_3380),
.B(n_47),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3405),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3390),
.B(n_1402),
.Y(n_3422)
);

NOR2x1_ASAP7_75t_L g3423 ( 
.A(n_3366),
.B(n_48),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3390),
.B(n_1403),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3365),
.Y(n_3425)
);

AND2x4_ASAP7_75t_L g3426 ( 
.A(n_3367),
.B(n_50),
.Y(n_3426)
);

HB1xp67_ASAP7_75t_L g3427 ( 
.A(n_3375),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3382),
.B(n_1405),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3384),
.B(n_1409),
.Y(n_3429)
);

INVxp67_ASAP7_75t_SL g3430 ( 
.A(n_3372),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3389),
.B(n_1413),
.Y(n_3431)
);

OR2x2_ASAP7_75t_L g3432 ( 
.A(n_3391),
.B(n_48),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3399),
.B(n_1415),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3400),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3402),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3379),
.Y(n_3436)
);

INVxp67_ASAP7_75t_L g3437 ( 
.A(n_3406),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_3394),
.Y(n_3438)
);

OR2x2_ASAP7_75t_L g3439 ( 
.A(n_3404),
.B(n_52),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3397),
.B(n_1417),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3378),
.B(n_1419),
.Y(n_3441)
);

OR2x2_ASAP7_75t_L g3442 ( 
.A(n_3408),
.B(n_52),
.Y(n_3442)
);

OR2x2_ASAP7_75t_L g3443 ( 
.A(n_3369),
.B(n_53),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3388),
.B(n_1422),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3386),
.B(n_1426),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3387),
.B(n_1427),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3371),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3396),
.B(n_1431),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3373),
.A2(n_1434),
.B1(n_1436),
.B2(n_1433),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3383),
.Y(n_3450)
);

OR2x2_ASAP7_75t_L g3451 ( 
.A(n_3374),
.B(n_54),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3393),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3392),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3395),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3381),
.B(n_1439),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3381),
.B(n_1441),
.Y(n_3456)
);

OR2x2_ASAP7_75t_L g3457 ( 
.A(n_3407),
.B(n_57),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3398),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3401),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3381),
.B(n_1447),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3401),
.Y(n_3461)
);

AND2x4_ASAP7_75t_L g3462 ( 
.A(n_3398),
.B(n_59),
.Y(n_3462)
);

OR2x2_ASAP7_75t_L g3463 ( 
.A(n_3407),
.B(n_58),
.Y(n_3463)
);

INVx1_ASAP7_75t_SL g3464 ( 
.A(n_3398),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3381),
.B(n_1453),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3381),
.B(n_1456),
.Y(n_3466)
);

AND4x1_ASAP7_75t_L g3467 ( 
.A(n_3372),
.B(n_60),
.C(n_58),
.D(n_59),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3401),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3381),
.B(n_1458),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3398),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3390),
.B(n_1461),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3381),
.B(n_1462),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3381),
.B(n_1465),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3381),
.B(n_1466),
.Y(n_3474)
);

INVx2_ASAP7_75t_SL g3475 ( 
.A(n_3368),
.Y(n_3475)
);

AND2x4_ASAP7_75t_SL g3476 ( 
.A(n_3384),
.B(n_61),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3401),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3401),
.Y(n_3478)
);

AOI211xp5_ASAP7_75t_L g3479 ( 
.A1(n_3420),
.A2(n_1471),
.B(n_1472),
.C(n_1470),
.Y(n_3479)
);

OAI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3415),
.A2(n_3423),
.B(n_3413),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3471),
.A2(n_1479),
.B(n_1473),
.Y(n_3481)
);

AOI211xp5_ASAP7_75t_L g3482 ( 
.A1(n_3464),
.A2(n_1484),
.B(n_1487),
.C(n_1480),
.Y(n_3482)
);

OAI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3458),
.A2(n_1489),
.B1(n_1493),
.B2(n_1488),
.Y(n_3483)
);

INVx1_ASAP7_75t_SL g3484 ( 
.A(n_3476),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3470),
.B(n_1495),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3438),
.Y(n_3486)
);

OAI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3437),
.A2(n_1502),
.B(n_1500),
.Y(n_3487)
);

AOI32xp33_ASAP7_75t_L g3488 ( 
.A1(n_3411),
.A2(n_3478),
.A3(n_3477),
.B1(n_3468),
.B2(n_3459),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3462),
.Y(n_3489)
);

AOI221xp5_ASAP7_75t_L g3490 ( 
.A1(n_3414),
.A2(n_1507),
.B1(n_1509),
.B2(n_1506),
.C(n_1503),
.Y(n_3490)
);

INVx1_ASAP7_75t_SL g3491 ( 
.A(n_3457),
.Y(n_3491)
);

OR2x2_ASAP7_75t_L g3492 ( 
.A(n_3410),
.B(n_63),
.Y(n_3492)
);

OAI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_3425),
.A2(n_1517),
.B1(n_1519),
.B2(n_1510),
.Y(n_3493)
);

OAI221xp5_ASAP7_75t_L g3494 ( 
.A1(n_3412),
.A2(n_1527),
.B1(n_1529),
.B2(n_1526),
.C(n_1520),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3452),
.B(n_1533),
.Y(n_3495)
);

AOI22xp33_ASAP7_75t_L g3496 ( 
.A1(n_3421),
.A2(n_1535),
.B1(n_1537),
.B2(n_1534),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3427),
.Y(n_3497)
);

OAI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_3434),
.A2(n_1539),
.B1(n_1540),
.B2(n_1538),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3461),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3426),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3463),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3435),
.B(n_1543),
.Y(n_3502)
);

INVx1_ASAP7_75t_SL g3503 ( 
.A(n_3432),
.Y(n_3503)
);

OAI22xp5_ASAP7_75t_L g3504 ( 
.A1(n_3416),
.A2(n_1545),
.B1(n_1546),
.B2(n_1544),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3430),
.A2(n_1552),
.B(n_1548),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3450),
.B(n_1553),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3441),
.B(n_1555),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3426),
.Y(n_3508)
);

OAI21xp33_ASAP7_75t_L g3509 ( 
.A1(n_3453),
.A2(n_1558),
.B(n_1557),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3444),
.B(n_1559),
.Y(n_3510)
);

AOI21xp33_ASAP7_75t_L g3511 ( 
.A1(n_3436),
.A2(n_1577),
.B(n_1576),
.Y(n_3511)
);

AOI22xp5_ASAP7_75t_L g3512 ( 
.A1(n_3454),
.A2(n_1584),
.B1(n_1585),
.B2(n_1579),
.Y(n_3512)
);

OAI211xp5_ASAP7_75t_SL g3513 ( 
.A1(n_3447),
.A2(n_1591),
.B(n_1593),
.C(n_1589),
.Y(n_3513)
);

AOI322xp5_ASAP7_75t_L g3514 ( 
.A1(n_3419),
.A2(n_1595),
.A3(n_70),
.B1(n_67),
.B2(n_69),
.C1(n_65),
.C2(n_66),
.Y(n_3514)
);

OAI32xp33_ASAP7_75t_L g3515 ( 
.A1(n_3422),
.A2(n_68),
.A3(n_71),
.B1(n_67),
.B2(n_70),
.Y(n_3515)
);

OAI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3455),
.A2(n_66),
.B(n_68),
.Y(n_3516)
);

AOI21xp33_ASAP7_75t_SL g3517 ( 
.A1(n_3429),
.A2(n_71),
.B(n_72),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3460),
.B(n_72),
.Y(n_3518)
);

INVx1_ASAP7_75t_SL g3519 ( 
.A(n_3469),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3472),
.B(n_73),
.Y(n_3520)
);

AOI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_3473),
.A2(n_3428),
.B1(n_3431),
.B2(n_3417),
.Y(n_3521)
);

OAI21xp33_ASAP7_75t_L g3522 ( 
.A1(n_3424),
.A2(n_73),
.B(n_74),
.Y(n_3522)
);

AOI221xp5_ASAP7_75t_L g3523 ( 
.A1(n_3449),
.A2(n_92),
.B1(n_101),
.B2(n_83),
.C(n_74),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3448),
.B(n_75),
.Y(n_3524)
);

OR2x2_ASAP7_75t_L g3525 ( 
.A(n_3456),
.B(n_75),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_SL g3526 ( 
.A(n_3467),
.B(n_76),
.Y(n_3526)
);

AOI211xp5_ASAP7_75t_SL g3527 ( 
.A1(n_3465),
.A2(n_80),
.B(n_77),
.C(n_79),
.Y(n_3527)
);

OAI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_3466),
.A2(n_81),
.B1(n_77),
.B2(n_80),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3474),
.B(n_81),
.Y(n_3529)
);

OAI21xp33_ASAP7_75t_L g3530 ( 
.A1(n_3440),
.A2(n_82),
.B(n_83),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_L g3531 ( 
.A1(n_3451),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_3531)
);

OAI221xp5_ASAP7_75t_L g3532 ( 
.A1(n_3439),
.A2(n_89),
.B1(n_85),
.B2(n_88),
.C(n_90),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3433),
.B(n_89),
.Y(n_3533)
);

OAI32xp33_ASAP7_75t_L g3534 ( 
.A1(n_3443),
.A2(n_93),
.A3(n_95),
.B1(n_92),
.B2(n_94),
.Y(n_3534)
);

AOI32xp33_ASAP7_75t_L g3535 ( 
.A1(n_3446),
.A2(n_94),
.A3(n_91),
.B1(n_93),
.B2(n_96),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3442),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3445),
.B(n_91),
.Y(n_3537)
);

INVx3_ASAP7_75t_L g3538 ( 
.A(n_3462),
.Y(n_3538)
);

A2O1A1Ixp33_ASAP7_75t_L g3539 ( 
.A1(n_3415),
.A2(n_99),
.B(n_96),
.C(n_97),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3475),
.Y(n_3540)
);

OAI21xp33_ASAP7_75t_SL g3541 ( 
.A1(n_3415),
.A2(n_101),
.B(n_102),
.Y(n_3541)
);

NAND3xp33_ASAP7_75t_SL g3542 ( 
.A(n_3420),
.B(n_103),
.C(n_104),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3464),
.B(n_103),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_3413),
.B(n_105),
.Y(n_3544)
);

AOI32xp33_ASAP7_75t_L g3545 ( 
.A1(n_3415),
.A2(n_112),
.A3(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3464),
.B(n_110),
.Y(n_3546)
);

OAI322xp33_ASAP7_75t_L g3547 ( 
.A1(n_3420),
.A2(n_124),
.A3(n_122),
.B1(n_118),
.B2(n_112),
.C1(n_117),
.C2(n_119),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3438),
.Y(n_3548)
);

AOI32xp33_ASAP7_75t_L g3549 ( 
.A1(n_3415),
.A2(n_127),
.A3(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3438),
.Y(n_3550)
);

AOI221xp5_ASAP7_75t_SL g3551 ( 
.A1(n_3464),
.A2(n_131),
.B1(n_125),
.B2(n_126),
.C(n_132),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3464),
.B(n_133),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3438),
.Y(n_3553)
);

AOI21xp33_ASAP7_75t_L g3554 ( 
.A1(n_3464),
.A2(n_134),
.B(n_135),
.Y(n_3554)
);

AOI22xp5_ASAP7_75t_SL g3555 ( 
.A1(n_3464),
.A2(n_138),
.B1(n_135),
.B2(n_137),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3471),
.A2(n_139),
.B(n_140),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3464),
.B(n_141),
.Y(n_3557)
);

AOI222xp33_ASAP7_75t_L g3558 ( 
.A1(n_3415),
.A2(n_170),
.B1(n_149),
.B2(n_179),
.C1(n_159),
.C2(n_142),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3475),
.Y(n_3559)
);

O2A1O1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3420),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3418),
.B(n_145),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3452),
.B(n_147),
.Y(n_3562)
);

AOI22xp33_ASAP7_75t_L g3563 ( 
.A1(n_3418),
.A2(n_151),
.B1(n_148),
.B2(n_149),
.Y(n_3563)
);

AOI33xp33_ASAP7_75t_L g3564 ( 
.A1(n_3464),
.A2(n_153),
.A3(n_155),
.B1(n_151),
.B2(n_152),
.B3(n_154),
.Y(n_3564)
);

NAND3xp33_ASAP7_75t_L g3565 ( 
.A(n_3415),
.B(n_152),
.C(n_156),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3464),
.B(n_162),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3438),
.Y(n_3567)
);

OAI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3464),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3438),
.Y(n_3569)
);

INVxp67_ASAP7_75t_L g3570 ( 
.A(n_3415),
.Y(n_3570)
);

NAND2x1_ASAP7_75t_L g3571 ( 
.A(n_3415),
.B(n_169),
.Y(n_3571)
);

INVx1_ASAP7_75t_SL g3572 ( 
.A(n_3464),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3438),
.Y(n_3573)
);

OAI21xp5_ASAP7_75t_SL g3574 ( 
.A1(n_3415),
.A2(n_169),
.B(n_170),
.Y(n_3574)
);

AOI322xp5_ASAP7_75t_L g3575 ( 
.A1(n_3415),
.A2(n_176),
.A3(n_175),
.B1(n_173),
.B2(n_171),
.C1(n_172),
.C2(n_174),
.Y(n_3575)
);

INVx1_ASAP7_75t_SL g3576 ( 
.A(n_3464),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3438),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3438),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3438),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3418),
.B(n_177),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3438),
.Y(n_3581)
);

AOI22xp5_ASAP7_75t_L g3582 ( 
.A1(n_3464),
.A2(n_187),
.B1(n_181),
.B2(n_184),
.Y(n_3582)
);

OAI21xp33_ASAP7_75t_L g3583 ( 
.A1(n_3418),
.A2(n_188),
.B(n_189),
.Y(n_3583)
);

AOI322xp5_ASAP7_75t_L g3584 ( 
.A1(n_3415),
.A2(n_194),
.A3(n_193),
.B1(n_191),
.B2(n_188),
.C1(n_189),
.C2(n_192),
.Y(n_3584)
);

INVxp67_ASAP7_75t_L g3585 ( 
.A(n_3415),
.Y(n_3585)
);

NAND3xp33_ASAP7_75t_L g3586 ( 
.A(n_3415),
.B(n_193),
.C(n_194),
.Y(n_3586)
);

OAI21xp33_ASAP7_75t_SL g3587 ( 
.A1(n_3415),
.A2(n_195),
.B(n_196),
.Y(n_3587)
);

AOI221x1_ASAP7_75t_L g3588 ( 
.A1(n_3410),
.A2(n_198),
.B1(n_195),
.B2(n_197),
.C(n_199),
.Y(n_3588)
);

CKINVDCx14_ASAP7_75t_R g3589 ( 
.A(n_3418),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3438),
.Y(n_3590)
);

OAI31xp33_ASAP7_75t_L g3591 ( 
.A1(n_3420),
.A2(n_200),
.A3(n_197),
.B(n_198),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3438),
.Y(n_3592)
);

OAI221xp5_ASAP7_75t_L g3593 ( 
.A1(n_3420),
.A2(n_205),
.B1(n_202),
.B2(n_204),
.C(n_206),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3538),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3508),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3589),
.B(n_3538),
.Y(n_3596)
);

NOR2xp33_ASAP7_75t_L g3597 ( 
.A(n_3541),
.B(n_204),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3500),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3572),
.B(n_3576),
.Y(n_3599)
);

NAND3x1_ASAP7_75t_L g3600 ( 
.A(n_3480),
.B(n_208),
.C(n_209),
.Y(n_3600)
);

INVxp33_ASAP7_75t_L g3601 ( 
.A(n_3526),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3587),
.B(n_210),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3489),
.Y(n_3603)
);

CKINVDCx20_ASAP7_75t_R g3604 ( 
.A(n_3484),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3561),
.B(n_211),
.Y(n_3605)
);

AND2x4_ASAP7_75t_L g3606 ( 
.A(n_3497),
.B(n_211),
.Y(n_3606)
);

NAND3xp33_ASAP7_75t_L g3607 ( 
.A(n_3570),
.B(n_214),
.C(n_215),
.Y(n_3607)
);

OAI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3585),
.A2(n_218),
.B(n_217),
.Y(n_3608)
);

INVxp67_ASAP7_75t_L g3609 ( 
.A(n_3571),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3543),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3486),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3548),
.Y(n_3612)
);

CKINVDCx20_ASAP7_75t_R g3613 ( 
.A(n_3544),
.Y(n_3613)
);

OAI31xp33_ASAP7_75t_L g3614 ( 
.A1(n_3574),
.A2(n_224),
.A3(n_222),
.B(n_223),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3555),
.B(n_222),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3550),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3553),
.Y(n_3617)
);

OR2x2_ASAP7_75t_L g3618 ( 
.A(n_3540),
.B(n_223),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_3551),
.B(n_3558),
.Y(n_3619)
);

AND2x4_ASAP7_75t_L g3620 ( 
.A(n_3567),
.B(n_225),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3569),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3580),
.B(n_226),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3575),
.B(n_227),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3559),
.B(n_229),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3584),
.B(n_229),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3573),
.B(n_230),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3577),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3578),
.B(n_230),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3579),
.B(n_231),
.Y(n_3629)
);

INVx2_ASAP7_75t_SL g3630 ( 
.A(n_3581),
.Y(n_3630)
);

INVx3_ASAP7_75t_L g3631 ( 
.A(n_3590),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3592),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3527),
.B(n_232),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3491),
.B(n_234),
.Y(n_3634)
);

HB1xp67_ASAP7_75t_L g3635 ( 
.A(n_3503),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3545),
.B(n_236),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3549),
.B(n_238),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3488),
.B(n_238),
.Y(n_3638)
);

INVx1_ASAP7_75t_SL g3639 ( 
.A(n_3519),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3546),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3552),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3557),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3566),
.Y(n_3643)
);

AND2x2_ASAP7_75t_L g3644 ( 
.A(n_3501),
.B(n_239),
.Y(n_3644)
);

NOR2x1_ASAP7_75t_L g3645 ( 
.A(n_3565),
.B(n_3586),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3583),
.B(n_239),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3562),
.B(n_242),
.Y(n_3647)
);

OR2x2_ASAP7_75t_L g3648 ( 
.A(n_3542),
.B(n_243),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3536),
.B(n_244),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3518),
.B(n_245),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3495),
.B(n_246),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3492),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3499),
.B(n_247),
.Y(n_3653)
);

INVx2_ASAP7_75t_SL g3654 ( 
.A(n_3520),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3524),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3539),
.B(n_248),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3525),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3506),
.B(n_248),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3521),
.B(n_249),
.Y(n_3659)
);

NAND2xp33_ASAP7_75t_L g3660 ( 
.A(n_3535),
.B(n_250),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3529),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3533),
.Y(n_3662)
);

INVx1_ASAP7_75t_SL g3663 ( 
.A(n_3537),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3502),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3516),
.B(n_3554),
.Y(n_3665)
);

INVxp67_ASAP7_75t_L g3666 ( 
.A(n_3593),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3485),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3588),
.B(n_251),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3564),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3522),
.B(n_255),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3568),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3591),
.B(n_257),
.Y(n_3672)
);

OAI22xp5_ASAP7_75t_L g3673 ( 
.A1(n_3563),
.A2(n_3582),
.B1(n_3494),
.B2(n_3531),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3556),
.B(n_257),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3507),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_SL g3676 ( 
.A(n_3560),
.B(n_259),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3510),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3528),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3534),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3515),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3599),
.B(n_3479),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3609),
.B(n_3530),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3635),
.Y(n_3683)
);

NOR2xp33_ASAP7_75t_L g3684 ( 
.A(n_3601),
.B(n_3509),
.Y(n_3684)
);

OAI22xp33_ASAP7_75t_L g3685 ( 
.A1(n_3638),
.A2(n_3623),
.B1(n_3625),
.B2(n_3668),
.Y(n_3685)
);

INVx1_ASAP7_75t_SL g3686 ( 
.A(n_3596),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3639),
.B(n_3482),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3603),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3597),
.B(n_3496),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3602),
.B(n_3547),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_SL g3691 ( 
.A(n_3614),
.B(n_3517),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3631),
.Y(n_3692)
);

NAND3xp33_ASAP7_75t_SL g3693 ( 
.A(n_3613),
.B(n_3514),
.C(n_3523),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3654),
.B(n_3512),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3630),
.B(n_3490),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3620),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3620),
.B(n_3487),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3619),
.B(n_3532),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_3633),
.B(n_3513),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3605),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3676),
.A2(n_3483),
.B(n_3493),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3606),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3634),
.Y(n_3703)
);

OR2x2_ASAP7_75t_L g3704 ( 
.A(n_3595),
.B(n_3504),
.Y(n_3704)
);

OR2x2_ASAP7_75t_L g3705 ( 
.A(n_3598),
.B(n_3498),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3651),
.B(n_3505),
.Y(n_3706)
);

NOR3xp33_ASAP7_75t_L g3707 ( 
.A(n_3666),
.B(n_3511),
.C(n_3481),
.Y(n_3707)
);

OR2x2_ASAP7_75t_L g3708 ( 
.A(n_3648),
.B(n_260),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3606),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3624),
.B(n_261),
.Y(n_3710)
);

NOR2xp33_ASAP7_75t_L g3711 ( 
.A(n_3663),
.B(n_261),
.Y(n_3711)
);

INVx1_ASAP7_75t_SL g3712 ( 
.A(n_3600),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3618),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3644),
.Y(n_3714)
);

NOR3xp33_ASAP7_75t_L g3715 ( 
.A(n_3673),
.B(n_263),
.C(n_264),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3622),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3680),
.B(n_263),
.Y(n_3717)
);

NAND2xp33_ASAP7_75t_SL g3718 ( 
.A(n_3615),
.B(n_265),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3649),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3653),
.Y(n_3720)
);

HB1xp67_ASAP7_75t_L g3721 ( 
.A(n_3610),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3650),
.Y(n_3722)
);

OR2x2_ASAP7_75t_L g3723 ( 
.A(n_3611),
.B(n_265),
.Y(n_3723)
);

NAND2xp33_ASAP7_75t_L g3724 ( 
.A(n_3645),
.B(n_266),
.Y(n_3724)
);

BUFx2_ASAP7_75t_L g3725 ( 
.A(n_3652),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_L g3726 ( 
.A(n_3669),
.B(n_268),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3671),
.B(n_3659),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3612),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3661),
.B(n_268),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3616),
.B(n_269),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3617),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3621),
.Y(n_3732)
);

NAND2xp33_ASAP7_75t_SL g3733 ( 
.A(n_3656),
.B(n_276),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3627),
.Y(n_3734)
);

NOR2x1_ASAP7_75t_L g3735 ( 
.A(n_3607),
.B(n_280),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3632),
.Y(n_3736)
);

HB1xp67_ASAP7_75t_L g3737 ( 
.A(n_3608),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3626),
.Y(n_3738)
);

AND2x4_ASAP7_75t_L g3739 ( 
.A(n_3657),
.B(n_280),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3628),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3665),
.B(n_281),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3629),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3658),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3646),
.B(n_282),
.Y(n_3744)
);

INVx2_ASAP7_75t_SL g3745 ( 
.A(n_3664),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3647),
.Y(n_3746)
);

OAI31xp33_ASAP7_75t_L g3747 ( 
.A1(n_3636),
.A2(n_3637),
.A3(n_3672),
.B(n_3678),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3670),
.B(n_283),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3655),
.B(n_284),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3640),
.B(n_285),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3641),
.B(n_285),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3674),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3642),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3643),
.B(n_287),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3662),
.B(n_289),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3675),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3677),
.B(n_292),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3667),
.Y(n_3758)
);

NOR2xp33_ASAP7_75t_L g3759 ( 
.A(n_3660),
.B(n_293),
.Y(n_3759)
);

INVxp67_ASAP7_75t_SL g3760 ( 
.A(n_3596),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3599),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_3594),
.B(n_293),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3599),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3599),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3599),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3599),
.B(n_294),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3599),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3599),
.Y(n_3768)
);

INVx1_ASAP7_75t_SL g3769 ( 
.A(n_3599),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3599),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3599),
.B(n_295),
.Y(n_3771)
);

OR2x2_ASAP7_75t_L g3772 ( 
.A(n_3594),
.B(n_296),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_SL g3773 ( 
.A(n_3599),
.B(n_297),
.Y(n_3773)
);

OR3x1_ASAP7_75t_L g3774 ( 
.A(n_3679),
.B(n_297),
.C(n_298),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3599),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3599),
.B(n_299),
.Y(n_3776)
);

OR2x2_ASAP7_75t_L g3777 ( 
.A(n_3594),
.B(n_300),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3599),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3604),
.Y(n_3779)
);

AND2x2_ASAP7_75t_SL g3780 ( 
.A(n_3599),
.B(n_301),
.Y(n_3780)
);

INVx1_ASAP7_75t_SL g3781 ( 
.A(n_3599),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3594),
.B(n_302),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3604),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3599),
.B(n_305),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3599),
.B(n_305),
.Y(n_3785)
);

INVxp67_ASAP7_75t_SL g3786 ( 
.A(n_3596),
.Y(n_3786)
);

HB1xp67_ASAP7_75t_L g3787 ( 
.A(n_3609),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3779),
.B(n_306),
.Y(n_3788)
);

OAI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3783),
.A2(n_3769),
.B1(n_3781),
.B2(n_3683),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3780),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3696),
.B(n_309),
.Y(n_3791)
);

NOR2x1_ASAP7_75t_L g3792 ( 
.A(n_3774),
.B(n_309),
.Y(n_3792)
);

NOR3xp33_ASAP7_75t_L g3793 ( 
.A(n_3685),
.B(n_321),
.C(n_310),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3787),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3702),
.B(n_310),
.Y(n_3795)
);

NOR3xp33_ASAP7_75t_L g3796 ( 
.A(n_3682),
.B(n_325),
.C(n_314),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_3709),
.B(n_3712),
.Y(n_3797)
);

OR2x2_ASAP7_75t_L g3798 ( 
.A(n_3761),
.B(n_315),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3776),
.B(n_316),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3763),
.B(n_317),
.Y(n_3800)
);

INVxp67_ASAP7_75t_L g3801 ( 
.A(n_3690),
.Y(n_3801)
);

NOR4xp25_ASAP7_75t_L g3802 ( 
.A(n_3693),
.B(n_320),
.C(n_318),
.D(n_319),
.Y(n_3802)
);

BUFx4f_ASAP7_75t_SL g3803 ( 
.A(n_3686),
.Y(n_3803)
);

NAND2xp33_ASAP7_75t_L g3804 ( 
.A(n_3721),
.B(n_318),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3784),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3764),
.B(n_323),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3765),
.B(n_326),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3767),
.B(n_326),
.Y(n_3808)
);

AOI21xp5_ASAP7_75t_L g3809 ( 
.A1(n_3724),
.A2(n_328),
.B(n_329),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3768),
.B(n_330),
.Y(n_3810)
);

NAND4xp25_ASAP7_75t_SL g3811 ( 
.A(n_3770),
.B(n_337),
.C(n_347),
.D(n_330),
.Y(n_3811)
);

OAI221xp5_ASAP7_75t_SL g3812 ( 
.A1(n_3747),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3775),
.B(n_332),
.Y(n_3813)
);

NOR2xp67_ASAP7_75t_L g3814 ( 
.A(n_3778),
.B(n_335),
.Y(n_3814)
);

NOR3x1_ASAP7_75t_L g3815 ( 
.A(n_3725),
.B(n_336),
.C(n_339),
.Y(n_3815)
);

INVx2_ASAP7_75t_SL g3816 ( 
.A(n_3739),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3691),
.A2(n_340),
.B(n_341),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3710),
.B(n_343),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3766),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3771),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3692),
.B(n_343),
.Y(n_3821)
);

AOI322xp5_ASAP7_75t_L g3822 ( 
.A1(n_3698),
.A2(n_3715),
.A3(n_3726),
.B1(n_3760),
.B2(n_3786),
.C1(n_3733),
.C2(n_3737),
.Y(n_3822)
);

NAND4xp25_ASAP7_75t_L g3823 ( 
.A(n_3684),
.B(n_350),
.C(n_344),
.D(n_345),
.Y(n_3823)
);

NAND4xp25_ASAP7_75t_L g3824 ( 
.A(n_3687),
.B(n_351),
.C(n_345),
.D(n_350),
.Y(n_3824)
);

NAND4xp25_ASAP7_75t_L g3825 ( 
.A(n_3681),
.B(n_356),
.C(n_352),
.D(n_355),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3727),
.B(n_357),
.Y(n_3826)
);

XNOR2xp5_ASAP7_75t_L g3827 ( 
.A(n_3703),
.B(n_357),
.Y(n_3827)
);

OR2x2_ASAP7_75t_L g3828 ( 
.A(n_3717),
.B(n_358),
.Y(n_3828)
);

NAND4xp75_ASAP7_75t_L g3829 ( 
.A(n_3735),
.B(n_361),
.C(n_358),
.D(n_360),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3741),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3700),
.B(n_364),
.Y(n_3831)
);

NOR3xp33_ASAP7_75t_L g3832 ( 
.A(n_3718),
.B(n_366),
.C(n_367),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3762),
.Y(n_3833)
);

AOI311xp33_ASAP7_75t_L g3834 ( 
.A1(n_3688),
.A2(n_373),
.A3(n_370),
.B(n_372),
.C(n_374),
.Y(n_3834)
);

NOR2xp67_ASAP7_75t_L g3835 ( 
.A(n_3745),
.B(n_373),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3772),
.Y(n_3836)
);

NAND3xp33_ASAP7_75t_L g3837 ( 
.A(n_3707),
.B(n_374),
.C(n_376),
.Y(n_3837)
);

AND2x4_ASAP7_75t_L g3838 ( 
.A(n_3714),
.B(n_377),
.Y(n_3838)
);

NAND3xp33_ASAP7_75t_L g3839 ( 
.A(n_3728),
.B(n_378),
.C(n_379),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3732),
.B(n_378),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3719),
.B(n_379),
.Y(n_3841)
);

AOI211xp5_ASAP7_75t_L g3842 ( 
.A1(n_3699),
.A2(n_383),
.B(n_380),
.C(n_382),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3720),
.B(n_380),
.Y(n_3843)
);

OAI211xp5_ASAP7_75t_L g3844 ( 
.A1(n_3701),
.A2(n_386),
.B(n_384),
.C(n_385),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3777),
.Y(n_3845)
);

NOR3xp33_ASAP7_75t_L g3846 ( 
.A(n_3689),
.B(n_386),
.C(n_387),
.Y(n_3846)
);

NAND4xp25_ASAP7_75t_SL g3847 ( 
.A(n_3695),
.B(n_389),
.C(n_387),
.D(n_388),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3759),
.B(n_392),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3757),
.B(n_393),
.Y(n_3849)
);

NOR2x1_ASAP7_75t_SL g3850 ( 
.A(n_3773),
.B(n_394),
.Y(n_3850)
);

NOR2xp33_ASAP7_75t_L g3851 ( 
.A(n_3803),
.B(n_3785),
.Y(n_3851)
);

NOR3xp33_ASAP7_75t_L g3852 ( 
.A(n_3789),
.B(n_3694),
.C(n_3713),
.Y(n_3852)
);

AOI221xp5_ASAP7_75t_L g3853 ( 
.A1(n_3802),
.A2(n_3731),
.B1(n_3736),
.B2(n_3734),
.C(n_3753),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3835),
.Y(n_3854)
);

AOI321xp33_ASAP7_75t_L g3855 ( 
.A1(n_3797),
.A2(n_3756),
.A3(n_3758),
.B1(n_3738),
.B2(n_3742),
.C(n_3740),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_SL g3856 ( 
.A(n_3792),
.B(n_3711),
.Y(n_3856)
);

O2A1O1Ixp5_ASAP7_75t_L g3857 ( 
.A1(n_3790),
.A2(n_3697),
.B(n_3706),
.C(n_3752),
.Y(n_3857)
);

AOI32xp33_ASAP7_75t_L g3858 ( 
.A1(n_3794),
.A2(n_3716),
.A3(n_3722),
.B1(n_3743),
.B2(n_3746),
.Y(n_3858)
);

AOI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3804),
.A2(n_3749),
.B(n_3729),
.Y(n_3859)
);

NOR2xp33_ASAP7_75t_L g3860 ( 
.A(n_3816),
.B(n_3708),
.Y(n_3860)
);

OAI21xp5_ASAP7_75t_SL g3861 ( 
.A1(n_3801),
.A2(n_3705),
.B(n_3704),
.Y(n_3861)
);

NAND4xp25_ASAP7_75t_SL g3862 ( 
.A(n_3822),
.B(n_3730),
.C(n_3751),
.D(n_3750),
.Y(n_3862)
);

XOR2xp5_ASAP7_75t_L g3863 ( 
.A(n_3827),
.B(n_3782),
.Y(n_3863)
);

OAI221xp5_ASAP7_75t_SL g3864 ( 
.A1(n_3830),
.A2(n_3754),
.B1(n_3755),
.B2(n_3744),
.C(n_3748),
.Y(n_3864)
);

AOI221xp5_ASAP7_75t_L g3865 ( 
.A1(n_3812),
.A2(n_3723),
.B1(n_398),
.B2(n_394),
.C(n_395),
.Y(n_3865)
);

AOI222xp33_ASAP7_75t_L g3866 ( 
.A1(n_3805),
.A2(n_401),
.B1(n_404),
.B2(n_398),
.C1(n_399),
.C2(n_402),
.Y(n_3866)
);

AOI221xp5_ASAP7_75t_L g3867 ( 
.A1(n_3793),
.A2(n_404),
.B1(n_401),
.B2(n_402),
.C(n_405),
.Y(n_3867)
);

AOI221xp5_ASAP7_75t_L g3868 ( 
.A1(n_3796),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.C(n_408),
.Y(n_3868)
);

INVx5_ASAP7_75t_L g3869 ( 
.A(n_3806),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3814),
.B(n_409),
.Y(n_3870)
);

AOI221xp5_ASAP7_75t_L g3871 ( 
.A1(n_3846),
.A2(n_3836),
.B1(n_3845),
.B2(n_3833),
.C(n_3837),
.Y(n_3871)
);

NOR2xp33_ASAP7_75t_L g3872 ( 
.A(n_3825),
.B(n_409),
.Y(n_3872)
);

AOI221xp5_ASAP7_75t_L g3873 ( 
.A1(n_3817),
.A2(n_413),
.B1(n_410),
.B2(n_412),
.C(n_414),
.Y(n_3873)
);

OAI211xp5_ASAP7_75t_L g3874 ( 
.A1(n_3844),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_3874)
);

NAND3xp33_ASAP7_75t_SL g3875 ( 
.A(n_3832),
.B(n_415),
.C(n_417),
.Y(n_3875)
);

AOI222xp33_ASAP7_75t_L g3876 ( 
.A1(n_3819),
.A2(n_423),
.B1(n_425),
.B2(n_418),
.C1(n_419),
.C2(n_424),
.Y(n_3876)
);

AOI221xp5_ASAP7_75t_L g3877 ( 
.A1(n_3847),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.C(n_430),
.Y(n_3877)
);

OA22x2_ASAP7_75t_L g3878 ( 
.A1(n_3826),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_3878)
);

AOI221xp5_ASAP7_75t_L g3879 ( 
.A1(n_3820),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.C(n_434),
.Y(n_3879)
);

OAI221xp5_ASAP7_75t_L g3880 ( 
.A1(n_3800),
.A2(n_441),
.B1(n_438),
.B2(n_439),
.C(n_442),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3824),
.B(n_438),
.Y(n_3881)
);

AOI221xp5_ASAP7_75t_SL g3882 ( 
.A1(n_3809),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.C(n_445),
.Y(n_3882)
);

AOI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3788),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_3883)
);

NAND3xp33_ASAP7_75t_SL g3884 ( 
.A(n_3842),
.B(n_448),
.C(n_450),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3810),
.A2(n_450),
.B(n_453),
.Y(n_3885)
);

NOR2xp33_ASAP7_75t_R g3886 ( 
.A(n_3811),
.B(n_453),
.Y(n_3886)
);

OAI211xp5_ASAP7_75t_L g3887 ( 
.A1(n_3834),
.A2(n_458),
.B(n_454),
.C(n_457),
.Y(n_3887)
);

AOI211xp5_ASAP7_75t_L g3888 ( 
.A1(n_3807),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_3888)
);

INVx2_ASAP7_75t_SL g3889 ( 
.A(n_3838),
.Y(n_3889)
);

AOI211xp5_ASAP7_75t_L g3890 ( 
.A1(n_3808),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_3890)
);

AOI221xp5_ASAP7_75t_L g3891 ( 
.A1(n_3813),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.C(n_464),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3799),
.B(n_464),
.Y(n_3892)
);

AOI31xp33_ASAP7_75t_L g3893 ( 
.A1(n_3791),
.A2(n_3831),
.A3(n_3843),
.B(n_3841),
.Y(n_3893)
);

A2O1A1O1Ixp25_ASAP7_75t_L g3894 ( 
.A1(n_3821),
.A2(n_468),
.B(n_465),
.C(n_466),
.D(n_469),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3889),
.B(n_3795),
.Y(n_3895)
);

AO22x2_ASAP7_75t_L g3896 ( 
.A1(n_3854),
.A2(n_3829),
.B1(n_3828),
.B2(n_3840),
.Y(n_3896)
);

NAND3xp33_ASAP7_75t_SL g3897 ( 
.A(n_3886),
.B(n_3848),
.C(n_3849),
.Y(n_3897)
);

OAI22xp33_ASAP7_75t_L g3898 ( 
.A1(n_3856),
.A2(n_3818),
.B1(n_3839),
.B2(n_3798),
.Y(n_3898)
);

AOI222xp33_ASAP7_75t_L g3899 ( 
.A1(n_3853),
.A2(n_3850),
.B1(n_3838),
.B2(n_3815),
.C1(n_3823),
.C2(n_468),
.Y(n_3899)
);

NAND3xp33_ASAP7_75t_L g3900 ( 
.A(n_3894),
.B(n_465),
.C(n_466),
.Y(n_3900)
);

NAND3xp33_ASAP7_75t_L g3901 ( 
.A(n_3852),
.B(n_469),
.C(n_471),
.Y(n_3901)
);

OAI31xp33_ASAP7_75t_SL g3902 ( 
.A1(n_3851),
.A2(n_473),
.A3(n_471),
.B(n_472),
.Y(n_3902)
);

AOI221xp5_ASAP7_75t_L g3903 ( 
.A1(n_3887),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.C(n_478),
.Y(n_3903)
);

AOI222xp33_ASAP7_75t_L g3904 ( 
.A1(n_3871),
.A2(n_478),
.B1(n_480),
.B2(n_475),
.C1(n_476),
.C2(n_479),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3878),
.Y(n_3905)
);

OAI211xp5_ASAP7_75t_L g3906 ( 
.A1(n_3861),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_3906)
);

AND4x2_ASAP7_75t_L g3907 ( 
.A(n_3859),
.B(n_485),
.C(n_481),
.D(n_484),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3892),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3860),
.A2(n_488),
.B1(n_484),
.B2(n_486),
.Y(n_3909)
);

AOI211xp5_ASAP7_75t_L g3910 ( 
.A1(n_3874),
.A2(n_493),
.B(n_489),
.C(n_491),
.Y(n_3910)
);

NAND4xp25_ASAP7_75t_SL g3911 ( 
.A(n_3865),
.B(n_494),
.C(n_491),
.D(n_493),
.Y(n_3911)
);

NOR3xp33_ASAP7_75t_L g3912 ( 
.A(n_3857),
.B(n_3862),
.C(n_3864),
.Y(n_3912)
);

AOI221xp5_ASAP7_75t_L g3913 ( 
.A1(n_3893),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.C(n_497),
.Y(n_3913)
);

OAI211xp5_ASAP7_75t_SL g3914 ( 
.A1(n_3858),
.A2(n_497),
.B(n_495),
.C(n_496),
.Y(n_3914)
);

AOI221xp5_ASAP7_75t_L g3915 ( 
.A1(n_3884),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.C(n_501),
.Y(n_3915)
);

OAI211xp5_ASAP7_75t_L g3916 ( 
.A1(n_3855),
.A2(n_506),
.B(n_503),
.C(n_505),
.Y(n_3916)
);

OAI221xp5_ASAP7_75t_SL g3917 ( 
.A1(n_3863),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.C(n_509),
.Y(n_3917)
);

OAI322xp33_ASAP7_75t_L g3918 ( 
.A1(n_3870),
.A2(n_507),
.A3(n_508),
.B1(n_510),
.B2(n_511),
.C1(n_512),
.C2(n_513),
.Y(n_3918)
);

INVxp33_ASAP7_75t_SL g3919 ( 
.A(n_3872),
.Y(n_3919)
);

AOI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3881),
.A2(n_515),
.B1(n_512),
.B2(n_514),
.Y(n_3920)
);

OAI21xp33_ASAP7_75t_L g3921 ( 
.A1(n_3875),
.A2(n_516),
.B(n_517),
.Y(n_3921)
);

AO22x2_ASAP7_75t_L g3922 ( 
.A1(n_3885),
.A2(n_519),
.B1(n_516),
.B2(n_518),
.Y(n_3922)
);

OAI221xp5_ASAP7_75t_L g3923 ( 
.A1(n_3882),
.A2(n_522),
.B1(n_519),
.B2(n_520),
.C(n_523),
.Y(n_3923)
);

CKINVDCx20_ASAP7_75t_R g3924 ( 
.A(n_3895),
.Y(n_3924)
);

OAI221xp5_ASAP7_75t_L g3925 ( 
.A1(n_3902),
.A2(n_3873),
.B1(n_3877),
.B2(n_3867),
.C(n_3868),
.Y(n_3925)
);

OAI21xp5_ASAP7_75t_SL g3926 ( 
.A1(n_3899),
.A2(n_3903),
.B(n_3916),
.Y(n_3926)
);

NAND3xp33_ASAP7_75t_L g3927 ( 
.A(n_3912),
.B(n_3869),
.C(n_3888),
.Y(n_3927)
);

INVxp67_ASAP7_75t_L g3928 ( 
.A(n_3896),
.Y(n_3928)
);

AOI221xp5_ASAP7_75t_L g3929 ( 
.A1(n_3898),
.A2(n_3880),
.B1(n_3891),
.B2(n_3879),
.C(n_3890),
.Y(n_3929)
);

OAI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_3900),
.A2(n_3883),
.B1(n_3866),
.B2(n_3876),
.Y(n_3930)
);

AOI21xp33_ASAP7_75t_L g3931 ( 
.A1(n_3921),
.A2(n_524),
.B(n_526),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3915),
.B(n_526),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3907),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3896),
.Y(n_3934)
);

AND2x4_ASAP7_75t_L g3935 ( 
.A(n_3908),
.B(n_527),
.Y(n_3935)
);

O2A1O1Ixp33_ASAP7_75t_L g3936 ( 
.A1(n_3914),
.A2(n_3906),
.B(n_3905),
.C(n_3923),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3922),
.Y(n_3937)
);

NAND4xp75_ASAP7_75t_L g3938 ( 
.A(n_3937),
.B(n_3913),
.C(n_3920),
.D(n_3919),
.Y(n_3938)
);

AND2x2_ASAP7_75t_L g3939 ( 
.A(n_3933),
.B(n_3910),
.Y(n_3939)
);

OAI221xp5_ASAP7_75t_L g3940 ( 
.A1(n_3928),
.A2(n_3901),
.B1(n_3904),
.B2(n_3917),
.C(n_3909),
.Y(n_3940)
);

OAI311xp33_ASAP7_75t_L g3941 ( 
.A1(n_3926),
.A2(n_3897),
.A3(n_3911),
.B1(n_3918),
.C1(n_530),
.Y(n_3941)
);

OAI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3934),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_3942)
);

OAI211xp5_ASAP7_75t_SL g3943 ( 
.A1(n_3929),
.A2(n_533),
.B(n_531),
.C(n_532),
.Y(n_3943)
);

AND2x4_ASAP7_75t_L g3944 ( 
.A(n_3924),
.B(n_533),
.Y(n_3944)
);

AOI221x1_ASAP7_75t_L g3945 ( 
.A1(n_3927),
.A2(n_537),
.B1(n_534),
.B2(n_536),
.C(n_538),
.Y(n_3945)
);

CKINVDCx5p33_ASAP7_75t_R g3946 ( 
.A(n_3939),
.Y(n_3946)
);

INVx1_ASAP7_75t_SL g3947 ( 
.A(n_3944),
.Y(n_3947)
);

INVx1_ASAP7_75t_SL g3948 ( 
.A(n_3938),
.Y(n_3948)
);

BUFx2_ASAP7_75t_L g3949 ( 
.A(n_3942),
.Y(n_3949)
);

NAND3xp33_ASAP7_75t_SL g3950 ( 
.A(n_3940),
.B(n_3936),
.C(n_3930),
.Y(n_3950)
);

CKINVDCx5p33_ASAP7_75t_R g3951 ( 
.A(n_3941),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3949),
.Y(n_3952)
);

OAI22x1_ASAP7_75t_L g3953 ( 
.A1(n_3951),
.A2(n_3932),
.B1(n_3935),
.B2(n_3943),
.Y(n_3953)
);

OAI22xp5_ASAP7_75t_L g3954 ( 
.A1(n_3948),
.A2(n_3925),
.B1(n_3931),
.B2(n_3945),
.Y(n_3954)
);

AOI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3952),
.A2(n_3950),
.B1(n_3946),
.B2(n_3947),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3953),
.B(n_536),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3956),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3957),
.Y(n_3958)
);

OAI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3958),
.A2(n_3955),
.B(n_3954),
.Y(n_3959)
);

INVx2_ASAP7_75t_SL g3960 ( 
.A(n_3959),
.Y(n_3960)
);

AOI21xp5_ASAP7_75t_L g3961 ( 
.A1(n_3960),
.A2(n_546),
.B(n_547),
.Y(n_3961)
);

AOI322xp5_ASAP7_75t_L g3962 ( 
.A1(n_3961),
.A2(n_548),
.A3(n_549),
.B1(n_550),
.B2(n_551),
.C1(n_552),
.C2(n_553),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3962),
.A2(n_551),
.B(n_553),
.Y(n_3963)
);

AOI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3963),
.A2(n_559),
.B1(n_554),
.B2(n_558),
.Y(n_3964)
);

AOI211xp5_ASAP7_75t_L g3965 ( 
.A1(n_3964),
.A2(n_560),
.B(n_558),
.C(n_559),
.Y(n_3965)
);


endmodule