module real_jpeg_16125_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_523),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_0),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_1),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_1),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_1),
.B(n_243),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_2),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_2),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_3),
.B(n_190),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_3),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_3),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_3),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_3),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_3),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_3),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_4),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_4),
.B(n_55),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_4),
.B(n_288),
.Y(n_287)
);

AND2x4_ASAP7_75t_SL g301 ( 
.A(n_4),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g337 ( 
.A(n_4),
.B(n_243),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_5),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_5),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_5),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_5),
.A2(n_12),
.B1(n_274),
.B2(n_279),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_5),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_7),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_7),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_8),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_8),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_8),
.Y(n_343)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_8),
.Y(n_431)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_9),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_9),
.Y(n_336)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_9),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_10),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_11),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_11),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_11),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_11),
.B(n_67),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_11),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_11),
.B(n_299),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_11),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_11),
.B(n_276),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_12),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_12),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_12),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_12),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_12),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_12),
.B(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_12),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_12),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g98 ( 
.A(n_13),
.B(n_78),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_13),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_13),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_13),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_13),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_13),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_13),
.B(n_446),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_15),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_15),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_15),
.B(n_377),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_15),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_15),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_15),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_15),
.B(n_486),
.Y(n_485)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_16),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_16),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_16),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_18),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_18),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_171),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_169),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_143),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_23),
.B(n_143),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_103),
.C(n_116),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_24),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_74),
.C(n_89),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_26),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.C(n_58),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_27),
.B(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_35),
.C(n_40),
.Y(n_114)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_31),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_32),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_34),
.A2(n_35),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_35),
.B(n_106),
.C(n_109),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_40),
.A2(n_41),
.B1(n_92),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_92),
.C(n_94),
.Y(n_91)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_42),
.Y(n_486)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_43),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_44),
.B(n_58),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.C(n_54),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_45),
.B(n_54),
.Y(n_187)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_49),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_50),
.B(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_53),
.Y(n_251)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_57),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_64),
.C(n_69),
.Y(n_115)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_62),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_73),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_74),
.B(n_89),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_83),
.C(n_88),
.Y(n_142)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_99),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_90),
.A2(n_91),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_92),
.B(n_189),
.C(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_92),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_92),
.A2(n_192),
.B1(n_198),
.B2(n_226),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_93),
.Y(n_440)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_93),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_94),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_94),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_94),
.A2(n_195),
.B1(n_287),
.B2(n_331),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_96),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_97),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_98),
.B(n_99),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_98),
.B(n_242),
.C(n_247),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_98),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_99),
.A2(n_209),
.B1(n_210),
.B2(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_103),
.A2(n_116),
.B1(n_117),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.C(n_115),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_106),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_108),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_121),
.C(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_132),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_120),
.C(n_132),
.Y(n_168)
);

XOR2x1_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_124),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_131),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_138),
.C(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_168),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_158),
.B2(n_159),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_154),
.Y(n_305)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_154),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_214),
.B(n_519),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_173),
.A2(n_521),
.B(n_522),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_SL g522 ( 
.A(n_174),
.B(n_177),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_183),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_199),
.C(n_211),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_194),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_186),
.B(n_188),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_225),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_194),
.B(n_315),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_195),
.B(n_284),
.C(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_211),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_209),
.C(n_210),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_208),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_208),
.Y(n_239)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_263),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_260),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g521 ( 
.A(n_217),
.B(n_260),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_218),
.B(n_220),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_222),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_240),
.C(n_257),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_223),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_238),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_224),
.B(n_227),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_228),
.A2(n_233),
.B1(n_234),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_228),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_230),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_232),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_233),
.B(n_409),
.C(n_410),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_233),
.A2(n_234),
.B1(n_409),
.B2(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_SL g323 ( 
.A(n_238),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_240),
.B(n_257),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_250),
.C(n_252),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_241),
.B(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_247),
.Y(n_271)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_246),
.Y(n_446)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_250),
.A2(n_252),
.B1(n_253),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_252),
.A2(n_253),
.B1(n_389),
.B2(n_390),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_253),
.B(n_384),
.C(n_389),
.Y(n_383)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AO21x2_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_359),
.B(n_516),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_353),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_318),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_266),
.B(n_318),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_311),
.Y(n_266)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_267),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_292),
.C(n_306),
.Y(n_267)
);

INVxp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.C(n_283),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_270),
.B(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_272),
.A2(n_273),
.B1(n_283),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_273),
.A2(n_375),
.B(n_378),
.Y(n_374)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_283),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_330),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_292),
.A2(n_307),
.B1(n_308),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_300),
.C(n_303),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.C(n_298),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_294),
.A2(n_298),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_294),
.B(n_424),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_296),
.B(n_371),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_298),
.Y(n_373)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_299),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_300),
.A2(n_301),
.B1(n_303),
.B2(n_349),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_357),
.C(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_325),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_319),
.A2(n_320),
.B1(n_323),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_347),
.C(n_350),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.C(n_338),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_329),
.B(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_332),
.B(n_338),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_337),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.C(n_344),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_339),
.A2(n_342),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_342),
.A2(n_406),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_342),
.B(n_470),
.C(n_474),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_343),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_344),
.B(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_350),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_353),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

AND2x2_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_354),
.B(n_356),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_416),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.C(n_396),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_362),
.B(n_366),
.Y(n_515)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.C(n_392),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_393),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_374),
.C(n_383),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_374),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_372),
.B(n_425),
.C(n_428),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx12f_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_384),
.B(n_502),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

XNOR2x1_ASAP7_75t_SL g458 ( 
.A(n_385),
.B(n_388),
.Y(n_458)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_385),
.A2(n_465),
.B1(n_466),
.B2(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.C(n_414),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_512),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_402),
.B(n_414),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.C(n_412),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_403),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_408),
.B(n_413),
.Y(n_507)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_409),
.Y(n_454)
);

XOR2x1_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.C(n_515),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_510),
.B(n_514),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_496),
.B(n_509),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_461),
.B(n_495),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_449),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_449),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_432),
.C(n_441),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_428),
.Y(n_424)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_432),
.A2(n_433),
.B1(n_441),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_439),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_434),
.B(n_439),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

AO22x1_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_445),
.B1(n_447),
.B2(n_448),
.Y(n_441)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_442),
.Y(n_447)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_445),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_447),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_455),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_451),
.B(n_452),
.C(n_455),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_458),
.C(n_459),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_489),
.B(n_494),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_463),
.A2(n_477),
.B(n_488),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_469),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_466),
.Y(n_483)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_484),
.B(n_487),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_482),
.Y(n_487)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_493),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_493),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_508),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_497),
.B(n_508),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_499),
.B1(n_505),
.B2(n_506),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_503),
.B2(n_504),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_504),
.C(n_505),
.Y(n_513)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_513),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);


endmodule