module fake_jpeg_553_n_153 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_153);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_0),
.CON(n_42),
.SN(n_42)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_14),
.Y(n_68)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_66),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_20),
.B1(n_15),
.B2(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_20),
.B1(n_15),
.B2(n_16),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_16),
.B1(n_30),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_16),
.B1(n_23),
.B2(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_7),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_14),
.B1(n_16),
.B2(n_5),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_38),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_3),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_5),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_90),
.Y(n_107)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_11),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_65),
.C(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_70),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_109),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_81),
.B(n_78),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_101),
.B(n_96),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_63),
.B1(n_57),
.B2(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_83),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_77),
.C(n_83),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_69),
.B1(n_64),
.B2(n_56),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

OAI21x1_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_102),
.B(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_91),
.B1(n_81),
.B2(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_115),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_70),
.B(n_79),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_122),
.B(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_86),
.B(n_88),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_90),
.B1(n_56),
.B2(n_64),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_109),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_123),
.B(n_105),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_103),
.C(n_107),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_131),
.C(n_70),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_107),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_113),
.B(n_122),
.C(n_116),
.D(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_132),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_118),
.B1(n_125),
.B2(n_120),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g142 ( 
.A(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_141),
.C(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_120),
.B1(n_99),
.B2(n_57),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_140),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_147),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_135),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_149),
.A2(n_150),
.B(n_141),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_149),
.B(n_142),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_146),
.Y(n_153)
);


endmodule