module fake_jpeg_28223_n_278 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_42),
.B(n_15),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_20),
.B1(n_14),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_52),
.B1(n_60),
.B2(n_18),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_50),
.B1(n_59),
.B2(n_56),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_33),
.B1(n_30),
.B2(n_29),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_55),
.B1(n_35),
.B2(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_33),
.B1(n_19),
.B2(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_59),
.B1(n_18),
.B2(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_34),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_32),
.A2(n_17),
.B1(n_16),
.B2(n_21),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_61),
.A2(n_40),
.B(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_66),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_12),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_81),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_28),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_78),
.B1(n_49),
.B2(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_80),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_35),
.C(n_37),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_101),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_102),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_93),
.Y(n_110)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_78),
.B1(n_74),
.B2(n_80),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_37),
.C(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_58),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_45),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_109),
.B(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_112),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_61),
.B(n_65),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_77),
.C(n_68),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_115),
.C(n_36),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_101),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_61),
.B(n_62),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_118),
.B(n_87),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_61),
.B(n_35),
.C(n_34),
.D(n_37),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_25),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_71),
.B1(n_49),
.B2(n_64),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_98),
.B1(n_84),
.B2(n_99),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_34),
.B(n_37),
.C(n_36),
.D(n_31),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_89),
.B(n_36),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_87),
.B1(n_89),
.B2(n_96),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_93),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_95),
.B1(n_91),
.B2(n_86),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_140),
.B1(n_124),
.B2(n_120),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_86),
.B(n_83),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_142),
.B(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_141),
.B1(n_117),
.B2(n_121),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_94),
.B1(n_49),
.B2(n_99),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_83),
.B1(n_99),
.B2(n_98),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_115),
.C(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_149),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_164),
.C(n_172),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_111),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_161),
.Y(n_182)
);

AOI21x1_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_109),
.B(n_114),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_163),
.B1(n_132),
.B2(n_137),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_111),
.B1(n_114),
.B2(n_110),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_110),
.C(n_106),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_25),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_124),
.B1(n_120),
.B2(n_96),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_167),
.B1(n_144),
.B2(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_96),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_31),
.C(n_54),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_161),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_149),
.C(n_137),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_183),
.C(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_188),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_132),
.C(n_141),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_140),
.B1(n_147),
.B2(n_82),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_82),
.B1(n_41),
.B2(n_48),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_82),
.B1(n_41),
.B2(n_48),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_31),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_195),
.C(n_152),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_48),
.B1(n_27),
.B2(n_25),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_27),
.C(n_15),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_214),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_152),
.C(n_173),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_206),
.C(n_180),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_204),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_207),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_173),
.C(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_212),
.B1(n_153),
.B2(n_156),
.Y(n_215)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_178),
.B1(n_182),
.B2(n_193),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_196),
.B1(n_209),
.B2(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_175),
.B1(n_183),
.B2(n_186),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_226),
.B1(n_197),
.B2(n_204),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_185),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_224),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_225),
.C(n_227),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_195),
.C(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_229),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_192),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_160),
.Y(n_225)
);

NAND4xp25_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_166),
.C(n_9),
.D(n_10),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_15),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_27),
.C(n_8),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_209),
.C(n_210),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_225),
.C(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_235),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_205),
.B1(n_220),
.B2(n_9),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_6),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_245),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_244),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_205),
.C(n_6),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_248),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_247),
.B(n_0),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_254),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_13),
.B(n_12),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_10),
.B(n_9),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_10),
.Y(n_254)
);

AOI221xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_238),
.B1(n_237),
.B2(n_242),
.C(n_234),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_1),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_262),
.B(n_1),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_0),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_0),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_1),
.B(n_2),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_250),
.B(n_3),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_3),
.C(n_5),
.Y(n_273)
);

NOR2x1p5_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_3),
.C(n_4),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_253),
.C(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_270),
.C(n_1),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_273),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_267),
.B(n_269),
.C(n_5),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_274),
.B(n_5),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_275),
.Y(n_278)
);


endmodule