module fake_netlist_5_1786_n_189 (n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_189);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_189;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_29;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_188;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_102;
wire n_64;
wire n_106;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVxp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVxp33_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_R g58 ( 
.A(n_38),
.B(n_0),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_0),
.B(n_1),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_35),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp67_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_29),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_41),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_45),
.B1(n_48),
.B2(n_40),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI21x1_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_63),
.B(n_57),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_63),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_63),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_57),
.B(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_36),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_57),
.B(n_48),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_68),
.B(n_61),
.C(n_49),
.Y(n_98)
);

AOI21x1_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_68),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_56),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_59),
.B(n_36),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_94),
.B(n_96),
.C(n_76),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_76),
.B(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_77),
.B(n_87),
.Y(n_108)
);

OAI21x1_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_86),
.B(n_49),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_82),
.C(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_64),
.B1(n_39),
.B2(n_43),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_100),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_R g114 ( 
.A(n_106),
.B(n_92),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_105),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_105),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_105),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_92),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_96),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_109),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_85),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_126),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_58),
.C(n_46),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_44),
.B1(n_124),
.B2(n_122),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_131),
.Y(n_144)
);

OAI221xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_103),
.B1(n_124),
.B2(n_128),
.C(n_127),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_103),
.B(n_138),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_131),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_114),
.B(n_127),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_147),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_122),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_114),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_149),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_145),
.C(n_36),
.Y(n_161)
);

OAI211xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_158),
.B(n_152),
.C(n_150),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_143),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_150),
.B1(n_157),
.B2(n_151),
.C(n_153),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_157),
.A2(n_109),
.B(n_4),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

OAI211xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_2),
.B(n_9),
.C(n_10),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_77),
.C(n_79),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_11),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_11),
.B(n_13),
.C(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_16),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_18),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_19),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_20),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_170),
.B(n_166),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_169),
.B(n_171),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_177),
.B1(n_176),
.B2(n_172),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_180),
.B1(n_178),
.B2(n_106),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_180),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_187),
.A2(n_186),
.B1(n_184),
.B2(n_79),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_79),
.B1(n_106),
.B2(n_104),
.Y(n_189)
);


endmodule