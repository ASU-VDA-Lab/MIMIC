module fake_netlist_6_4602_n_2469 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2469);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2469;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2468;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_2127;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_1207;
wire n_811;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2357;
wire n_2025;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_107),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_48),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_121),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_132),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_18),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_83),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_8),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_143),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_122),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_99),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_142),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_84),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_88),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_71),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_105),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_69),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_226),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_194),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_89),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_160),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_29),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_133),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_187),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_13),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_125),
.Y(n_278)
);

BUFx8_ASAP7_75t_SL g279 ( 
.A(n_97),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_107),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_94),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_152),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_34),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_147),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_46),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_124),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_199),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_77),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_14),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_193),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_118),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_73),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_21),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_39),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_227),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_154),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_97),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_212),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_218),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_228),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_214),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_205),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_176),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_164),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_88),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_67),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_105),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_30),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_229),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_104),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_204),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_173),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_76),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_80),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_85),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_54),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_84),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_72),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_71),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_56),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_23),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_100),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_113),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_151),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_18),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_101),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_19),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_119),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_159),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_211),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_69),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_102),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_63),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_134),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_40),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_58),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_45),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_115),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_12),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_23),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_170),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_215),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_213),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_129),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_31),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_149),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_189),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_108),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_200),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_44),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_174),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_185),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_28),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_180),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_25),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_51),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_92),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_145),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_47),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_104),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_230),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_178),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_202),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_128),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_127),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_49),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_153),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_168),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_49),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_27),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_17),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_137),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_91),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_148),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_41),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_63),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_51),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_96),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_156),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_186),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_39),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_90),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_9),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_57),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_222),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_98),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_96),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_20),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_198),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_22),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_74),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_33),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_32),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_86),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_74),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_232),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_48),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_221),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_184),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_231),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_191),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_65),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_210),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_68),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_120),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_155),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_172),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_24),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_4),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_10),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_55),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_1),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_192),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_100),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_58),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_8),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_80),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_41),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_62),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_46),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_19),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_95),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_108),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_75),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_112),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_224),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_235),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_66),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_141),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_83),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_38),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_45),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_36),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_44),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_76),
.Y(n_441)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_60),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_181),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_68),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_40),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_52),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_81),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_162),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_93),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_24),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_94),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_131),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_53),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_27),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_91),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_166),
.Y(n_456)
);

BUFx2_ASAP7_75t_SL g457 ( 
.A(n_220),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_17),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_196),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_158),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_78),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_161),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_0),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_263),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_279),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_244),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_238),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_240),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_311),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_311),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_311),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_248),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_311),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_311),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_311),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_309),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_241),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_250),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_415),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_251),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_252),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_244),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_313),
.B(n_0),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_311),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_311),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_264),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_309),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_245),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_275),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g490 ( 
.A(n_236),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_311),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_424),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_283),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_354),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_285),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_442),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_287),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_321),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_288),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_294),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_302),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_304),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_305),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_255),
.B(n_1),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_245),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_442),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_314),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_246),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_442),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_328),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_321),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_317),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_329),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_333),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_255),
.B(n_2),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_352),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_335),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_R g525 ( 
.A(n_269),
.B(n_116),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_388),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_388),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_339),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_388),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_388),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_326),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_356),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_249),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_237),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_253),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_237),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_326),
.B(n_2),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_284),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_272),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_347),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_284),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_254),
.B(n_291),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_254),
.B(n_3),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_348),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_323),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_349),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_351),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_357),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_323),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_306),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_303),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_374),
.B(n_4),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_325),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_325),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_366),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_367),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_368),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_372),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_253),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_412),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_373),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_377),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_385),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_391),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_256),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_404),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_405),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_406),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_281),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_256),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_407),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_409),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_303),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_262),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_262),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_411),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_268),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_419),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_431),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_268),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_270),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_270),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_273),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_433),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_273),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_435),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_456),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_274),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_460),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_462),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_274),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_550),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_470),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_524),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_467),
.B(n_463),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_542),
.B(n_291),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_346),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_468),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_470),
.Y(n_600)
);

NOR2xp67_ASAP7_75t_L g601 ( 
.A(n_469),
.B(n_239),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_464),
.B(n_259),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_517),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_477),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_470),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_469),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_551),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_479),
.B(n_507),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_524),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_471),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_547),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_471),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_500),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_550),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_550),
.B(n_346),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_478),
.B(n_258),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_480),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_558),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_543),
.B(n_432),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_474),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_526),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_474),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_551),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_522),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_563),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_532),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_552),
.B(n_374),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_526),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_475),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_527),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_529),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_475),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_481),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_529),
.B(n_432),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_484),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_484),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_567),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_530),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_485),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_530),
.B(n_560),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_565),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_565),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_570),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_569),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_486),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_485),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_574),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_491),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_491),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_572),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_576),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_493),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_575),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_492),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_584),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_573),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_575),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_493),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_497),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_492),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_497),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_498),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_577),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_500),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_577),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_498),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_586),
.Y(n_674)
);

CKINVDCx16_ASAP7_75t_R g675 ( 
.A(n_479),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_R g676 ( 
.A(n_487),
.B(n_461),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_580),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_516),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_552),
.B(n_242),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_580),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_489),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_494),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_503),
.Y(n_683)
);

BUFx8_ASAP7_75t_L g684 ( 
.A(n_516),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_503),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_539),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_507),
.B(n_343),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_581),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_496),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_594),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_608),
.B(n_593),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_593),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_649),
.B(n_495),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_622),
.B(n_490),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_592),
.B(n_499),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_649),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_623),
.Y(n_697)
);

BUFx4f_ASAP7_75t_L g698 ( 
.A(n_606),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_623),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_623),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_686),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_679),
.B(n_560),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_592),
.B(n_615),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_602),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_594),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_600),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_622),
.B(n_501),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_592),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_606),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_594),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_602),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_625),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_625),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_608),
.B(n_502),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_592),
.B(n_504),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_598),
.A2(n_597),
.B(n_483),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_671),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_606),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_605),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_599),
.B(n_505),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_671),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_606),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_636),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_636),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_604),
.B(n_506),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_689),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_636),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_639),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_639),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_678),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_615),
.B(n_511),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_639),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_605),
.Y(n_734)
);

NAND3x1_ASAP7_75t_L g735 ( 
.A(n_598),
.B(n_277),
.C(n_276),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_678),
.B(n_512),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_597),
.B(n_533),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_640),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_679),
.A2(n_476),
.B1(n_560),
.B2(n_537),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_615),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_605),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_640),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_620),
.B(n_515),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_640),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_615),
.B(n_466),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_651),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_686),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_606),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_606),
.Y(n_749)
);

XNOR2xp5_ASAP7_75t_L g750 ( 
.A(n_602),
.B(n_408),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_596),
.B(n_495),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_600),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_661),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_651),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_596),
.B(n_518),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_689),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_630),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_612),
.B(n_520),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_619),
.B(n_523),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_611),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_630),
.Y(n_763)
);

INVx4_ASAP7_75t_SL g764 ( 
.A(n_611),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_600),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_630),
.B(n_466),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_637),
.B(n_528),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_600),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_651),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_644),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_650),
.B(n_540),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_681),
.B(n_544),
.Y(n_772)
);

INVx4_ASAP7_75t_SL g773 ( 
.A(n_611),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_653),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_653),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_679),
.B(n_482),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_616),
.B(n_546),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_612),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_616),
.B(n_548),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_653),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_616),
.B(n_555),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_659),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_659),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_659),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_676),
.Y(n_787)
);

XNOR2xp5_ASAP7_75t_L g788 ( 
.A(n_661),
.B(n_430),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_611),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_616),
.B(n_482),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_687),
.B(n_557),
.C(n_556),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_682),
.B(n_561),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_665),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_665),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_616),
.B(n_508),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_601),
.B(n_562),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_665),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_687),
.B(n_564),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_674),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_607),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_666),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_666),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_611),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_644),
.B(n_457),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_619),
.B(n_566),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_675),
.B(n_568),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_601),
.B(n_571),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_668),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_614),
.Y(n_810)
);

INVx4_ASAP7_75t_SL g811 ( 
.A(n_613),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_613),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_613),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_645),
.B(n_508),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_645),
.B(n_535),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_668),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_613),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_613),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_675),
.B(n_578),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_668),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_674),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_646),
.B(n_535),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_669),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_669),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_614),
.B(n_579),
.Y(n_825)
);

AND2x2_ASAP7_75t_SL g826 ( 
.A(n_638),
.B(n_334),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_607),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_646),
.B(n_559),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_669),
.B(n_587),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_676),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_614),
.A2(n_590),
.B1(n_589),
.B2(n_472),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_683),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_683),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_647),
.B(n_472),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_647),
.B(n_472),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_638),
.B(n_334),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_648),
.A2(n_537),
.B1(n_521),
.B2(n_265),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_683),
.B(n_509),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_685),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_614),
.B(n_472),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_667),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_R g842 ( 
.A(n_621),
.B(n_465),
.Y(n_842)
);

CKINVDCx14_ASAP7_75t_R g843 ( 
.A(n_667),
.Y(n_843)
);

OR2x2_ASAP7_75t_SL g844 ( 
.A(n_614),
.B(n_276),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_685),
.B(n_509),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_684),
.B(n_525),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_685),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_648),
.A2(n_521),
.B1(n_559),
.B2(n_459),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_607),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_613),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_607),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_690),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_690),
.Y(n_853)
);

AND2x6_ASAP7_75t_SL g854 ( 
.A(n_807),
.B(n_277),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_706),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_SL g856 ( 
.A1(n_750),
.A2(n_627),
.B1(n_629),
.B2(n_603),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_708),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_716),
.A2(n_694),
.B(n_707),
.C(n_790),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_714),
.B(n_684),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_708),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_705),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_706),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_770),
.B(n_613),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_696),
.B(n_621),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_706),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_628),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_745),
.B(n_617),
.Y(n_867)
);

AND2x6_ASAP7_75t_L g868 ( 
.A(n_790),
.B(n_242),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_765),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_765),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_798),
.B(n_684),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_778),
.B(n_684),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_759),
.A2(n_402),
.B1(n_684),
.B2(n_459),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_765),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_778),
.B(n_628),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_826),
.A2(n_247),
.B1(n_257),
.B2(n_243),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_745),
.B(n_617),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_826),
.A2(n_247),
.B1(n_257),
.B2(n_243),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_SL g879 ( 
.A(n_810),
.B(n_641),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_705),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_710),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_755),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_810),
.Y(n_883)
);

OAI22xp33_ASAP7_75t_L g884 ( 
.A1(n_691),
.A2(n_278),
.B1(n_292),
.B2(n_267),
.Y(n_884)
);

AND2x6_ASAP7_75t_SL g885 ( 
.A(n_720),
.B(n_286),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_836),
.B(n_267),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_759),
.A2(n_658),
.B(n_660),
.C(n_652),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_799),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_760),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_745),
.B(n_617),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_795),
.B(n_617),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_778),
.B(n_652),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_717),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_795),
.A2(n_457),
.B1(n_413),
.B2(n_292),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_800),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_836),
.B(n_617),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_763),
.B(n_641),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_800),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_766),
.B(n_655),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_702),
.B(n_617),
.Y(n_900)
);

AND2x6_ASAP7_75t_SL g901 ( 
.A(n_726),
.B(n_286),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_702),
.B(n_617),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_710),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_766),
.A2(n_513),
.B(n_514),
.C(n_510),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_815),
.B(n_618),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_693),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_766),
.B(n_658),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_815),
.B(n_618),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_815),
.B(n_655),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_787),
.B(n_657),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_740),
.B(n_618),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_740),
.B(n_618),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_743),
.B(n_657),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_767),
.B(n_662),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_842),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_779),
.A2(n_298),
.B1(n_299),
.B2(n_278),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_800),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_829),
.B(n_618),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_814),
.B(n_618),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_830),
.B(n_662),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_814),
.B(n_618),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_771),
.B(n_772),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_737),
.B(n_834),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_721),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_792),
.B(n_603),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_781),
.A2(n_298),
.B1(n_308),
.B2(n_299),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_783),
.A2(n_691),
.B1(n_805),
.B2(n_822),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_SL g928 ( 
.A1(n_750),
.A2(n_629),
.B1(n_627),
.B2(n_445),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_R g929 ( 
.A(n_780),
.B(n_436),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_737),
.B(n_343),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_721),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_822),
.B(n_633),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_736),
.B(n_583),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_791),
.B(n_488),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_703),
.A2(n_609),
.B(n_607),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_827),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_691),
.B(n_295),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_827),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_828),
.A2(n_513),
.B(n_514),
.C(n_510),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_691),
.A2(n_308),
.B1(n_359),
.B2(n_316),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_828),
.B(n_633),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_719),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_835),
.B(n_343),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_796),
.B(n_307),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_731),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_736),
.B(n_731),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_808),
.B(n_312),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_719),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_805),
.A2(n_697),
.B1(n_700),
.B2(n_699),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_805),
.B(n_660),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_827),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_780),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_851),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_734),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_805),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_695),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_SL g957 ( 
.A(n_727),
.B(n_449),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_851),
.B(n_633),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_851),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_715),
.B(n_633),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_732),
.B(n_850),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_697),
.B(n_633),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_699),
.B(n_633),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_698),
.A2(n_626),
.B(n_609),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_698),
.A2(n_626),
.B(n_609),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_739),
.B(n_307),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_755),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_752),
.A2(n_316),
.B1(n_363),
.B2(n_359),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_700),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_713),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_713),
.A2(n_363),
.B1(n_379),
.B2(n_369),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_848),
.B(n_664),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_757),
.B(n_355),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_722),
.B(n_633),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_837),
.A2(n_670),
.B(n_672),
.C(n_664),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_761),
.A2(n_369),
.B1(n_384),
.B2(n_379),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_722),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_724),
.B(n_643),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_724),
.B(n_643),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_725),
.A2(n_384),
.B1(n_448),
.B2(n_395),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_725),
.B(n_643),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_728),
.B(n_643),
.Y(n_982)
);

OAI221xp5_ASAP7_75t_L g983 ( 
.A1(n_840),
.A2(n_398),
.B1(n_300),
.B2(n_315),
.C(n_289),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_806),
.B(n_307),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_728),
.B(n_643),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_831),
.B(n_307),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_846),
.B(n_307),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_729),
.B(n_643),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_729),
.B(n_643),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_730),
.A2(n_448),
.B1(n_452),
.B2(n_395),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_701),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_SL g992 ( 
.A(n_701),
.B(n_266),
.C(n_261),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_727),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_730),
.B(n_654),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_727),
.B(n_758),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_734),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_SL g997 ( 
.A1(n_782),
.A2(n_793),
.B(n_794),
.C(n_784),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_758),
.B(n_443),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_733),
.B(n_654),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_733),
.B(n_738),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_819),
.A2(n_452),
.B1(n_672),
.B2(n_670),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_738),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_825),
.A2(n_290),
.B(n_289),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_742),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_758),
.B(n_443),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_SL g1006 ( 
.A1(n_704),
.A2(n_453),
.B1(n_451),
.B2(n_360),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_844),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_742),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_744),
.Y(n_1009)
);

AND2x6_ASAP7_75t_SL g1010 ( 
.A(n_788),
.B(n_290),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_782),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_744),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_841),
.B(n_396),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_774),
.B(n_654),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_711),
.B(n_438),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_L g1016 ( 
.A(n_718),
.B(n_303),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_821),
.B(n_271),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_774),
.B(n_654),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_776),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_741),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_784),
.B(n_677),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_747),
.B(n_280),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_776),
.B(n_654),
.Y(n_1023)
);

NOR2xp67_ASAP7_75t_L g1024 ( 
.A(n_747),
.B(n_677),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_785),
.B(n_786),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_741),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_858),
.B(n_922),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_857),
.B(n_680),
.Y(n_1028)
);

AND2x6_ASAP7_75t_L g1029 ( 
.A(n_950),
.B(n_718),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_886),
.B(n_718),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_869),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_857),
.B(n_680),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_969),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_855),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_855),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_969),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_862),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_862),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_865),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_924),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_886),
.B(n_718),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_860),
.B(n_688),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_869),
.Y(n_1044)
);

AND3x2_ASAP7_75t_SL g1045 ( 
.A(n_1006),
.B(n_1010),
.C(n_884),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_871),
.B(n_844),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_869),
.Y(n_1047)
);

INVx3_ASAP7_75t_SL g1048 ( 
.A(n_952),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_SL g1049 ( 
.A(n_928),
.B(n_788),
.C(n_293),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_956),
.B(n_907),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_956),
.B(n_785),
.Y(n_1051)
);

INVx5_ASAP7_75t_L g1052 ( 
.A(n_868),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_907),
.B(n_786),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_970),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_924),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_927),
.B(n_718),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_882),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_865),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_946),
.B(n_583),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_923),
.B(n_843),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_882),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_892),
.B(n_802),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_872),
.B(n_735),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_946),
.B(n_531),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_937),
.B(n_712),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_993),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_931),
.B(n_531),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_870),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_870),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_950),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_919),
.B(n_749),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_874),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_1013),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_970),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_892),
.B(n_688),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_874),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_895),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_947),
.B(n_802),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_868),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_955),
.B(n_735),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_906),
.B(n_746),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_875),
.B(n_756),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_895),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_977),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_SL g1085 ( 
.A(n_952),
.B(n_991),
.C(n_920),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_866),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_921),
.B(n_932),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_898),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_941),
.B(n_803),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_SL g1090 ( 
.A1(n_957),
.A2(n_360),
.B1(n_441),
.B2(n_260),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_868),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_898),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_977),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_991),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1002),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_897),
.B(n_769),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_993),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_917),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_931),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_868),
.A2(n_809),
.B1(n_820),
.B2(n_803),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_945),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1002),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_945),
.B(n_260),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_967),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_893),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_917),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_866),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_SL g1108 ( 
.A(n_929),
.B(n_297),
.C(n_282),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_891),
.B(n_809),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_973),
.B(n_310),
.C(n_301),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_R g1111 ( 
.A(n_889),
.B(n_318),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_900),
.B(n_820),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1015),
.B(n_832),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_905),
.B(n_749),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_967),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_902),
.B(n_832),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_936),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1008),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_950),
.B(n_764),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_955),
.B(n_764),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_972),
.B(n_839),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_868),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_933),
.B(n_260),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_936),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_972),
.B(n_839),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_938),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_1007),
.B(n_764),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_888),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_883),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_938),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_SL g1131 ( 
.A(n_910),
.B(n_320),
.C(n_319),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_868),
.A2(n_847),
.B1(n_794),
.B2(n_797),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_933),
.B(n_360),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_908),
.B(n_749),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1007),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_896),
.B(n_749),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_867),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_R g1138 ( 
.A(n_889),
.B(n_322),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_899),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_L g1140 ( 
.A(n_876),
.B(n_749),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_949),
.B(n_775),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_951),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_878),
.B(n_847),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_961),
.B(n_793),
.Y(n_1144)
);

INVx8_ASAP7_75t_L g1145 ( 
.A(n_1021),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_915),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_877),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_863),
.B(n_797),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_959),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_856),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_1021),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1024),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_959),
.B(n_764),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_890),
.B(n_775),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1008),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1009),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_915),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_909),
.B(n_581),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1009),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_918),
.B(n_775),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_934),
.B(n_801),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_913),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_1017),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_953),
.B(n_773),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1012),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1011),
.B(n_801),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_854),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1022),
.B(n_441),
.Y(n_1169)
);

NOR3xp33_ASAP7_75t_SL g1170 ( 
.A(n_864),
.B(n_327),
.C(n_324),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_930),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1012),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_1011),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_966),
.A2(n_823),
.B1(n_824),
.B2(n_816),
.Y(n_1174)
);

NOR2x1p5_ASAP7_75t_L g1175 ( 
.A(n_995),
.B(n_330),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_859),
.B(n_443),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_987),
.B(n_773),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_960),
.B(n_775),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1019),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1001),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_852),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_SL g1182 ( 
.A(n_983),
.B(n_340),
.C(n_331),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_SL g1183 ( 
.A(n_1003),
.B(n_345),
.C(n_342),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_887),
.B(n_816),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_883),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1019),
.B(n_823),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_885),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_904),
.B(n_775),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_914),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_879),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1004),
.B(n_824),
.Y(n_1191)
);

OR2x2_ASAP7_75t_SL g1192 ( 
.A(n_901),
.B(n_296),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_883),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_852),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_R g1195 ( 
.A(n_925),
.B(n_353),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_984),
.A2(n_723),
.B1(n_777),
.B2(n_751),
.Y(n_1196)
);

AND2x6_ASAP7_75t_L g1197 ( 
.A(n_873),
.B(n_789),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_853),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_853),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_943),
.B(n_441),
.Y(n_1200)
);

XNOR2xp5_ASAP7_75t_L g1201 ( 
.A(n_992),
.B(n_117),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_939),
.B(n_894),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_861),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_958),
.B(n_789),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_975),
.B(n_833),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_861),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_880),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_968),
.B(n_753),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_880),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_986),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_881),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_881),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_903),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_903),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_940),
.B(n_362),
.C(n_358),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_942),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_942),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_948),
.B(n_833),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_948),
.B(n_954),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_954),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_996),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_996),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_L g1223 ( 
.A(n_1066),
.B(n_998),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_L g1224 ( 
.A1(n_1027),
.A2(n_944),
.B(n_997),
.C(n_1005),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1033),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1067),
.B(n_916),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1033),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1113),
.B(n_1000),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1087),
.A2(n_698),
.B(n_911),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1161),
.A2(n_1178),
.B(n_1136),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1163),
.A2(n_976),
.B1(n_365),
.B2(n_376),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1152),
.A2(n_1180),
.B1(n_1145),
.B2(n_1163),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1037),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1113),
.B(n_1025),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1096),
.B(n_1020),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1094),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1096),
.B(n_1020),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1119),
.Y(n_1238)
);

AND2x6_ASAP7_75t_L g1239 ( 
.A(n_1122),
.B(n_1026),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1164),
.A2(n_926),
.B1(n_1016),
.B2(n_1026),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1119),
.Y(n_1241)
);

OAI22x1_ASAP7_75t_L g1242 ( 
.A1(n_1189),
.A2(n_378),
.B1(n_381),
.B2(n_364),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1205),
.A2(n_963),
.A3(n_974),
.B(n_962),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1161),
.A2(n_912),
.B(n_935),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1152),
.B(n_978),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1119),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1037),
.Y(n_1247)
);

INVx5_ASAP7_75t_L g1248 ( 
.A(n_1029),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1054),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1050),
.B(n_971),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1094),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1136),
.A2(n_1141),
.B(n_1202),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1178),
.A2(n_981),
.B(n_979),
.Y(n_1253)
);

NOR2x1_ASAP7_75t_SL g1254 ( 
.A(n_1079),
.B(n_789),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1141),
.A2(n_1125),
.B(n_1121),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1188),
.A2(n_985),
.B(n_982),
.Y(n_1256)
);

OA22x2_ASAP7_75t_L g1257 ( 
.A1(n_1189),
.A2(n_332),
.B1(n_336),
.B2(n_296),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1140),
.A2(n_751),
.B(n_723),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1152),
.B(n_723),
.Y(n_1259)
);

NOR4xp25_ASAP7_75t_L g1260 ( 
.A(n_1110),
.B(n_1169),
.C(n_1073),
.D(n_1108),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1105),
.B(n_980),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1044),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1065),
.B(n_990),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1188),
.A2(n_989),
.B(n_988),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1065),
.B(n_994),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1054),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1075),
.B(n_999),
.Y(n_1267)
);

NAND2x1_ASAP7_75t_L g1268 ( 
.A(n_1044),
.B(n_789),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1046),
.A2(n_336),
.B(n_337),
.C(n_332),
.Y(n_1269)
);

AND2x2_ASAP7_75t_SL g1270 ( 
.A(n_1091),
.B(n_1140),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1204),
.A2(n_1018),
.B(n_1014),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1128),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1145),
.A2(n_1023),
.B1(n_965),
.B2(n_964),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1204),
.A2(n_845),
.B(n_838),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_SL g1275 ( 
.A1(n_1184),
.A2(n_1016),
.B(n_370),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1075),
.B(n_753),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1086),
.B(n_582),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1030),
.A2(n_768),
.B(n_754),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1030),
.A2(n_768),
.B(n_754),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1123),
.B(n_582),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1091),
.A2(n_338),
.B(n_337),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1074),
.A2(n_338),
.A3(n_383),
.B(n_392),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1084),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1070),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1075),
.B(n_849),
.Y(n_1285)
);

NOR2x1_ASAP7_75t_L g1286 ( 
.A(n_1066),
.B(n_751),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1078),
.B(n_849),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1084),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1071),
.A2(n_610),
.B(n_595),
.Y(n_1289)
);

BUFx8_ASAP7_75t_L g1290 ( 
.A(n_1061),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1081),
.B(n_595),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1071),
.A2(n_624),
.B(n_610),
.Y(n_1292)
);

BUFx5_ASAP7_75t_L g1293 ( 
.A(n_1029),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1173),
.A2(n_818),
.B(n_777),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1081),
.B(n_624),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1107),
.B(n_386),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_SL g1297 ( 
.A1(n_1056),
.A2(n_591),
.B(n_585),
.C(n_588),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1093),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1093),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1059),
.B(n_585),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1042),
.A2(n_1062),
.B(n_1053),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1048),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1079),
.B(n_777),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1056),
.A2(n_632),
.B(n_631),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1095),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1173),
.A2(n_818),
.B(n_812),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1145),
.B(n_631),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1155),
.A2(n_634),
.B(n_632),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1102),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1133),
.B(n_588),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1046),
.A2(n_361),
.B(n_447),
.C(n_446),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1173),
.A2(n_818),
.B(n_812),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1042),
.A2(n_519),
.B(n_634),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1173),
.A2(n_812),
.B(n_789),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1109),
.A2(n_813),
.B(n_812),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1155),
.A2(n_642),
.B(n_635),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1145),
.B(n_635),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1102),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1048),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1082),
.A2(n_429),
.B(n_344),
.C(n_350),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1044),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1162),
.B(n_642),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1144),
.A2(n_1089),
.B(n_1079),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1079),
.A2(n_813),
.B(n_812),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1051),
.B(n_813),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1082),
.B(n_813),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1035),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1112),
.A2(n_519),
.B(n_609),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1114),
.A2(n_573),
.B(n_609),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1060),
.A2(n_1139),
.B1(n_1063),
.B2(n_1210),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1114),
.A2(n_656),
.B(n_626),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1134),
.A2(n_656),
.B(n_626),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1035),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1137),
.B(n_813),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1118),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1103),
.B(n_591),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1137),
.B(n_817),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_SL g1338 ( 
.A1(n_1091),
.A2(n_344),
.B(n_341),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1079),
.A2(n_817),
.B(n_748),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1179),
.A2(n_1156),
.B(n_1157),
.C(n_1118),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1134),
.A2(n_656),
.B(n_626),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1116),
.A2(n_817),
.B(n_748),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1156),
.Y(n_1343)
);

NAND2x1_ASAP7_75t_L g1344 ( 
.A(n_1047),
.B(n_817),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1130),
.A2(n_663),
.B(n_656),
.Y(n_1345)
);

BUFx8_ASAP7_75t_L g1346 ( 
.A(n_1104),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1149),
.A2(n_817),
.B(n_748),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1130),
.A2(n_663),
.B(n_656),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1130),
.A2(n_663),
.B(n_536),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1186),
.A2(n_1160),
.B(n_1157),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1090),
.A2(n_350),
.B(n_341),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1060),
.Y(n_1352)
);

INVx6_ASAP7_75t_L g1353 ( 
.A(n_1035),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1137),
.B(n_1148),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1137),
.B(n_654),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1052),
.A2(n_748),
.B(n_709),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1160),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1166),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1115),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1052),
.A2(n_748),
.B(n_709),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1166),
.A2(n_1172),
.B1(n_1148),
.B2(n_1052),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1052),
.B(n_1070),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1172),
.Y(n_1363)
);

AO21x1_ASAP7_75t_L g1364 ( 
.A1(n_1143),
.A2(n_371),
.B(n_361),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1070),
.B(n_709),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1035),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1219),
.A2(n_663),
.B(n_709),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1148),
.A2(n_443),
.B1(n_387),
.B2(n_389),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1142),
.A2(n_663),
.B(n_536),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1148),
.B(n_1028),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1028),
.B(n_654),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1047),
.A2(n_762),
.B(n_709),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1047),
.A2(n_804),
.B(n_762),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_SL g1374 ( 
.A(n_1097),
.Y(n_1374)
);

AOI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1064),
.A2(n_1171),
.B(n_1200),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1028),
.B(n_673),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1194),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1212),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1132),
.A2(n_804),
.B(n_762),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1195),
.B(n_534),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1142),
.A2(n_538),
.B(n_534),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1032),
.B(n_673),
.Y(n_1382)
);

INVx5_ASAP7_75t_L g1383 ( 
.A(n_1029),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1032),
.B(n_673),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1034),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1043),
.B(n_673),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1036),
.A2(n_429),
.A3(n_371),
.B(n_380),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1236),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1272),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1275),
.A2(n_1191),
.B(n_1218),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1228),
.B(n_1043),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1336),
.B(n_1280),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1263),
.A2(n_1183),
.B(n_1182),
.C(n_1215),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1225),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1225),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1252),
.A2(n_1208),
.B(n_1196),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1275),
.A2(n_1142),
.B(n_1167),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1378),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1247),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1247),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1283),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1369),
.A2(n_1031),
.B(n_1207),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1369),
.A2(n_1031),
.B(n_1207),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1277),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1248),
.B(n_1122),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1378),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1262),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1234),
.B(n_1043),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1375),
.A2(n_1153),
.B(n_1063),
.C(n_1190),
.Y(n_1409)
);

OR2x6_ASAP7_75t_SL g1410 ( 
.A(n_1232),
.B(n_1146),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1353),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1283),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1310),
.B(n_1226),
.Y(n_1413)
);

CKINVDCx12_ASAP7_75t_R g1414 ( 
.A(n_1300),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1236),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1224),
.A2(n_1100),
.B(n_1174),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1354),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1290),
.A2(n_1195),
.B1(n_1151),
.B2(n_1045),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1231),
.A2(n_1063),
.B1(n_1080),
.B2(n_1135),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1244),
.A2(n_1329),
.B(n_1332),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1244),
.A2(n_1031),
.B(n_1207),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1265),
.B(n_1370),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1298),
.B(n_1063),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1298),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1364),
.A2(n_1311),
.A3(n_1269),
.B(n_1340),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1367),
.A2(n_1039),
.B(n_1038),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1323),
.A2(n_1176),
.B(n_1209),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1238),
.B(n_1070),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1305),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1270),
.A2(n_1176),
.B1(n_1055),
.B2(n_1099),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1329),
.A2(n_1221),
.B(n_1198),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1305),
.Y(n_1432)
);

CKINVDCx14_ASAP7_75t_R g1433 ( 
.A(n_1251),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1332),
.A2(n_1221),
.B(n_1198),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1224),
.A2(n_1216),
.B(n_1213),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1248),
.B(n_1122),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1359),
.B(n_1146),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1255),
.A2(n_1222),
.B(n_1058),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1269),
.A2(n_1131),
.B(n_1170),
.C(n_1159),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1341),
.A2(n_1230),
.B(n_1349),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1341),
.A2(n_1221),
.B(n_1217),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1304),
.A2(n_1068),
.B(n_1040),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1353),
.Y(n_1443)
);

INVx5_ASAP7_75t_L g1444 ( 
.A(n_1248),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1357),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1304),
.A2(n_1072),
.B(n_1069),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1248),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_L g1448 ( 
.A(n_1238),
.B(n_1041),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1229),
.A2(n_1176),
.B(n_1077),
.Y(n_1449)
);

AO31x2_ASAP7_75t_L g1450 ( 
.A1(n_1311),
.A2(n_1340),
.A3(n_1320),
.B(n_1273),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1230),
.A2(n_1083),
.B(n_1076),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1261),
.A2(n_1085),
.B(n_1049),
.C(n_1101),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1380),
.A2(n_1080),
.B1(n_1176),
.B2(n_1175),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1256),
.A2(n_1092),
.B(n_1088),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1301),
.A2(n_1106),
.B(n_1098),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1235),
.B(n_1158),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1327),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1357),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1326),
.A2(n_1124),
.B(n_1117),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1256),
.A2(n_1217),
.B(n_1194),
.Y(n_1460)
);

AOI211xp5_ASAP7_75t_L g1461 ( 
.A1(n_1351),
.A2(n_1201),
.B(n_1168),
.C(n_1138),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1377),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1327),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1330),
.A2(n_1045),
.B(n_1185),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1377),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1250),
.A2(n_1147),
.B(n_1126),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1264),
.A2(n_1220),
.B(n_1150),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1257),
.A2(n_1080),
.B1(n_1158),
.B2(n_1151),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1240),
.A2(n_1220),
.B(n_1177),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1257),
.A2(n_1080),
.B1(n_1197),
.B2(n_1127),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1237),
.B(n_1127),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1291),
.B(n_1127),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_L g1473 ( 
.A(n_1241),
.B(n_1211),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1284),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1227),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1264),
.A2(n_541),
.B(n_538),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1295),
.B(n_1212),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1383),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1383),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1267),
.A2(n_1177),
.B(n_1197),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1241),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1233),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1289),
.A2(n_545),
.B(n_541),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1246),
.B(n_1120),
.Y(n_1484)
);

BUFx12f_ASAP7_75t_L g1485 ( 
.A(n_1290),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1249),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1260),
.B(n_1029),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1271),
.A2(n_549),
.B(n_545),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1266),
.Y(n_1489)
);

OAI222xp33_ASAP7_75t_L g1490 ( 
.A1(n_1368),
.A2(n_428),
.B1(n_390),
.B2(n_394),
.C1(n_399),
.C2(n_400),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1383),
.B(n_1122),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1383),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1246),
.B(n_1120),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1251),
.Y(n_1494)
);

BUFx4f_ASAP7_75t_L g1495 ( 
.A(n_1284),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1271),
.A2(n_553),
.B(n_549),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1319),
.A2(n_1193),
.B1(n_1129),
.B2(n_1057),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1284),
.B(n_1120),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1284),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1253),
.A2(n_554),
.B(n_553),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1258),
.A2(n_1214),
.B(n_1211),
.Y(n_1501)
);

INVx6_ASAP7_75t_L g1502 ( 
.A(n_1333),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1262),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1352),
.B(n_1057),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1245),
.A2(n_1177),
.B(n_1197),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1353),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1288),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1322),
.B(n_1287),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1299),
.Y(n_1509)
);

AOI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1315),
.A2(n_1154),
.B(n_1165),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1313),
.A2(n_1154),
.B(n_1165),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1253),
.A2(n_554),
.B(n_380),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1296),
.A2(n_1129),
.B1(n_1097),
.B2(n_382),
.C(n_383),
.Y(n_1513)
);

INVx8_ASAP7_75t_L g1514 ( 
.A(n_1239),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1381),
.A2(n_382),
.B(n_375),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1321),
.Y(n_1516)
);

A2O1A1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1320),
.A2(n_1165),
.B(n_1154),
.C(n_1206),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_SL g1518 ( 
.A(n_1361),
.B(n_1181),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1302),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1296),
.A2(n_375),
.B(n_446),
.C(n_447),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1333),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1345),
.A2(n_393),
.B(n_392),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1309),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1318),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1335),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1345),
.A2(n_1348),
.B(n_1292),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1343),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1242),
.A2(n_1111),
.B1(n_1138),
.B2(n_1029),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1348),
.A2(n_397),
.B(n_393),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1362),
.B(n_1211),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1358),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1302),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1270),
.A2(n_1352),
.B1(n_1363),
.B2(n_1223),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1362),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1289),
.A2(n_1292),
.B(n_1308),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1290),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1346),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1308),
.A2(n_417),
.B(n_397),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1276),
.B(n_1181),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1350),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1385),
.A2(n_1197),
.B1(n_1187),
.B2(n_1214),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1366),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1350),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1350),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1285),
.B(n_1181),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1282),
.Y(n_1546)
);

AO31x2_ASAP7_75t_L g1547 ( 
.A1(n_1325),
.A2(n_1214),
.A3(n_458),
.B(n_455),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1239),
.Y(n_1548)
);

NAND2x1p5_ASAP7_75t_L g1549 ( 
.A(n_1321),
.B(n_1181),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1328),
.A2(n_1111),
.B(n_420),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1387),
.B(n_1199),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1316),
.A2(n_420),
.B(n_417),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1316),
.A2(n_458),
.B(n_455),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1346),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1293),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1254),
.A2(n_1206),
.B(n_1203),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1274),
.A2(n_437),
.B(n_401),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1346),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1282),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1331),
.A2(n_1274),
.B(n_1297),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1307),
.B(n_1199),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1366),
.Y(n_1562)
);

AO21x1_ASAP7_75t_L g1563 ( 
.A1(n_1245),
.A2(n_437),
.B(n_1197),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1293),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1374),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1243),
.B(n_1317),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1347),
.A2(n_1206),
.B(n_1203),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1387),
.B(n_1199),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1293),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1282),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1278),
.A2(n_1279),
.B(n_1342),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1417),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1388),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1413),
.A2(n_1187),
.B1(n_454),
.B2(n_425),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1498),
.B(n_1286),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1389),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1475),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1498),
.B(n_1334),
.Y(n_1578)
);

INVx4_ASAP7_75t_SL g1579 ( 
.A(n_1548),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1413),
.A2(n_421),
.B1(n_444),
.B2(n_450),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1456),
.B(n_1293),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1392),
.B(n_1422),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1418),
.A2(n_418),
.B1(n_439),
.B2(n_434),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1475),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1513),
.A2(n_1374),
.B1(n_1281),
.B2(n_1338),
.Y(n_1585)
);

OAI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1520),
.A2(n_403),
.B(n_440),
.C(n_427),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1482),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1395),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1395),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1391),
.A2(n_414),
.B1(n_426),
.B2(n_423),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1482),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1392),
.B(n_1387),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1486),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1501),
.A2(n_1303),
.B(n_1355),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1408),
.A2(n_1468),
.B1(n_1508),
.B2(n_1453),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1464),
.A2(n_410),
.B1(n_416),
.B2(n_422),
.C1(n_1192),
.C2(n_443),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1423),
.B(n_1387),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1404),
.A2(n_1259),
.B1(n_1384),
.B2(n_1382),
.Y(n_1598)
);

INVx8_ASAP7_75t_L g1599 ( 
.A(n_1514),
.Y(n_1599)
);

BUFx8_ASAP7_75t_SL g1600 ( 
.A(n_1485),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1422),
.B(n_1371),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1398),
.B(n_1376),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1486),
.Y(n_1603)
);

INVx6_ASAP7_75t_L g1604 ( 
.A(n_1502),
.Y(n_1604)
);

CKINVDCx6p67_ASAP7_75t_R g1605 ( 
.A(n_1485),
.Y(n_1605)
);

OAI211xp5_ASAP7_75t_L g1606 ( 
.A1(n_1468),
.A2(n_1386),
.B(n_1337),
.C(n_1199),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1535),
.A2(n_1314),
.B(n_1324),
.Y(n_1607)
);

NAND2x1_ASAP7_75t_L g1608 ( 
.A(n_1530),
.B(n_1239),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1424),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1417),
.B(n_1243),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1416),
.A2(n_1303),
.B(n_1379),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1388),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1495),
.Y(n_1613)
);

CKINVDCx11_ASAP7_75t_R g1614 ( 
.A(n_1536),
.Y(n_1614)
);

OR2x6_ASAP7_75t_SL g1615 ( 
.A(n_1415),
.B(n_1293),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1495),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1472),
.B(n_1243),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1424),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1512),
.A2(n_1306),
.B(n_1312),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1524),
.Y(n_1620)
);

CKINVDCx8_ASAP7_75t_R g1621 ( 
.A(n_1415),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1470),
.A2(n_1259),
.B1(n_1206),
.B2(n_1203),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1550),
.A2(n_303),
.B1(n_370),
.B2(n_1203),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1477),
.B(n_1243),
.Y(n_1624)
);

BUFx8_ASAP7_75t_L g1625 ( 
.A(n_1536),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1550),
.A2(n_303),
.B1(n_370),
.B2(n_1239),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1406),
.B(n_303),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1537),
.A2(n_1293),
.B1(n_1239),
.B2(n_370),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1477),
.B(n_1365),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1432),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1556),
.A2(n_1294),
.B(n_1268),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1550),
.A2(n_370),
.B1(n_303),
.B2(n_1344),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1406),
.B(n_303),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1389),
.B(n_303),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1470),
.A2(n_370),
.B1(n_1365),
.B2(n_673),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1432),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1461),
.B(n_370),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1445),
.Y(n_1638)
);

OAI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1541),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1437),
.B(n_370),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1524),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1517),
.A2(n_1339),
.B(n_1356),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1537),
.A2(n_370),
.B1(n_7),
.B2(n_9),
.Y(n_1643)
);

NAND2x1_ASAP7_75t_L g1644 ( 
.A(n_1530),
.B(n_1372),
.Y(n_1644)
);

NAND2xp33_ASAP7_75t_R g1645 ( 
.A(n_1494),
.B(n_123),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1419),
.A2(n_673),
.B1(n_10),
.B2(n_11),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1518),
.A2(n_1373),
.B(n_1360),
.Y(n_1647)
);

OAI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1541),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_15),
.Y(n_1648)
);

OR2x6_ASAP7_75t_L g1649 ( 
.A(n_1514),
.B(n_126),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1514),
.B(n_135),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1525),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1533),
.A2(n_804),
.B1(n_762),
.B2(n_20),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1471),
.B(n_15),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1409),
.B(n_773),
.Y(n_1654)
);

NAND2xp33_ASAP7_75t_L g1655 ( 
.A(n_1528),
.B(n_762),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1494),
.B(n_16),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1393),
.B(n_16),
.Y(n_1657)
);

BUFx2_ASAP7_75t_SL g1658 ( 
.A(n_1444),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_SL g1659 ( 
.A(n_1554),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1533),
.A2(n_804),
.B1(n_22),
.B2(n_25),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1487),
.A2(n_21),
.B1(n_26),
.B2(n_29),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1498),
.B(n_136),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1532),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1445),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1504),
.A2(n_1563),
.B1(n_1466),
.B2(n_1558),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1563),
.A2(n_1554),
.B1(n_1558),
.B2(n_1497),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1514),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1439),
.B(n_33),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1518),
.A2(n_804),
.B(n_811),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1414),
.A2(n_811),
.B1(n_773),
.B2(n_36),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1525),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1414),
.A2(n_811),
.B1(n_35),
.B2(n_37),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1457),
.B(n_34),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1458),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1489),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1489),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1527),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1514),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1527),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1458),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1463),
.B(n_53),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1530),
.B(n_233),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1430),
.A2(n_54),
.B(n_55),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1519),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1452),
.A2(n_811),
.B(n_59),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1428),
.B(n_225),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1433),
.A2(n_1565),
.B1(n_1444),
.B2(n_1548),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_L g1688 ( 
.A(n_1444),
.B(n_56),
.Y(n_1688)
);

CKINVDCx6p67_ASAP7_75t_R g1689 ( 
.A(n_1562),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1531),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1506),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1444),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1507),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1531),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1394),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1532),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1507),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1428),
.B(n_1448),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1474),
.Y(n_1699)
);

INVx6_ASAP7_75t_L g1700 ( 
.A(n_1502),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1509),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1539),
.B(n_64),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1448),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1509),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1428),
.A2(n_1545),
.B1(n_1539),
.B2(n_1480),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1530),
.B(n_140),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1523),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1396),
.A2(n_146),
.B(n_219),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1562),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1545),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1438),
.A2(n_79),
.B(n_81),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1484),
.B(n_1493),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_SL g1713 ( 
.A(n_1444),
.B(n_157),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1484),
.A2(n_82),
.B1(n_87),
.B2(n_89),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1523),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1394),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1399),
.Y(n_1717)
);

NAND2xp33_ASAP7_75t_L g1718 ( 
.A(n_1444),
.B(n_82),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_R g1719 ( 
.A(n_1447),
.B(n_223),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1566),
.A2(n_87),
.B1(n_90),
.B2(n_93),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1490),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.C(n_101),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1566),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_SL g1723 ( 
.A1(n_1546),
.A2(n_103),
.B(n_106),
.C(n_109),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1400),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1534),
.Y(n_1725)
);

OR2x6_ASAP7_75t_L g1726 ( 
.A(n_1530),
.B(n_182),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1410),
.A2(n_109),
.B1(n_110),
.B2(n_138),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1400),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1401),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1396),
.A2(n_110),
.B1(n_217),
.B2(n_144),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1505),
.B(n_139),
.C(n_150),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1410),
.A2(n_169),
.B1(n_171),
.B2(n_175),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1401),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1493),
.B(n_177),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1412),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1499),
.Y(n_1736)
);

OAI211xp5_ASAP7_75t_L g1737 ( 
.A1(n_1469),
.A2(n_179),
.B(n_188),
.C(n_190),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1412),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1429),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1396),
.A2(n_216),
.B1(n_195),
.B2(n_203),
.Y(n_1740)
);

NAND3x1_ASAP7_75t_L g1741 ( 
.A(n_1551),
.B(n_206),
.C(n_207),
.Y(n_1741)
);

CKINVDCx16_ASAP7_75t_R g1742 ( 
.A(n_1411),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1462),
.B(n_209),
.Y(n_1743)
);

INVx6_ASAP7_75t_L g1744 ( 
.A(n_1502),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1551),
.A2(n_1568),
.B1(n_1511),
.B2(n_1473),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1462),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_SL g1747 ( 
.A(n_1561),
.B(n_1481),
.C(n_1435),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1546),
.A2(n_1570),
.B1(n_1559),
.B2(n_1455),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1465),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1559),
.A2(n_1570),
.B1(n_1455),
.B2(n_1568),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1465),
.Y(n_1751)
);

INVx4_ASAP7_75t_SL g1752 ( 
.A(n_1548),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1481),
.B(n_1407),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1455),
.A2(n_1511),
.B1(n_1451),
.B2(n_1426),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1511),
.A2(n_1451),
.B1(n_1426),
.B2(n_1454),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1502),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1411),
.B(n_1443),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1547),
.Y(n_1758)
);

BUFx12f_ASAP7_75t_L g1759 ( 
.A(n_1521),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1451),
.A2(n_1426),
.B1(n_1454),
.B2(n_1442),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1503),
.B(n_1443),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1547),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1451),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1548),
.B(n_1569),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1543),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1450),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1454),
.A2(n_1446),
.B1(n_1442),
.B2(n_1544),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1548),
.A2(n_1534),
.B1(n_1495),
.B2(n_1521),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1542),
.B(n_1521),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1577),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1583),
.A2(n_1473),
.B1(n_1521),
.B2(n_1405),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1584),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1721),
.A2(n_1454),
.B1(n_1446),
.B2(n_1442),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1711),
.A2(n_1571),
.B(n_1390),
.Y(n_1774)
);

AOI222xp33_ASAP7_75t_L g1775 ( 
.A1(n_1646),
.A2(n_1540),
.B1(n_1534),
.B2(n_1542),
.C1(n_1516),
.C2(n_1543),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1582),
.B(n_1425),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1596),
.A2(n_1442),
.B1(n_1446),
.B2(n_1534),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1583),
.A2(n_1491),
.B1(n_1436),
.B2(n_1405),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1646),
.A2(n_1405),
.B(n_1436),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1661),
.A2(n_1446),
.B1(n_1534),
.B2(n_1557),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1587),
.Y(n_1781)
);

OAI211xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1574),
.A2(n_1540),
.B(n_1544),
.C(n_1516),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1661),
.A2(n_1722),
.B1(n_1720),
.B2(n_1685),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1699),
.Y(n_1785)
);

OAI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1645),
.A2(n_1478),
.B1(n_1492),
.B2(n_1447),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1595),
.B(n_1425),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1668),
.B(n_1516),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1639),
.A2(n_1555),
.B1(n_1564),
.B2(n_1479),
.C(n_1492),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1574),
.A2(n_1449),
.B1(n_1427),
.B2(n_1549),
.C(n_1436),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1634),
.B(n_1547),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1712),
.B(n_1547),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1698),
.B(n_1447),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1696),
.A2(n_1557),
.B(n_1449),
.C(n_1427),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1720),
.A2(n_1557),
.B1(n_1390),
.B2(n_1552),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1645),
.A2(n_1478),
.B1(n_1479),
.B2(n_1492),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1591),
.Y(n_1797)
);

OAI222xp33_ASAP7_75t_L g1798 ( 
.A1(n_1643),
.A2(n_1459),
.B1(n_1549),
.B2(n_1491),
.C1(n_1478),
.C2(n_1479),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1722),
.A2(n_1557),
.B1(n_1552),
.B2(n_1397),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1597),
.B(n_1425),
.Y(n_1800)
);

OAI211xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1580),
.A2(n_1564),
.B(n_1555),
.C(n_1425),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1639),
.A2(n_1648),
.B1(n_1683),
.B2(n_1580),
.C(n_1675),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1675),
.A2(n_1552),
.B1(n_1397),
.B2(n_1467),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1593),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1676),
.A2(n_1450),
.B1(n_1549),
.B2(n_1569),
.C(n_1491),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1603),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1627),
.B(n_1450),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1676),
.A2(n_1552),
.B1(n_1467),
.B2(n_1571),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1697),
.A2(n_1460),
.B1(n_1553),
.B2(n_1538),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1697),
.A2(n_1460),
.B1(n_1553),
.B2(n_1538),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1707),
.A2(n_1483),
.B1(n_1476),
.B2(n_1515),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1595),
.A2(n_1569),
.B1(n_1459),
.B2(n_1510),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1613),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1688),
.A2(n_1567),
.B1(n_1515),
.B2(n_1450),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1707),
.A2(n_1483),
.B1(n_1476),
.B2(n_1496),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1657),
.A2(n_1483),
.B1(n_1500),
.B2(n_1496),
.Y(n_1816)
);

OAI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1590),
.A2(n_1678),
.B1(n_1667),
.B2(n_1718),
.C(n_1730),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_SL g1818 ( 
.A1(n_1730),
.A2(n_1450),
.B(n_1510),
.C(n_1567),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1633),
.B(n_1488),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1760),
.A2(n_1560),
.B(n_1500),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1666),
.A2(n_1483),
.B1(n_1529),
.B2(n_1522),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1703),
.B(n_1560),
.C(n_1421),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1613),
.Y(n_1823)
);

AOI331xp33_ASAP7_75t_L g1824 ( 
.A1(n_1590),
.A2(n_1421),
.A3(n_1440),
.B1(n_1420),
.B2(n_1441),
.B3(n_1434),
.C1(n_1402),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1637),
.B(n_1402),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1620),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1695),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1714),
.A2(n_1403),
.B1(n_1526),
.B2(n_1434),
.C(n_1441),
.Y(n_1828)
);

NAND2xp33_ASAP7_75t_R g1829 ( 
.A(n_1682),
.B(n_1403),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1660),
.A2(n_1431),
.B1(n_1526),
.B2(n_1723),
.C(n_1727),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1723),
.A2(n_1431),
.B1(n_1710),
.B2(n_1652),
.C(n_1665),
.Y(n_1831)
);

AO21x1_ASAP7_75t_L g1832 ( 
.A1(n_1719),
.A2(n_1581),
.B(n_1654),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1665),
.A2(n_1586),
.B1(n_1740),
.B2(n_1653),
.C(n_1640),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1695),
.Y(n_1834)
);

AOI222xp33_ASAP7_75t_L g1835 ( 
.A1(n_1740),
.A2(n_1656),
.B1(n_1655),
.B2(n_1666),
.C1(n_1606),
.C2(n_1702),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1613),
.Y(n_1836)
);

BUFx8_ASAP7_75t_SL g1837 ( 
.A(n_1600),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1732),
.A2(n_1737),
.B1(n_1731),
.B2(n_1682),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1576),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1611),
.A2(n_1642),
.B(n_1594),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1601),
.B(n_1602),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1672),
.A2(n_1682),
.B1(n_1726),
.B2(n_1706),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1708),
.A2(n_1598),
.B1(n_1691),
.B2(n_1623),
.C(n_1635),
.Y(n_1843)
);

OA21x2_ASAP7_75t_L g1844 ( 
.A1(n_1760),
.A2(n_1767),
.B(n_1755),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1641),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1759),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1585),
.A2(n_1719),
.B1(n_1741),
.B2(n_1605),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1613),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1706),
.A2(n_1726),
.B1(n_1684),
.B2(n_1581),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1572),
.B(n_1673),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1654),
.A2(n_1747),
.B(n_1632),
.Y(n_1851)
);

OAI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1670),
.A2(n_1635),
.B1(n_1626),
.B2(n_1632),
.C(n_1623),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1576),
.Y(n_1853)
);

AO22x2_ASAP7_75t_L g1854 ( 
.A1(n_1758),
.A2(n_1762),
.B1(n_1624),
.B2(n_1610),
.Y(n_1854)
);

AOI222xp33_ASAP7_75t_L g1855 ( 
.A1(n_1659),
.A2(n_1681),
.B1(n_1622),
.B2(n_1614),
.C1(n_1625),
.C2(n_1626),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1651),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1706),
.A2(n_1726),
.B1(n_1649),
.B2(n_1650),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1622),
.A2(n_1734),
.B(n_1629),
.C(n_1686),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1572),
.B(n_1698),
.Y(n_1859)
);

OAI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1687),
.A2(n_1621),
.B(n_1617),
.C(n_1705),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1649),
.A2(n_1650),
.B1(n_1659),
.B2(n_1663),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1649),
.A2(n_1650),
.B1(n_1625),
.B2(n_1662),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1647),
.A2(n_1631),
.B(n_1608),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1578),
.B(n_1769),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1701),
.B(n_1704),
.Y(n_1865)
);

AOI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1662),
.A2(n_1686),
.B1(n_1766),
.B2(n_1713),
.C1(n_1715),
.C2(n_1677),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1578),
.A2(n_1693),
.B1(n_1690),
.B2(n_1671),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1607),
.A2(n_1644),
.B(n_1767),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1679),
.A2(n_1694),
.B1(n_1766),
.B2(n_1575),
.Y(n_1869)
);

OA21x2_ASAP7_75t_L g1870 ( 
.A1(n_1755),
.A2(n_1754),
.B(n_1748),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_SL g1871 ( 
.A1(n_1658),
.A2(n_1599),
.B1(n_1736),
.B2(n_1709),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1716),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1615),
.A2(n_1768),
.B1(n_1742),
.B2(n_1689),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1717),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1745),
.A2(n_1628),
.B1(n_1573),
.B2(n_1612),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1757),
.B(n_1756),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1575),
.A2(n_1728),
.B1(n_1746),
.B2(n_1729),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1724),
.A2(n_1735),
.B1(n_1738),
.B2(n_1739),
.Y(n_1878)
);

OAI211xp5_ASAP7_75t_L g1879 ( 
.A1(n_1753),
.A2(n_1750),
.B(n_1761),
.C(n_1754),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1604),
.A2(n_1744),
.B1(n_1700),
.B2(n_1616),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1588),
.B(n_1636),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1733),
.B(n_1749),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1733),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1750),
.A2(n_1748),
.B1(n_1749),
.B2(n_1751),
.C(n_1763),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1674),
.B(n_1751),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1604),
.A2(n_1744),
.B1(n_1700),
.B2(n_1616),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1599),
.A2(n_1616),
.B1(n_1744),
.B2(n_1604),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1616),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1743),
.A2(n_1664),
.B1(n_1589),
.B2(n_1638),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1763),
.A2(n_1664),
.B1(n_1680),
.B2(n_1609),
.C(n_1618),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1609),
.B(n_1630),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1618),
.A2(n_1680),
.B1(n_1630),
.B2(n_1638),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1700),
.A2(n_1599),
.B1(n_1725),
.B2(n_1692),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1579),
.B(n_1752),
.Y(n_1894)
);

NAND3xp33_ASAP7_75t_L g1895 ( 
.A(n_1692),
.B(n_1764),
.C(n_1619),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1579),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1579),
.B(n_1752),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1764),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1752),
.B(n_1764),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1669),
.A2(n_1027),
.B(n_1611),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1619),
.B(n_1582),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1619),
.A2(n_1721),
.B1(n_1596),
.B2(n_1711),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1699),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1709),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1577),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1582),
.B(n_1413),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_SL g1907 ( 
.A1(n_1688),
.A2(n_957),
.B1(n_1718),
.B2(n_1732),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_1759),
.Y(n_1908)
);

OAI211xp5_ASAP7_75t_SL g1909 ( 
.A1(n_1596),
.A2(n_1090),
.B(n_1513),
.C(n_1583),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1582),
.B(n_1413),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1698),
.B(n_1579),
.Y(n_1911)
);

NAND2x1_ASAP7_75t_L g1912 ( 
.A(n_1692),
.B(n_1764),
.Y(n_1912)
);

OAI211xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1596),
.A2(n_1090),
.B(n_1513),
.C(n_1583),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1582),
.B(n_1413),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1684),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1582),
.B(n_1413),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1572),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1583),
.A2(n_1163),
.B1(n_1189),
.B2(n_1418),
.Y(n_1921)
);

OAI21x1_ASAP7_75t_SL g1922 ( 
.A1(n_1711),
.A2(n_1685),
.B(n_1487),
.Y(n_1922)
);

AO31x2_ASAP7_75t_L g1923 ( 
.A1(n_1758),
.A2(n_1762),
.A3(n_1546),
.B(n_1570),
.Y(n_1923)
);

AO31x2_ASAP7_75t_L g1924 ( 
.A1(n_1758),
.A2(n_1762),
.A3(n_1546),
.B(n_1570),
.Y(n_1924)
);

AOI222xp33_ASAP7_75t_L g1925 ( 
.A1(n_1721),
.A2(n_1646),
.B1(n_1711),
.B2(n_1661),
.C1(n_937),
.C2(n_1583),
.Y(n_1925)
);

OAI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1645),
.A2(n_957),
.B1(n_1189),
.B2(n_1163),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1582),
.B(n_1413),
.Y(n_1927)
);

OAI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1645),
.A2(n_957),
.B1(n_1189),
.B2(n_1163),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1583),
.A2(n_1163),
.B1(n_1189),
.B2(n_1418),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1582),
.B(n_1413),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1582),
.B(n_1572),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1721),
.A2(n_1520),
.B1(n_1639),
.B2(n_922),
.C(n_694),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1684),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1583),
.A2(n_922),
.B1(n_1090),
.B2(n_957),
.C(n_973),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1721),
.A2(n_1520),
.B1(n_1639),
.B2(n_922),
.C(n_694),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1940)
);

OAI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1645),
.A2(n_957),
.B1(n_1189),
.B2(n_1163),
.Y(n_1941)
);

AO221x2_ASAP7_75t_L g1942 ( 
.A1(n_1639),
.A2(n_1648),
.B1(n_1727),
.B2(n_1711),
.C(n_1464),
.Y(n_1942)
);

AOI222xp33_ASAP7_75t_L g1943 ( 
.A1(n_1721),
.A2(n_1646),
.B1(n_1711),
.B2(n_1661),
.C1(n_937),
.C2(n_1583),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1582),
.B(n_1572),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1765),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1611),
.A2(n_1027),
.B(n_859),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1721),
.A2(n_1596),
.B1(n_1711),
.B2(n_1661),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1923),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1920),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1933),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1827),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1923),
.Y(n_1952)
);

AO31x2_ASAP7_75t_L g1953 ( 
.A1(n_1812),
.A2(n_1821),
.A3(n_1840),
.B(n_1900),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1944),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1923),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1776),
.B(n_1939),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1923),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1841),
.B(n_1854),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1906),
.B(n_1910),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1800),
.B(n_1783),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1898),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1924),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1834),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1834),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1807),
.B(n_1792),
.Y(n_1965)
);

INVx4_ASAP7_75t_R g1966 ( 
.A(n_1894),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1924),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1870),
.B(n_1791),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1870),
.B(n_1854),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1870),
.B(n_1854),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1844),
.B(n_1770),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1844),
.B(n_1772),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1872),
.B(n_1874),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1924),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1844),
.B(n_1781),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1901),
.B(n_1924),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1883),
.B(n_1895),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1797),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1898),
.Y(n_1979)
);

NAND2xp33_ASAP7_75t_L g1980 ( 
.A(n_1914),
.B(n_1915),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1804),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1806),
.Y(n_1982)
);

NAND4xp25_ASAP7_75t_L g1983 ( 
.A(n_1914),
.B(n_1947),
.C(n_1930),
.D(n_1916),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1917),
.B(n_1919),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1942),
.A2(n_1947),
.B1(n_1936),
.B2(n_1931),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1826),
.B(n_1845),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1856),
.B(n_1905),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1825),
.B(n_1850),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1884),
.B(n_1869),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1787),
.B(n_1859),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1882),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1945),
.B(n_1819),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1865),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1868),
.Y(n_1994)
);

NOR2x1_ASAP7_75t_L g1995 ( 
.A(n_1782),
.B(n_1786),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1891),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1879),
.B(n_1927),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1932),
.B(n_1839),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1878),
.B(n_1877),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1868),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1785),
.B(n_1903),
.Y(n_2001)
);

NOR2x1_ASAP7_75t_SL g2002 ( 
.A(n_1860),
.B(n_1794),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1885),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1918),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1878),
.B(n_1877),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1881),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1864),
.B(n_1876),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1829),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1867),
.B(n_1774),
.Y(n_2009)
);

AOI211xp5_ASAP7_75t_L g2010 ( 
.A1(n_1937),
.A2(n_1909),
.B(n_1913),
.C(n_1928),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1935),
.Y(n_2011)
);

BUFx3_ASAP7_75t_L g2012 ( 
.A(n_1912),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1820),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1892),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1853),
.B(n_1822),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1892),
.B(n_1780),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1780),
.B(n_1788),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1820),
.B(n_1832),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1788),
.B(n_1849),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1890),
.Y(n_2020)
);

BUFx3_ASAP7_75t_L g2021 ( 
.A(n_1911),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1849),
.B(n_1818),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1801),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1818),
.B(n_1851),
.Y(n_2024)
);

INVx2_ASAP7_75t_R g2025 ( 
.A(n_1896),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1828),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1790),
.Y(n_2027)
);

OAI211xp5_ASAP7_75t_L g2028 ( 
.A1(n_1915),
.A2(n_1930),
.B(n_1931),
.C(n_1936),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1889),
.B(n_1773),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1773),
.B(n_1796),
.Y(n_2030)
);

INVxp67_ASAP7_75t_L g2031 ( 
.A(n_1829),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1793),
.B(n_1808),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1863),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1946),
.B(n_1902),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1793),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1808),
.B(n_1799),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1799),
.B(n_1795),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1795),
.B(n_1803),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1803),
.Y(n_2039)
);

AOI31xp33_ASAP7_75t_L g2040 ( 
.A1(n_1907),
.A2(n_1784),
.A3(n_1916),
.B(n_1940),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1922),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1911),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1926),
.B(n_1941),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_1942),
.A2(n_1940),
.B1(n_1784),
.B2(n_1925),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1814),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1899),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1942),
.A2(n_1943),
.B1(n_1938),
.B2(n_1934),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1830),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1809),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1902),
.B(n_1777),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1816),
.A2(n_1810),
.B(n_1809),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1810),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1873),
.B(n_1816),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1980),
.A2(n_1817),
.B1(n_1802),
.B2(n_1838),
.Y(n_2054)
);

AND2x4_ASAP7_75t_SL g2055 ( 
.A(n_1961),
.B(n_1857),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1950),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1983),
.A2(n_1842),
.B1(n_1833),
.B2(n_1857),
.Y(n_2057)
);

OR2x2_ASAP7_75t_L g2058 ( 
.A(n_1958),
.B(n_1875),
.Y(n_2058)
);

BUFx2_ASAP7_75t_L g2059 ( 
.A(n_1977),
.Y(n_2059)
);

OAI33xp33_ASAP7_75t_L g2060 ( 
.A1(n_1983),
.A2(n_2048),
.A3(n_1958),
.B1(n_1997),
.B2(n_2034),
.B3(n_2024),
.Y(n_2060)
);

INVx5_ASAP7_75t_SL g2061 ( 
.A(n_1961),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_1954),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1960),
.B(n_1866),
.Y(n_2063)
);

AO21x2_ASAP7_75t_L g2064 ( 
.A1(n_2034),
.A2(n_1847),
.B(n_1798),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_2012),
.Y(n_2065)
);

AO21x2_ASAP7_75t_L g2066 ( 
.A1(n_1948),
.A2(n_1824),
.B(n_1779),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_2047),
.A2(n_1842),
.B1(n_1862),
.B2(n_1861),
.Y(n_2067)
);

OAI31xp33_ASAP7_75t_L g2068 ( 
.A1(n_2028),
.A2(n_1929),
.A3(n_1921),
.B(n_1777),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2028),
.A2(n_1861),
.B(n_1835),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1960),
.B(n_1855),
.Y(n_2070)
);

OR2x6_ASAP7_75t_L g2071 ( 
.A(n_2008),
.B(n_1897),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1959),
.B(n_1904),
.Y(n_2072)
);

OAI31xp33_ASAP7_75t_SL g2073 ( 
.A1(n_2043),
.A2(n_1831),
.A3(n_1871),
.B(n_1843),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1998),
.B(n_1775),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_2044),
.A2(n_1852),
.B1(n_1862),
.B2(n_1771),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1990),
.B(n_1976),
.Y(n_2076)
);

AO21x2_ASAP7_75t_L g2077 ( 
.A1(n_1948),
.A2(n_1778),
.B(n_1886),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1995),
.B(n_1837),
.Y(n_2078)
);

OAI211xp5_ASAP7_75t_SL g2079 ( 
.A1(n_2010),
.A2(n_1858),
.B(n_1880),
.C(n_1893),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1990),
.B(n_1815),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1978),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1985),
.A2(n_1789),
.B1(n_1805),
.B2(n_1908),
.Y(n_2082)
);

AOI211xp5_ASAP7_75t_L g2083 ( 
.A1(n_2010),
.A2(n_1846),
.B(n_1908),
.C(n_1848),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2035),
.B(n_1893),
.Y(n_2084)
);

OAI332xp33_ASAP7_75t_L g2085 ( 
.A1(n_2048),
.A2(n_1837),
.A3(n_1887),
.B1(n_1811),
.B2(n_1815),
.B3(n_1846),
.C1(n_1823),
.C2(n_1848),
.Y(n_2085)
);

OAI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2024),
.A2(n_1811),
.B(n_1836),
.C(n_1888),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_1976),
.B(n_1888),
.Y(n_2087)
);

CKINVDCx16_ASAP7_75t_R g2088 ( 
.A(n_2021),
.Y(n_2088)
);

INVx1_ASAP7_75t_SL g2089 ( 
.A(n_1998),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1984),
.B(n_1848),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1978),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1951),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_1949),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_2001),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_1971),
.B(n_1972),
.Y(n_2095)
);

OAI31xp33_ASAP7_75t_L g2096 ( 
.A1(n_2050),
.A2(n_1813),
.A3(n_1823),
.B(n_1848),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1965),
.B(n_1813),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2050),
.A2(n_1813),
.B1(n_1823),
.B2(n_1989),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2040),
.A2(n_1813),
.B(n_1823),
.Y(n_2099)
);

AOI221xp5_ASAP7_75t_L g2100 ( 
.A1(n_2040),
.A2(n_2026),
.B1(n_2017),
.B2(n_1989),
.C(n_2027),
.Y(n_2100)
);

OAI31xp33_ASAP7_75t_L g2101 ( 
.A1(n_2023),
.A2(n_2030),
.A3(n_2027),
.B(n_2037),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2017),
.A2(n_2019),
.B1(n_2030),
.B2(n_2041),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_1949),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2019),
.A2(n_2041),
.B1(n_2009),
.B2(n_2045),
.Y(n_2104)
);

NAND2xp33_ASAP7_75t_R g2105 ( 
.A(n_1997),
.B(n_1969),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1981),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1995),
.A2(n_2041),
.B(n_2022),
.Y(n_2107)
);

OAI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2022),
.A2(n_2026),
.B1(n_2027),
.B2(n_2053),
.C(n_2045),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_1979),
.Y(n_2109)
);

OAI31xp33_ASAP7_75t_L g2110 ( 
.A1(n_2023),
.A2(n_2037),
.A3(n_2029),
.B(n_2053),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_SL g2111 ( 
.A1(n_2002),
.A2(n_2036),
.B1(n_2009),
.B2(n_1999),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1971),
.B(n_1972),
.Y(n_2112)
);

AOI33xp33_ASAP7_75t_L g2113 ( 
.A1(n_1969),
.A2(n_1970),
.A3(n_2026),
.B1(n_2020),
.B2(n_2052),
.B3(n_2049),
.Y(n_2113)
);

OAI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2029),
.A2(n_2008),
.B(n_2031),
.C(n_2036),
.Y(n_2114)
);

INVx4_ASAP7_75t_L g2115 ( 
.A(n_2012),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1968),
.B(n_1988),
.Y(n_2116)
);

OA21x2_ASAP7_75t_L g2117 ( 
.A1(n_2013),
.A2(n_1974),
.B(n_1955),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1981),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_1999),
.A2(n_2005),
.B1(n_2020),
.B2(n_2016),
.Y(n_2119)
);

NOR2x1p5_ASAP7_75t_L g2120 ( 
.A(n_2012),
.B(n_2021),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2005),
.A2(n_2046),
.B1(n_2032),
.B2(n_2016),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1963),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_1977),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1963),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_1975),
.B(n_1970),
.Y(n_2125)
);

NAND2xp33_ASAP7_75t_SL g2126 ( 
.A(n_2042),
.B(n_1961),
.Y(n_2126)
);

AND2x6_ASAP7_75t_SL g2127 ( 
.A(n_2007),
.B(n_1956),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1964),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1956),
.B(n_2006),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2006),
.B(n_2003),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1977),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1982),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2003),
.B(n_1991),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_2032),
.A2(n_2052),
.B1(n_2049),
.B2(n_2038),
.Y(n_2134)
);

AOI211xp5_ASAP7_75t_L g2135 ( 
.A1(n_2038),
.A2(n_2031),
.B(n_2015),
.C(n_2039),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2081),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2116),
.B(n_1975),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_2117),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2081),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2076),
.B(n_1993),
.Y(n_2140)
);

HB1xp67_ASAP7_75t_L g2141 ( 
.A(n_2095),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2091),
.Y(n_2142)
);

NAND2x1p5_ASAP7_75t_L g2143 ( 
.A(n_2115),
.B(n_2018),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2125),
.B(n_2018),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_2120),
.B(n_1994),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2091),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2125),
.B(n_2013),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2112),
.B(n_2015),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2120),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2106),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2112),
.B(n_1977),
.Y(n_2151)
);

AOI221xp5_ASAP7_75t_L g2152 ( 
.A1(n_2060),
.A2(n_2039),
.B1(n_2004),
.B2(n_2011),
.C(n_2014),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2106),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2076),
.B(n_1993),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2059),
.B(n_1974),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_2078),
.B(n_2007),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2118),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2059),
.B(n_1962),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2129),
.B(n_1991),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2135),
.B(n_1996),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2117),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_2078),
.B(n_2035),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2118),
.Y(n_2163)
);

OAI33xp33_ASAP7_75t_L g2164 ( 
.A1(n_2067),
.A2(n_1962),
.A3(n_1957),
.B1(n_1955),
.B2(n_1986),
.B3(n_1973),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2123),
.B(n_1957),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2131),
.B(n_1952),
.Y(n_2166)
);

INVx1_ASAP7_75t_SL g2167 ( 
.A(n_2089),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2117),
.B(n_1952),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2135),
.B(n_1996),
.Y(n_2169)
);

NOR3xp33_ASAP7_75t_L g2170 ( 
.A(n_2069),
.B(n_2033),
.C(n_2014),
.Y(n_2170)
);

INVx1_ASAP7_75t_SL g2171 ( 
.A(n_2087),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2132),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2117),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2132),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2133),
.B(n_1992),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2066),
.B(n_1967),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2066),
.B(n_1967),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2130),
.B(n_1992),
.Y(n_2178)
);

NAND2x1_ASAP7_75t_L g2179 ( 
.A(n_2115),
.B(n_1966),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2092),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2066),
.B(n_2000),
.Y(n_2181)
);

INVxp67_ASAP7_75t_L g2182 ( 
.A(n_2107),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2122),
.B(n_2051),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2056),
.B(n_1953),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_2071),
.B(n_1994),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2124),
.B(n_2051),
.Y(n_2186)
);

AND2x2_ASAP7_75t_SL g2187 ( 
.A(n_2113),
.B(n_2051),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2071),
.B(n_1994),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2128),
.B(n_2097),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2093),
.B(n_1987),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_2167),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2138),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2144),
.B(n_2087),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2144),
.B(n_2080),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_2167),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2136),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2184),
.B(n_2080),
.Y(n_2197)
);

OAI21xp33_ASAP7_75t_L g2198 ( 
.A1(n_2170),
.A2(n_2073),
.B(n_2182),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2182),
.B(n_2063),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2184),
.B(n_2103),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2136),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_2149),
.B(n_2071),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2139),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2160),
.B(n_2063),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2139),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2160),
.B(n_2119),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2138),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2138),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2138),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_2169),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2161),
.Y(n_2211)
);

OAI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_2187),
.A2(n_2057),
.B1(n_2054),
.B2(n_2111),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2142),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2151),
.B(n_2071),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2142),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2148),
.B(n_2062),
.Y(n_2216)
);

OR2x6_ASAP7_75t_L g2217 ( 
.A(n_2179),
.B(n_2071),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2161),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2148),
.B(n_2169),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2141),
.B(n_2058),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2146),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2141),
.B(n_2058),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2155),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2146),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2155),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2150),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2151),
.B(n_2088),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2150),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2151),
.B(n_2088),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_2156),
.B(n_2094),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_2190),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2153),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2190),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2153),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2162),
.B(n_2072),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2161),
.Y(n_2236)
);

INVxp67_ASAP7_75t_SL g2237 ( 
.A(n_2143),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2149),
.B(n_2097),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2152),
.B(n_2119),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2149),
.B(n_2137),
.Y(n_2240)
);

OR2x6_ASAP7_75t_L g2241 ( 
.A(n_2179),
.B(n_2143),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2171),
.B(n_2121),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2171),
.B(n_2134),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2157),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2157),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2163),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2152),
.B(n_2110),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2211),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2210),
.B(n_2110),
.Y(n_2249)
);

AND4x1_ASAP7_75t_L g2250 ( 
.A(n_2198),
.B(n_2083),
.C(n_2068),
.D(n_2101),
.Y(n_2250)
);

INVxp67_ASAP7_75t_SL g2251 ( 
.A(n_2220),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_2220),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2214),
.B(n_2145),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2196),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2222),
.Y(n_2255)
);

INVxp33_ASAP7_75t_L g2256 ( 
.A(n_2230),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_2206),
.B(n_2108),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2199),
.Y(n_2258)
);

INVx2_ASAP7_75t_SL g2259 ( 
.A(n_2240),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2196),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2228),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2228),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_2219),
.B(n_2140),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2247),
.B(n_2170),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2222),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2214),
.B(n_2145),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2204),
.B(n_2101),
.Y(n_2267)
);

OAI222xp33_ASAP7_75t_L g2268 ( 
.A1(n_2239),
.A2(n_2102),
.B1(n_2104),
.B2(n_2098),
.C1(n_2075),
.C2(n_2070),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2240),
.B(n_2145),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2202),
.B(n_2145),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2211),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2235),
.B(n_2159),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2218),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_2219),
.B(n_2197),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2233),
.B(n_2187),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2191),
.B(n_2187),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2202),
.B(n_2217),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_SL g2278 ( 
.A(n_2212),
.Y(n_2278)
);

NOR3xp33_ASAP7_75t_L g2279 ( 
.A(n_2195),
.B(n_2100),
.C(n_2079),
.Y(n_2279)
);

NOR2x1_ASAP7_75t_L g2280 ( 
.A(n_2241),
.B(n_2217),
.Y(n_2280)
);

AOI221x1_ASAP7_75t_SL g2281 ( 
.A1(n_2202),
.A2(n_2083),
.B1(n_2140),
.B2(n_2154),
.C(n_2159),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2217),
.B(n_2145),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2231),
.B(n_2154),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2218),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2232),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2217),
.B(n_2137),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_2241),
.Y(n_2287)
);

OR2x2_ASAP7_75t_L g2288 ( 
.A(n_2197),
.B(n_2194),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2232),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2216),
.B(n_2137),
.Y(n_2290)
);

NAND2xp33_ASAP7_75t_R g2291 ( 
.A(n_2243),
.B(n_2099),
.Y(n_2291)
);

NAND2x1p5_ASAP7_75t_L g2292 ( 
.A(n_2227),
.B(n_2115),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2243),
.B(n_2147),
.Y(n_2293)
);

AOI221xp5_ASAP7_75t_L g2294 ( 
.A1(n_2237),
.A2(n_2164),
.B1(n_2181),
.B2(n_2177),
.C(n_2176),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2194),
.B(n_2183),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2200),
.B(n_2183),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_2241),
.Y(n_2297)
);

NAND2xp33_ASAP7_75t_SL g2298 ( 
.A(n_2227),
.B(n_2105),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2236),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2234),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2229),
.B(n_2147),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2242),
.Y(n_2302)
);

OAI21xp33_ASAP7_75t_L g2303 ( 
.A1(n_2264),
.A2(n_2242),
.B(n_2082),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_2278),
.Y(n_2304)
);

OAI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2268),
.A2(n_2068),
.B(n_2181),
.Y(n_2305)
);

NAND3xp33_ASAP7_75t_L g2306 ( 
.A(n_2250),
.B(n_2176),
.C(n_2177),
.Y(n_2306)
);

NAND2x1p5_ASAP7_75t_L g2307 ( 
.A(n_2280),
.B(n_2176),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_SL g2308 ( 
.A1(n_2257),
.A2(n_2002),
.B1(n_2064),
.B2(n_2114),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2254),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2272),
.B(n_2238),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2254),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_2256),
.B(n_2267),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2280),
.B(n_2241),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2260),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2260),
.Y(n_2315)
);

AOI221xp5_ASAP7_75t_L g2316 ( 
.A1(n_2281),
.A2(n_2164),
.B1(n_2181),
.B2(n_2177),
.C(n_2085),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2259),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2261),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2259),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2258),
.B(n_2216),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2281),
.B(n_2302),
.Y(n_2321)
);

O2A1O1Ixp5_ASAP7_75t_L g2322 ( 
.A1(n_2298),
.A2(n_2126),
.B(n_2086),
.C(n_2229),
.Y(n_2322)
);

NAND2xp33_ASAP7_75t_L g2323 ( 
.A(n_2279),
.B(n_2070),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2250),
.B(n_2238),
.Y(n_2324)
);

AOI31xp33_ASAP7_75t_L g2325 ( 
.A1(n_2291),
.A2(n_2143),
.A3(n_2098),
.B(n_2074),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2248),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2292),
.B(n_2223),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2261),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2262),
.Y(n_2329)
);

OAI21xp33_ASAP7_75t_L g2330 ( 
.A1(n_2249),
.A2(n_2055),
.B(n_2200),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2248),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2249),
.A2(n_2297),
.B1(n_2294),
.B2(n_2277),
.Y(n_2332)
);

INVx1_ASAP7_75t_SL g2333 ( 
.A(n_2252),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2276),
.A2(n_2085),
.B(n_2064),
.Y(n_2334)
);

AOI221xp5_ASAP7_75t_L g2335 ( 
.A1(n_2275),
.A2(n_2225),
.B1(n_2224),
.B2(n_2244),
.C(n_2205),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2262),
.Y(n_2336)
);

INVx2_ASAP7_75t_SL g2337 ( 
.A(n_2292),
.Y(n_2337)
);

INVxp33_ASAP7_75t_L g2338 ( 
.A(n_2292),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2263),
.B(n_2175),
.Y(n_2339)
);

INVxp33_ASAP7_75t_L g2340 ( 
.A(n_2277),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2275),
.A2(n_2143),
.B1(n_2055),
.B2(n_2193),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2251),
.A2(n_2064),
.B(n_2090),
.Y(n_2342)
);

AOI22xp33_ASAP7_75t_L g2343 ( 
.A1(n_2286),
.A2(n_2282),
.B1(n_2287),
.B2(n_2293),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2248),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2309),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_SL g2346 ( 
.A1(n_2305),
.A2(n_2287),
.B1(n_2282),
.B2(n_2255),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2309),
.Y(n_2347)
);

AOI222xp33_ASAP7_75t_L g2348 ( 
.A1(n_2323),
.A2(n_2265),
.B1(n_2293),
.B2(n_2283),
.C1(n_2286),
.C2(n_2290),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2340),
.B(n_2253),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2311),
.Y(n_2350)
);

AOI311xp33_ASAP7_75t_L g2351 ( 
.A1(n_2316),
.A2(n_2285),
.A3(n_2300),
.B(n_2289),
.C(n_2245),
.Y(n_2351)
);

INVx1_ASAP7_75t_SL g2352 ( 
.A(n_2304),
.Y(n_2352)
);

AOI222xp33_ASAP7_75t_L g2353 ( 
.A1(n_2323),
.A2(n_2287),
.B1(n_2301),
.B2(n_2270),
.C1(n_2168),
.C2(n_2269),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2332),
.A2(n_2287),
.B1(n_2270),
.B2(n_2269),
.Y(n_2354)
);

NAND2x1_ASAP7_75t_SL g2355 ( 
.A(n_2313),
.B(n_2327),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2308),
.B(n_2322),
.Y(n_2356)
);

NAND4xp75_ASAP7_75t_L g2357 ( 
.A(n_2313),
.B(n_2096),
.C(n_2253),
.D(n_2266),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2307),
.Y(n_2358)
);

AOI31xp33_ASAP7_75t_L g2359 ( 
.A1(n_2324),
.A2(n_2274),
.A3(n_2288),
.B(n_2263),
.Y(n_2359)
);

OAI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2306),
.A2(n_2274),
.B1(n_2288),
.B2(n_2295),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2333),
.B(n_2310),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2311),
.Y(n_2362)
);

AOI222xp33_ASAP7_75t_L g2363 ( 
.A1(n_2303),
.A2(n_2301),
.B1(n_2168),
.B2(n_2289),
.C1(n_2285),
.C2(n_2300),
.Y(n_2363)
);

OAI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2334),
.A2(n_2096),
.B(n_2168),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2312),
.B(n_2266),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2321),
.B(n_2295),
.Y(n_2366)
);

AOI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2330),
.A2(n_2185),
.B1(n_2188),
.B2(n_2084),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2314),
.Y(n_2368)
);

AOI222xp33_ASAP7_75t_L g2369 ( 
.A1(n_2335),
.A2(n_2186),
.B1(n_2183),
.B2(n_2166),
.C1(n_2158),
.C2(n_2155),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2320),
.B(n_2193),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2314),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2339),
.B(n_2234),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2318),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_SL g2374 ( 
.A(n_2307),
.B(n_2065),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2343),
.A2(n_2185),
.B1(n_2188),
.B2(n_2084),
.Y(n_2375)
);

NOR3xp33_ASAP7_75t_SL g2376 ( 
.A(n_2356),
.B(n_2341),
.C(n_2342),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2345),
.Y(n_2377)
);

AOI21xp33_ASAP7_75t_L g2378 ( 
.A1(n_2359),
.A2(n_2338),
.B(n_2337),
.Y(n_2378)
);

OR3x1_ASAP7_75t_L g2379 ( 
.A(n_2355),
.B(n_2315),
.C(n_2329),
.Y(n_2379)
);

NOR3xp33_ASAP7_75t_SL g2380 ( 
.A(n_2366),
.B(n_2328),
.C(n_2318),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2347),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2361),
.B(n_2317),
.Y(n_2382)
);

INVx1_ASAP7_75t_SL g2383 ( 
.A(n_2352),
.Y(n_2383)
);

AOI21xp33_ASAP7_75t_L g2384 ( 
.A1(n_2346),
.A2(n_2348),
.B(n_2354),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2350),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2362),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2364),
.B(n_2325),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2370),
.B(n_2317),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2368),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2371),
.Y(n_2390)
);

XNOR2xp5_ASAP7_75t_L g2391 ( 
.A(n_2357),
.B(n_2307),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2349),
.B(n_2319),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2373),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2372),
.Y(n_2394)
);

INVxp67_ASAP7_75t_L g2395 ( 
.A(n_2365),
.Y(n_2395)
);

INVx2_ASAP7_75t_SL g2396 ( 
.A(n_2358),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2372),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2353),
.B(n_2319),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_R g2399 ( 
.A(n_2358),
.B(n_2337),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2383),
.B(n_2360),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2387),
.B(n_2364),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2395),
.B(n_2360),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2395),
.B(n_2363),
.Y(n_2403)
);

NOR3xp33_ASAP7_75t_L g2404 ( 
.A(n_2384),
.B(n_2367),
.C(n_2375),
.Y(n_2404)
);

AOI211xp5_ASAP7_75t_L g2405 ( 
.A1(n_2391),
.A2(n_2374),
.B(n_2351),
.C(n_2327),
.Y(n_2405)
);

NOR3xp33_ASAP7_75t_L g2406 ( 
.A(n_2378),
.B(n_2328),
.C(n_2336),
.Y(n_2406)
);

AOI211xp5_ASAP7_75t_L g2407 ( 
.A1(n_2398),
.A2(n_2336),
.B(n_2329),
.C(n_2331),
.Y(n_2407)
);

NOR3xp33_ASAP7_75t_L g2408 ( 
.A(n_2392),
.B(n_2326),
.C(n_2344),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2396),
.B(n_2369),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2380),
.B(n_2344),
.Y(n_2410)
);

XNOR2x1_ASAP7_75t_L g2411 ( 
.A(n_2382),
.B(n_2185),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2377),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_L g2413 ( 
.A(n_2380),
.B(n_2331),
.C(n_2326),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2394),
.B(n_2296),
.Y(n_2414)
);

AO22x2_ASAP7_75t_L g2415 ( 
.A1(n_2401),
.A2(n_2389),
.B1(n_2385),
.B2(n_2393),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2404),
.A2(n_2379),
.B1(n_2376),
.B2(n_2388),
.Y(n_2416)
);

AOI21xp33_ASAP7_75t_SL g2417 ( 
.A1(n_2400),
.A2(n_2397),
.B(n_2390),
.Y(n_2417)
);

NAND4xp25_ASAP7_75t_SL g2418 ( 
.A(n_2405),
.B(n_2376),
.C(n_2386),
.D(n_2381),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2402),
.B(n_2296),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2406),
.B(n_2399),
.Y(n_2420)
);

NOR2xp67_ASAP7_75t_L g2421 ( 
.A(n_2413),
.B(n_2399),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_R g2422 ( 
.A(n_2412),
.B(n_2127),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2409),
.B(n_2271),
.Y(n_2423)
);

AOI221xp5_ASAP7_75t_L g2424 ( 
.A1(n_2403),
.A2(n_2299),
.B1(n_2284),
.B2(n_2273),
.C(n_2271),
.Y(n_2424)
);

A2O1A1Ixp33_ASAP7_75t_L g2425 ( 
.A1(n_2410),
.A2(n_2299),
.B(n_2284),
.C(n_2273),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2407),
.A2(n_2299),
.B(n_2284),
.Y(n_2426)
);

NOR2xp67_ASAP7_75t_L g2427 ( 
.A(n_2414),
.B(n_2271),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2408),
.B(n_2411),
.Y(n_2428)
);

OAI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2416),
.A2(n_2273),
.B1(n_2245),
.B2(n_2192),
.Y(n_2429)
);

CKINVDCx6p67_ASAP7_75t_R g2430 ( 
.A(n_2420),
.Y(n_2430)
);

NAND2xp33_ASAP7_75t_SL g2431 ( 
.A(n_2422),
.B(n_2065),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_R g2432 ( 
.A(n_2418),
.B(n_2127),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_SL g2433 ( 
.A(n_2421),
.B(n_2192),
.Y(n_2433)
);

CKINVDCx20_ASAP7_75t_R g2434 ( 
.A(n_2428),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2427),
.Y(n_2435)
);

AOI322xp5_ASAP7_75t_L g2436 ( 
.A1(n_2423),
.A2(n_2207),
.A3(n_2208),
.B1(n_2209),
.B2(n_2173),
.C1(n_2166),
.C2(n_2158),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2415),
.B(n_2201),
.Y(n_2437)
);

NOR3xp33_ASAP7_75t_L g2438 ( 
.A(n_2435),
.B(n_2417),
.C(n_2419),
.Y(n_2438)
);

AOI211xp5_ASAP7_75t_L g2439 ( 
.A1(n_2432),
.A2(n_2426),
.B(n_2424),
.C(n_2415),
.Y(n_2439)
);

NOR2x1_ASAP7_75t_L g2440 ( 
.A(n_2434),
.B(n_2425),
.Y(n_2440)
);

XOR2x1_ASAP7_75t_L g2441 ( 
.A(n_2430),
.B(n_2429),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2433),
.B(n_2189),
.Y(n_2442)
);

NOR3xp33_ASAP7_75t_L g2443 ( 
.A(n_2431),
.B(n_2207),
.C(n_2208),
.Y(n_2443)
);

OAI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2437),
.A2(n_2209),
.B(n_2236),
.Y(n_2444)
);

NOR2x1_ASAP7_75t_L g2445 ( 
.A(n_2436),
.B(n_2203),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2440),
.B(n_2189),
.Y(n_2446)
);

HB1xp67_ASAP7_75t_L g2447 ( 
.A(n_2441),
.Y(n_2447)
);

OAI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2439),
.A2(n_2246),
.B1(n_2226),
.B2(n_2213),
.Y(n_2448)
);

NAND3xp33_ASAP7_75t_SL g2449 ( 
.A(n_2438),
.B(n_2186),
.C(n_2166),
.Y(n_2449)
);

OAI221xp5_ASAP7_75t_SL g2450 ( 
.A1(n_2443),
.A2(n_2158),
.B1(n_2221),
.B2(n_2215),
.C(n_2186),
.Y(n_2450)
);

INVx5_ASAP7_75t_L g2451 ( 
.A(n_2442),
.Y(n_2451)
);

AOI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2444),
.A2(n_2173),
.B1(n_2185),
.B2(n_2188),
.C(n_2174),
.Y(n_2452)
);

BUFx4f_ASAP7_75t_SL g2453 ( 
.A(n_2447),
.Y(n_2453)
);

NOR3xp33_ASAP7_75t_L g2454 ( 
.A(n_2448),
.B(n_2445),
.C(n_2175),
.Y(n_2454)
);

NOR3xp33_ASAP7_75t_L g2455 ( 
.A(n_2449),
.B(n_2188),
.C(n_2185),
.Y(n_2455)
);

NOR3xp33_ASAP7_75t_L g2456 ( 
.A(n_2446),
.B(n_2188),
.C(n_2178),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2451),
.Y(n_2457)
);

NOR2x1p5_ASAP7_75t_L g2458 ( 
.A(n_2457),
.B(n_2451),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2454),
.A2(n_2450),
.B(n_2452),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2458),
.A2(n_2453),
.B1(n_2456),
.B2(n_2455),
.Y(n_2460)
);

INVxp67_ASAP7_75t_L g2461 ( 
.A(n_2460),
.Y(n_2461)
);

OAI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2460),
.A2(n_2459),
.B(n_2178),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2462),
.A2(n_2173),
.B(n_1986),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2461),
.B(n_2163),
.Y(n_2464)
);

AOI21xp33_ASAP7_75t_SL g2465 ( 
.A1(n_2464),
.A2(n_2077),
.B(n_2180),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2463),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_SL g2467 ( 
.A1(n_2466),
.A2(n_2109),
.B1(n_2061),
.B2(n_2165),
.Y(n_2467)
);

OAI221xp5_ASAP7_75t_R g2468 ( 
.A1(n_2467),
.A2(n_2465),
.B1(n_2025),
.B2(n_1966),
.C(n_2061),
.Y(n_2468)
);

AOI211xp5_ASAP7_75t_L g2469 ( 
.A1(n_2468),
.A2(n_2174),
.B(n_2172),
.C(n_1961),
.Y(n_2469)
);


endmodule