module fake_jpeg_16763_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_2),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_52),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_2),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_67),
.B1(n_66),
.B2(n_54),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_103)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_67),
.B1(n_66),
.B2(n_64),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_98),
.B1(n_103),
.B2(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_59),
.B1(n_63),
.B2(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_6),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_60),
.C(n_49),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_85),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_65),
.B1(n_60),
.B2(n_59),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_57),
.B1(n_53),
.B2(n_50),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_48),
.B1(n_65),
.B2(n_20),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_113),
.A3(n_17),
.B1(n_46),
.B2(n_34),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_18),
.B1(n_40),
.B2(n_38),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_110),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_16),
.B1(n_36),
.B2(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_4),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_100),
.B1(n_113),
.B2(n_27),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_121),
.Y(n_130)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_124),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_6),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_7),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_124),
.B1(n_116),
.B2(n_123),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_133),
.A2(n_125),
.B1(n_122),
.B2(n_106),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_129),
.B(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_133),
.B(n_26),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_135),
.C(n_110),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_139),
.A2(n_141),
.B(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_146),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_144),
.B1(n_95),
.B2(n_120),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_145),
.C(n_148),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.C(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_149),
.B(n_7),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_21),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_15),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_23),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_14),
.C(n_32),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_13),
.C(n_30),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_28),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_8),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_99),
.B1(n_111),
.B2(n_11),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);


endmodule