module fake_jpeg_3215_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_65),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_58),
.B(n_78),
.Y(n_130)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_74),
.Y(n_165)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g137 ( 
.A(n_76),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_91),
.B(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g177 ( 
.A(n_103),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_15),
.B(n_26),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_104),
.A2(n_30),
.B(n_37),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_105),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_145),
.Y(n_166)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_58),
.B(n_34),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_49),
.A2(n_26),
.B1(n_34),
.B2(n_42),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_24),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_34),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_50),
.B(n_42),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_42),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_155),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_26),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_5),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_70),
.A2(n_47),
.B1(n_30),
.B2(n_24),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_70),
.B(n_23),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_163),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_98),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_99),
.B(n_23),
.C(n_28),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_47),
.Y(n_172)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_101),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_174),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_30),
.B1(n_47),
.B2(n_24),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_159),
.B1(n_20),
.B2(n_21),
.Y(n_227)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_137),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_192),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_105),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_100),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_29),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_200),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_139),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_106),
.B(n_110),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_144),
.B(n_43),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_206),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_207),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_43),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_212),
.Y(n_229)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

BUFx4f_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_132),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_107),
.B(n_29),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_109),
.B(n_129),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_21),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_122),
.B1(n_125),
.B2(n_112),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_235),
.B1(n_250),
.B2(n_193),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_138),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_139),
.C(n_121),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_238),
.C(n_209),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_173),
.Y(n_234)
);

BUFx16f_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_175),
.A2(n_122),
.B1(n_125),
.B2(n_151),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_136),
.C(n_117),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_239),
.B(n_188),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_190),
.A2(n_113),
.B1(n_141),
.B2(n_63),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_195),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_255),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_182),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_220),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_254),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_233),
.B(n_217),
.C(n_229),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_212),
.B1(n_214),
.B2(n_200),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_241),
.B1(n_236),
.B2(n_240),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_264),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_174),
.B1(n_166),
.B2(n_113),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_273),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_174),
.B1(n_141),
.B2(n_167),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_223),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_270),
.Y(n_292)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_262),
.A2(n_224),
.B1(n_248),
.B2(n_222),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_127),
.B1(n_131),
.B2(n_133),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_213),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_187),
.B(n_29),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_265),
.A2(n_253),
.B(n_281),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_220),
.Y(n_266)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_280),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_170),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_268),
.B(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_204),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_231),
.B(n_128),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_271),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_250),
.A2(n_157),
.B1(n_135),
.B2(n_133),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_277),
.B1(n_279),
.B2(n_281),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_131),
.B1(n_79),
.B2(n_72),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_225),
.B(n_184),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_283),
.Y(n_288)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_227),
.A2(n_135),
.B1(n_157),
.B2(n_52),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_247),
.B(n_197),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_227),
.A2(n_230),
.B1(n_247),
.B2(n_240),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_221),
.B(n_171),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_221),
.B(n_189),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_285),
.B(n_279),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_256),
.B1(n_258),
.B2(n_252),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_287),
.A2(n_315),
.B1(n_277),
.B2(n_272),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_236),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_289),
.B(n_306),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_253),
.Y(n_318)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_227),
.A3(n_251),
.B1(n_215),
.B2(n_242),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_258),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_177),
.C(n_222),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_298),
.C(n_299),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_215),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_219),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_219),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_307),
.C(n_265),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_304),
.A2(n_274),
.B1(n_262),
.B2(n_266),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_305),
.A2(n_265),
.B(n_269),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_244),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_244),
.C(n_117),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

INVx13_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_242),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_310),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_257),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_224),
.B1(n_178),
.B2(n_202),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_320),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_312),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_321),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_344),
.B1(n_320),
.B2(n_345),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_253),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_291),
.A2(n_271),
.B1(n_264),
.B2(n_269),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_294),
.B1(n_301),
.B2(n_303),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_268),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_337),
.C(n_343),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_308),
.B(n_259),
.Y(n_328)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_328),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_308),
.B(n_259),
.Y(n_329)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_330),
.A2(n_254),
.B1(n_216),
.B2(n_286),
.Y(n_383)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_302),
.Y(n_332)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_291),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_342),
.Y(n_351)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_335),
.A2(n_305),
.B(n_294),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_282),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_271),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_349),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_312),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_266),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_287),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_345),
.Y(n_354)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_293),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_348),
.Y(n_353)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_269),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_307),
.C(n_301),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_352),
.A2(n_376),
.B1(n_383),
.B2(n_344),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_298),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_356),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_297),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_374),
.C(n_350),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_311),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_363),
.C(n_375),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_322),
.A2(n_290),
.B1(n_284),
.B2(n_269),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_362),
.A2(n_330),
.B1(n_318),
.B2(n_323),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_319),
.B(n_311),
.Y(n_363)
);

OAI21xp33_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_372),
.B(n_348),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_365),
.A2(n_249),
.B1(n_237),
.B2(n_346),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_284),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_273),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_324),
.A2(n_290),
.B(n_315),
.C(n_313),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_339),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_379),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_273),
.C(n_160),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_321),
.B(n_316),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_328),
.A2(n_290),
.B1(n_300),
.B2(n_263),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_342),
.B(n_248),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_336),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_329),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_399),
.Y(n_427)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_387),
.A2(n_376),
.B1(n_378),
.B2(n_380),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_323),
.C(n_318),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_391),
.C(n_398),
.Y(n_416)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_335),
.C(n_332),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_392),
.A2(n_362),
.B1(n_372),
.B2(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_367),
.A2(n_357),
.B(n_364),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_394),
.A2(n_411),
.B1(n_415),
.B2(n_383),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_331),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_408),
.Y(n_420)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_334),
.C(n_347),
.Y(n_398)
);

XOR2x2_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_326),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_405),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_326),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_403),
.B(n_404),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_326),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_384),
.B(n_263),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_357),
.B(n_340),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_37),
.B(n_45),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_384),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_338),
.C(n_160),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_410),
.C(n_412),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_352),
.B(n_216),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_346),
.B(n_261),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_201),
.C(n_185),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_366),
.B(n_368),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_414),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_249),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_370),
.C(n_371),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_423),
.C(n_431),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_402),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_142),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_371),
.C(n_368),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_429),
.B1(n_430),
.B2(n_436),
.Y(n_450)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_387),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_401),
.A2(n_378),
.B1(n_382),
.B2(n_380),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_407),
.A2(n_382),
.B1(n_237),
.B2(n_211),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_206),
.C(n_187),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_237),
.C(n_243),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_403),
.C(n_391),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_388),
.B(n_261),
.CI(n_124),
.CON(n_435),
.SN(n_435)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_400),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_196),
.B1(n_207),
.B2(n_132),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_8),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_SL g461 ( 
.A1(n_438),
.A2(n_28),
.B(n_46),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_440),
.A2(n_412),
.B(n_45),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_448),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_419),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_409),
.C(n_404),
.Y(n_447)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_399),
.C(n_405),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_452),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_111),
.C(n_61),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_436),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_142),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_454),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_53),
.C(n_62),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_420),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_455),
.A2(n_461),
.B(n_463),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_83),
.C(n_69),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_456),
.B(n_457),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_439),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_424),
.A2(n_151),
.B(n_43),
.Y(n_458)
);

AO21x1_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_460),
.B(n_19),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_433),
.A2(n_74),
.B1(n_68),
.B2(n_45),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_462),
.C(n_465),
.Y(n_482)
);

OAI321xp33_ASAP7_75t_L g460 ( 
.A1(n_438),
.A2(n_37),
.A3(n_28),
.B1(n_46),
.B2(n_20),
.C(n_21),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_430),
.A2(n_143),
.B1(n_193),
.B2(n_46),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_12),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_416),
.B(n_20),
.C(n_19),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_467),
.B(n_474),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_417),
.C(n_432),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_472),
.Y(n_498)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_470),
.Y(n_489)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_431),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_417),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_443),
.A2(n_426),
.B(n_434),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_25),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_421),
.C(n_437),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_477),
.B(n_479),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_434),
.C(n_440),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_442),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_484),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_441),
.C(n_435),
.Y(n_484)
);

NAND2x1_ASAP7_75t_SL g485 ( 
.A(n_464),
.B(n_435),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_479),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_456),
.B(n_446),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_486),
.A2(n_471),
.B1(n_8),
.B2(n_10),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_473),
.A2(n_467),
.B(n_485),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_495),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_483),
.A2(n_450),
.B(n_458),
.Y(n_488)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_492),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_480),
.A2(n_448),
.B1(n_451),
.B2(n_454),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_5),
.B1(n_11),
.B2(n_2),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_143),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_193),
.C(n_143),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_499),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_19),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_142),
.C(n_27),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_502),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_0),
.C(n_1),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_476),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_504),
.B(n_508),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_489),
.A2(n_480),
.B1(n_475),
.B2(n_482),
.Y(n_505)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_505),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_466),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_475),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_512),
.B(n_516),
.Y(n_522)
);

AOI321xp33_ASAP7_75t_L g513 ( 
.A1(n_490),
.A2(n_5),
.A3(n_11),
.B1(n_10),
.B2(n_12),
.C(n_4),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_513),
.Y(n_518)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_499),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_497),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_525),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_511),
.A2(n_510),
.B(n_491),
.Y(n_520)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_520),
.A2(n_526),
.B(n_517),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_503),
.A2(n_488),
.B(n_501),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_521),
.B(n_506),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_496),
.C(n_500),
.Y(n_525)
);

AOI322xp5_ASAP7_75t_L g526 ( 
.A1(n_505),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.C1(n_502),
.C2(n_514),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_527),
.A2(n_530),
.B(n_531),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_506),
.C(n_507),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_528),
.B(n_532),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_524),
.B(n_0),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_529),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_4),
.C(n_0),
.Y(n_532)
);

INVx11_ASAP7_75t_L g533 ( 
.A(n_521),
.Y(n_533)
);

AOI21xp33_ASAP7_75t_L g537 ( 
.A1(n_533),
.A2(n_522),
.B(n_518),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_536),
.A2(n_533),
.B(n_2),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_528),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_539),
.C(n_534),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_540),
.B(n_535),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_2),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_2),
.Y(n_543)
);


endmodule