module fake_ariane_3005_n_805 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_805);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_805;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_783;
wire n_675;

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_94),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_76),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_0),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_36),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_91),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_63),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_43),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_55),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_21),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_89),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_50),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_32),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_4),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_52),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_110),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_19),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_71),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_18),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_98),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_141),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_48),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_6),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_112),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_8),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_93),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_33),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_13),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_73),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_84),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_0),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_189),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_165),
.A2(n_69),
.B(n_157),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_213),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_1),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_200),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_184),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_1),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_2),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_2),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

CKINVDCx11_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_160),
.B(n_3),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_169),
.A2(n_74),
.B(n_155),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_3),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_166),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_175),
.B(n_5),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g255 ( 
.A(n_187),
.B(n_7),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_193),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_195),
.B(n_7),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_226),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_258),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_239),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_201),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_232),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_219),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_215),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_227),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_227),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_237),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_R g275 ( 
.A(n_231),
.B(n_162),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_231),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_R g279 ( 
.A(n_231),
.B(n_170),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_242),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_R g285 ( 
.A(n_250),
.B(n_171),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_246),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_229),
.B(n_173),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_183),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_234),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_245),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_236),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_254),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_216),
.B(n_185),
.Y(n_299)
);

NOR2x1p5_ASAP7_75t_L g300 ( 
.A(n_217),
.B(n_209),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_222),
.B(n_188),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_251),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_228),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_R g304 ( 
.A(n_234),
.B(n_190),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_228),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_255),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_217),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_256),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_248),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_292),
.A2(n_256),
.B1(n_248),
.B2(n_255),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_233),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_284),
.B(n_233),
.Y(n_318)
);

NOR2x1p5_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_244),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_244),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_252),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_289),
.Y(n_322)
);

NAND2xp33_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_252),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_269),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_257),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_257),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_211),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_R g332 ( 
.A(n_260),
.B(n_197),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_269),
.B(n_274),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_265),
.B(n_238),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_267),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_249),
.C(n_238),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_277),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_220),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_270),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_293),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_221),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_285),
.B(n_235),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_268),
.B(n_235),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_198),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_285),
.B(n_203),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_275),
.B(n_204),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_275),
.B(n_221),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_221),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_263),
.B(n_207),
.Y(n_360)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_271),
.B(n_223),
.Y(n_361)
);

BUFx8_ASAP7_75t_L g362 ( 
.A(n_261),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_284),
.B(n_208),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_277),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_223),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_302),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_264),
.B(n_210),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_262),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_298),
.B(n_182),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g373 ( 
.A(n_292),
.B(n_159),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_322),
.B(n_247),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_312),
.A2(n_182),
.B1(n_223),
.B2(n_224),
.Y(n_378)
);

CKINVDCx8_ASAP7_75t_R g379 ( 
.A(n_322),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_8),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_342),
.A2(n_182),
.B1(n_10),
.B2(n_11),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_327),
.B(n_182),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_9),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_9),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_330),
.A2(n_182),
.B1(n_12),
.B2(n_13),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_330),
.B(n_182),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_331),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_14),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_320),
.B(n_15),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_336),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_15),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_325),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_309),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_331),
.A2(n_22),
.B(n_23),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_310),
.B(n_24),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_341),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_25),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_309),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_405)
);

BUFx12f_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_354),
.B(n_29),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_354),
.B(n_31),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_357),
.B(n_34),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_35),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_315),
.B(n_37),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_373),
.A2(n_158),
.B1(n_39),
.B2(n_40),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_323),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_314),
.B(n_44),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_367),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_311),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_369),
.B(n_45),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_365),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_366),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_343),
.Y(n_426)
);

NOR2x1p5_ASAP7_75t_L g427 ( 
.A(n_364),
.B(n_154),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_354),
.B(n_46),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_354),
.B(n_47),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_363),
.B(n_51),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_351),
.B(n_53),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_311),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_319),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_350),
.B(n_54),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_372),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_317),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_317),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_L g442 ( 
.A(n_317),
.B(n_60),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_317),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_391),
.A2(n_318),
.B(n_349),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_351),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_386),
.A2(n_355),
.B1(n_356),
.B2(n_370),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_390),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_344),
.B(n_370),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_441),
.A2(n_358),
.B(n_352),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_443),
.A2(n_348),
.B(n_313),
.Y(n_454)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_407),
.A2(n_348),
.B(n_313),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_348),
.Y(n_456)
);

O2A1O1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_396),
.A2(n_394),
.B(n_382),
.C(n_392),
.Y(n_457)
);

O2A1O1Ixp33_ASAP7_75t_SL g458 ( 
.A1(n_410),
.A2(n_428),
.B(n_430),
.C(n_400),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_402),
.A2(n_411),
.B(n_431),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_313),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_L g462 ( 
.A1(n_389),
.A2(n_311),
.B(n_62),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_61),
.C(n_64),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_65),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_384),
.A2(n_66),
.B(n_67),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_411),
.A2(n_438),
.B(n_377),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_409),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_389),
.A2(n_68),
.B1(n_75),
.B2(n_77),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_SL g469 ( 
.A1(n_383),
.A2(n_78),
.B(n_79),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_377),
.A2(n_80),
.B(n_81),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_424),
.B(n_82),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_424),
.B(n_83),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_401),
.B(n_85),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_442),
.A2(n_407),
.B(n_440),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_379),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_401),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_435),
.B(n_412),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_86),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_436),
.A2(n_87),
.B(n_90),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_397),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_385),
.A2(n_92),
.B(n_95),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_383),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_393),
.A2(n_103),
.B(n_108),
.C(n_109),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_395),
.B(n_111),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_387),
.B(n_153),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_115),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_399),
.A2(n_117),
.B(n_119),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_121),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_423),
.B(n_123),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_426),
.Y(n_496)
);

O2A1O1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_414),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_497)
);

NAND2x1p5_ASAP7_75t_L g498 ( 
.A(n_420),
.B(n_128),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_421),
.A2(n_416),
.B(n_398),
.C(n_405),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_415),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_452),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_452),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_461),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_478),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_466),
.A2(n_378),
.B(n_416),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_485),
.Y(n_511)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_499),
.A2(n_398),
.B(n_405),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_427),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_480),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_415),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_419),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_490),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_480),
.B(n_425),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_459),
.A2(n_381),
.B(n_439),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_479),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_464),
.B(n_129),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_477),
.B(n_132),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_467),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_449),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_455),
.A2(n_134),
.B(n_135),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_444),
.A2(n_137),
.B(n_139),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_477),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_474),
.A2(n_140),
.B(n_142),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_475),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_454),
.A2(n_143),
.B(n_144),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_448),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_491),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_500),
.B(n_145),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_146),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_493),
.A2(n_147),
.B(n_148),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_483),
.B(n_150),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_492),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_481),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_488),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_471),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_457),
.B(n_151),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_494),
.B(n_152),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_472),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_537),
.A2(n_462),
.B(n_469),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_504),
.B(n_447),
.Y(n_555)
);

AO21x1_ASAP7_75t_SL g556 ( 
.A1(n_550),
.A2(n_470),
.B(n_468),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_507),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_510),
.A2(n_451),
.B(n_465),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_512),
.A2(n_486),
.B1(n_463),
.B2(n_495),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_516),
.B(n_487),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_534),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

BUFx2_ASAP7_75t_SL g563 ( 
.A(n_533),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_505),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_509),
.B(n_484),
.Y(n_565)
);

CKINVDCx11_ASAP7_75t_R g566 ( 
.A(n_525),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g567 ( 
.A1(n_510),
.A2(n_450),
.B(n_482),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_505),
.B(n_458),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_505),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_525),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_519),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_549),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_519),
.B(n_497),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_541),
.B(n_548),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_508),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_523),
.A2(n_526),
.B1(n_522),
.B2(n_545),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_523),
.B(n_522),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_531),
.B(n_517),
.Y(n_580)
);

BUFx12f_ASAP7_75t_L g581 ( 
.A(n_536),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_531),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_540),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_512),
.A2(n_523),
.B1(n_526),
.B2(n_522),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_549),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_536),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_518),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_535),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_539),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

INVx8_ASAP7_75t_L g595 ( 
.A(n_526),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_527),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_SL g597 ( 
.A(n_589),
.B(n_552),
.C(n_529),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_555),
.A2(n_526),
.B1(n_547),
.B2(n_546),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_555),
.B(n_526),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_561),
.B(n_522),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_544),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_566),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_546),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_R g605 ( 
.A(n_589),
.B(n_539),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_524),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_SL g608 ( 
.A(n_578),
.B(n_551),
.C(n_513),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_584),
.A2(n_549),
.B1(n_513),
.B2(n_527),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_590),
.B(n_534),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_R g611 ( 
.A(n_562),
.B(n_503),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_572),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_584),
.B(n_503),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_579),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_582),
.B(n_549),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_584),
.A2(n_560),
.B1(n_585),
.B2(n_554),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_563),
.B(n_530),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_566),
.B(n_530),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_571),
.B(n_503),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_596),
.B(n_506),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_576),
.B(n_506),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_584),
.A2(n_543),
.B1(n_524),
.B2(n_528),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_584),
.B(n_579),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_543),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_577),
.B(n_506),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_R g627 ( 
.A(n_579),
.B(n_514),
.Y(n_627)
);

O2A1O1Ixp33_ASAP7_75t_SL g628 ( 
.A1(n_575),
.A2(n_514),
.B(n_520),
.C(n_542),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_586),
.A2(n_579),
.B1(n_574),
.B2(n_591),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_583),
.B(n_514),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_587),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_520),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_570),
.B(n_528),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_581),
.B(n_532),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_553),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_R g636 ( 
.A(n_573),
.B(n_532),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_592),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_565),
.B(n_535),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_585),
.B(n_542),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_556),
.A2(n_521),
.B1(n_574),
.B2(n_594),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_573),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_595),
.A2(n_521),
.B1(n_593),
.B2(n_588),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_SL g644 ( 
.A(n_553),
.B(n_564),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_559),
.B(n_553),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_553),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_621),
.B(n_588),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_639),
.B(n_588),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_640),
.B(n_573),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_637),
.Y(n_650)
);

AO21x2_ASAP7_75t_L g651 ( 
.A1(n_597),
.A2(n_592),
.B(n_567),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_607),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_558),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_570),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_626),
.B(n_558),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_604),
.B(n_570),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_641),
.B(n_568),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_638),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_638),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_612),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_630),
.B(n_564),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_604),
.B(n_564),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_616),
.A2(n_564),
.B1(n_595),
.B2(n_599),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_597),
.A2(n_595),
.B(n_645),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_603),
.B(n_595),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_610),
.B(n_619),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_633),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_614),
.B(n_642),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_614),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_631),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_618),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_615),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_615),
.Y(n_673)
);

OAI332xp33_ASAP7_75t_L g674 ( 
.A1(n_605),
.A2(n_611),
.A3(n_620),
.B1(n_608),
.B2(n_598),
.B3(n_634),
.C1(n_617),
.C2(n_636),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_646),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_633),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_598),
.A2(n_629),
.B1(n_624),
.B2(n_602),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_642),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_629),
.B(n_601),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_643),
.B(n_613),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_628),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_643),
.B(n_613),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_606),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_635),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_650),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_650),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_678),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_649),
.B(n_608),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_649),
.B(n_606),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_652),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_666),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_652),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_648),
.B(n_606),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_648),
.B(n_623),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_670),
.B(n_600),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_668),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_668),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_672),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_672),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_653),
.B(n_625),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_653),
.B(n_635),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_660),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_685),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_680),
.A2(n_683),
.B1(n_657),
.B2(n_664),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_673),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_656),
.B(n_635),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_655),
.B(n_632),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_680),
.B(n_632),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_671),
.B(n_632),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_655),
.B(n_609),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_673),
.B(n_644),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_669),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_669),
.B(n_627),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_647),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_647),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_658),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_716),
.B(n_667),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_697),
.B(n_667),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_697),
.B(n_683),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_688),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_686),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_713),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_SL g724 ( 
.A1(n_705),
.A2(n_675),
.B1(n_665),
.B2(n_677),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_698),
.B(n_676),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_699),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_700),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_706),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_692),
.B(n_698),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_686),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_702),
.B(n_676),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_687),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_712),
.B(n_715),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_691),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_687),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_702),
.B(n_679),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_717),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_717),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_701),
.B(n_679),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_711),
.B(n_659),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_720),
.B(n_689),
.Y(n_741)
);

OAI33xp33_ASAP7_75t_L g742 ( 
.A1(n_724),
.A2(n_733),
.A3(n_723),
.B1(n_729),
.B2(n_726),
.B3(n_728),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_720),
.B(n_689),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_734),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_738),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_734),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_722),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_721),
.A2(n_696),
.B(n_675),
.C(n_710),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_736),
.B(n_701),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_736),
.A2(n_696),
.B1(n_695),
.B2(n_711),
.Y(n_750)
);

INVxp33_ASAP7_75t_L g751 ( 
.A(n_731),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_750),
.B(n_738),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_L g753 ( 
.A1(n_750),
.A2(n_740),
.B1(n_727),
.B2(n_714),
.C(n_722),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_743),
.A2(n_704),
.B1(n_739),
.B2(n_737),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_745),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_742),
.A2(n_695),
.B1(n_709),
.B2(n_739),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_741),
.B(n_735),
.Y(n_757)
);

XNOR2xp5_ASAP7_75t_L g758 ( 
.A(n_743),
.B(n_709),
.Y(n_758)
);

AND2x4_ASAP7_75t_SL g759 ( 
.A(n_756),
.B(n_749),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_L g760 ( 
.A1(n_752),
.A2(n_748),
.B(n_682),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_758),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_754),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_757),
.B(n_732),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_753),
.B(n_748),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_760),
.A2(n_674),
.B(n_751),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_762),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_761),
.Y(n_768)
);

AOI211xp5_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_682),
.B(n_707),
.C(n_708),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_767),
.B(n_763),
.C(n_764),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_768),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_766),
.A2(n_759),
.B1(n_657),
.B2(n_709),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_R g773 ( 
.A(n_771),
.B(n_704),
.Y(n_773)
);

OAI211xp5_ASAP7_75t_L g774 ( 
.A1(n_770),
.A2(n_769),
.B(n_704),
.C(n_685),
.Y(n_774)
);

AOI221xp5_ASAP7_75t_L g775 ( 
.A1(n_772),
.A2(n_747),
.B1(n_746),
.B2(n_744),
.C(n_730),
.Y(n_775)
);

AOI222xp33_ASAP7_75t_L g776 ( 
.A1(n_771),
.A2(n_730),
.B1(n_663),
.B2(n_725),
.C1(n_662),
.C2(n_693),
.Y(n_776)
);

NOR2x1p5_ASAP7_75t_L g777 ( 
.A(n_773),
.B(n_774),
.Y(n_777)
);

NOR2x1_ASAP7_75t_L g778 ( 
.A(n_776),
.B(n_651),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_775),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_773),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_773),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_777),
.A2(n_719),
.B1(n_718),
.B2(n_725),
.Y(n_782)
);

NAND2x1p5_ASAP7_75t_L g783 ( 
.A(n_781),
.B(n_714),
.Y(n_783)
);

AO22x2_ASAP7_75t_L g784 ( 
.A1(n_780),
.A2(n_731),
.B1(n_684),
.B2(n_654),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_779),
.B(n_661),
.C(n_708),
.Y(n_785)
);

NAND4xp75_ASAP7_75t_L g786 ( 
.A(n_778),
.B(n_694),
.C(n_690),
.D(n_661),
.Y(n_786)
);

NOR2x1p5_ASAP7_75t_L g787 ( 
.A(n_781),
.B(n_654),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_SL g788 ( 
.A(n_787),
.B(n_782),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_783),
.B(n_694),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_785),
.B(n_651),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_786),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_SL g792 ( 
.A(n_791),
.B(n_784),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_789),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_790),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_788),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_795),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_793),
.A2(n_684),
.B1(n_654),
.B2(n_658),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_794),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_796),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_798),
.A2(n_792),
.B1(n_659),
.B2(n_681),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_799),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_801),
.B(n_800),
.Y(n_802)
);

AOI21x1_ASAP7_75t_L g803 ( 
.A1(n_802),
.A2(n_797),
.B(n_690),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_803),
.B(n_681),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_804),
.A2(n_651),
.B1(n_703),
.B2(n_691),
.Y(n_805)
);


endmodule