module real_jpeg_31522_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_0),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_0),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_0),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_146),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_1),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_1),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_1),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_2),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_2),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_2),
.B(n_210),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_2),
.B(n_480),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_493),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_3),
.B(n_494),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_7),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_7),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_7),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_7),
.B(n_376),
.Y(n_375)
);

NAND2x1_ASAP7_75t_L g438 ( 
.A(n_7),
.B(n_439),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_7),
.B(n_50),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_8),
.B(n_123),
.Y(n_122)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_8),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_8),
.B(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_8),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_8),
.B(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_9),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_9),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_131),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g163 ( 
.A(n_9),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_9),
.B(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_9),
.B(n_190),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_9),
.B(n_467),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_12),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_12),
.B(n_112),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_12),
.B(n_288),
.Y(n_287)
);

NAND2x1_ASAP7_75t_L g300 ( 
.A(n_12),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_12),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_12),
.B(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_14),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_176),
.Y(n_175)
);

AND2x4_ASAP7_75t_SL g284 ( 
.A(n_14),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_14),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_14),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_14),
.B(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_15),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_16),
.B(n_82),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_16),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_16),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_16),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_16),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_16),
.B(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_17),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_454),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_445),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_245),
.C(n_357),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_195),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_147),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_25),
.B(n_147),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_74),
.C(n_98),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_27),
.A2(n_74),
.B1(n_75),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_27),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_46),
.Y(n_27)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_28),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_41),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_30),
.A2(n_31),
.B1(n_464),
.B2(n_468),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_31),
.B(n_36),
.C(n_41),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_31),
.B(n_36),
.C(n_41),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_34),
.Y(n_164)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_40),
.Y(n_482)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_44),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_45),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_47),
.B(n_58),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_47),
.B(n_58),
.Y(n_194)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_53),
.Y(n_97)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_53),
.A2(n_54),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_54),
.B(n_206),
.C(n_209),
.Y(n_382)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.C(n_70),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_70),
.B2(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_60),
.B(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_60),
.A2(n_61),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_60),
.B(n_132),
.C(n_420),
.Y(n_470)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_63),
.Y(n_216)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_63),
.Y(n_285)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_63),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_64),
.Y(n_265)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_68),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_73),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_73),
.Y(n_378)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_97),
.Y(n_75)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_76),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_91),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_81),
.B(n_85),
.C(n_91),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_81),
.B(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2x1_ASAP7_75t_L g346 ( 
.A(n_85),
.B(n_91),
.Y(n_346)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_95),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_96),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_97),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_98),
.B(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_128),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_110),
.B1(n_126),
.B2(n_127),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_108),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_104),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_104),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_107),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_108),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_109),
.Y(n_233)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_126),
.C(n_128),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_118),
.C(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_116),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_116),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2x2_ASAP7_75t_L g386 ( 
.A(n_119),
.B(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_119),
.B(n_206),
.C(n_389),
.Y(n_441)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.C(n_142),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_129),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_174),
.B1(n_175),
.B2(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_130),
.B(n_175),
.C(n_180),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_130),
.A2(n_132),
.B1(n_178),
.B2(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_SL g283 ( 
.A(n_131),
.Y(n_283)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_132),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_132),
.A2(n_267),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_132),
.B(n_400),
.C(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_169),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_149),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_155),
.C(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_165),
.C(n_225),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx4f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_159),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_162),
.A2(n_163),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_197),
.B(n_199),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_192),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_183),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_183),
.C(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_179),
.B2(n_180),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_191),
.C(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_195),
.A2(n_447),
.B(n_448),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_196),
.B(n_200),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_201),
.B(n_360),
.C(n_361),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_228),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_203),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_204),
.B(n_213),
.C(n_227),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_206),
.B(n_257),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_206),
.A2(n_207),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_208),
.A2(n_209),
.B1(n_479),
.B2(n_483),
.Y(n_478)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_220),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_215),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_217),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_219),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_221),
.B(n_393),
.C(n_394),
.Y(n_392)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_225),
.B(n_428),
.C(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_228),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_229),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_232),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_234),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_235),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_236)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g402 ( 
.A(n_242),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_243),
.B(n_370),
.C(n_371),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_244),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_271),
.B(n_356),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_268),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_247),
.B(n_268),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.C(n_255),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_248),
.B(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.C(n_266),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_256),
.B(n_260),
.Y(n_348)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_266),
.B(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_267),
.B(n_396),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_350),
.B(n_355),
.Y(n_271)
);

OAI21x1_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_338),
.B(n_349),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_306),
.B(n_337),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_290),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_275),
.B(n_290),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.C(n_286),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_276),
.A2(n_277),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_284),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_295),
.C(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_300),
.C(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_330),
.B(n_336),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_319),
.B(n_329),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_313),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_341),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_345),
.C(n_347),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_354),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_357),
.A2(n_446),
.B(n_449),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_362),
.B1(n_408),
.B2(n_411),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_359),
.B(n_363),
.Y(n_452)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_383),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_403),
.C(n_410),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_369),
.C(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2x2_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_382),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_379),
.B2(n_381),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_374),
.B(n_381),
.C(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_379),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_379),
.B(n_438),
.Y(n_437)
);

MAJx2_ASAP7_75t_L g475 ( 
.A(n_381),
.B(n_438),
.C(n_440),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_403),
.B2(n_407),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_391),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_386),
.B(n_392),
.C(n_395),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_397),
.Y(n_432)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_403),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.C(n_406),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_412),
.B(n_451),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_434),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_416),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_424),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_417),
.B(n_426),
.C(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_431),
.B2(n_433),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

XOR2x2_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_428),
.Y(n_429)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_431),
.Y(n_433)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_433),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_434),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_444),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_443),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_436),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_436)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_437),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_452),
.B(n_453),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_491),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_486),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_SL g492 ( 
.A(n_456),
.B(n_486),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_461),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.C(n_460),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_473),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_469),
.Y(n_462)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_464),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_484),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.C(n_490),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);


endmodule