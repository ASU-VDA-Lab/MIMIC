module fake_ariane_3275_n_1360 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1360);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1360;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1356;
wire n_1341;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g314 ( 
.A(n_126),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_114),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_171),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_150),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_106),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_109),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_103),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_214),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_180),
.Y(n_327)
);

CKINVDCx12_ASAP7_75t_R g328 ( 
.A(n_239),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_275),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_59),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_183),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_233),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_145),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_230),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_92),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_266),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_228),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_283),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_167),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_277),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_37),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_140),
.Y(n_344)
);

BUFx8_ASAP7_75t_SL g345 ( 
.A(n_163),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_221),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_191),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_206),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_159),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_74),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_54),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_187),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_116),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_274),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_241),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_35),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_225),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_172),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_200),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_184),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_101),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_31),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_153),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_189),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_202),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_197),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_7),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_246),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_14),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_287),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_278),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_82),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_182),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_9),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_271),
.Y(n_379)
);

BUFx8_ASAP7_75t_SL g380 ( 
.A(n_113),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_284),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_71),
.Y(n_382)
);

BUFx8_ASAP7_75t_SL g383 ( 
.A(n_165),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_128),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_144),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_20),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_7),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_80),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_91),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_178),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_127),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_115),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_25),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_16),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_254),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_207),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_204),
.B(n_273),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_134),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_272),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_186),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_293),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_3),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_55),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_268),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_64),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_12),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_89),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_104),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_48),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_276),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_286),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_15),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_100),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_211),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_75),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_296),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_62),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_232),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_94),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_302),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_195),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_21),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_298),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_108),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_168),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_31),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_235),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_236),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_305),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_65),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_117),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_303),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_73),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_280),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_37),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_216),
.B(n_174),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_205),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_179),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_111),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_215),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_224),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_4),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_21),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_1),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_212),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_264),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_102),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_57),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_253),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_190),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_267),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_16),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_49),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_67),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_259),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_56),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_209),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_161),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_248),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_97),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_257),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_289),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_148),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_155),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_226),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_63),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_141),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_240),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_48),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_28),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_164),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_17),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_223),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_238),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_14),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_143),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_22),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_255),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_213),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_300),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_310),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_234),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_311),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_93),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_53),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_188),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_90),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_256),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_218),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_125),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_251),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_219),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_250),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_22),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_265),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_262),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_129),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_270),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_78),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_44),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_5),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_27),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_220),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_131),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_42),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_281),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_119),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_198),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_45),
.Y(n_511)
);

BUFx8_ASAP7_75t_SL g512 ( 
.A(n_170),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_43),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_288),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_6),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_36),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_269),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_30),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_139),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_17),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_26),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_146),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_137),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_157),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_173),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_142),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_4),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_0),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_345),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_411),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_325),
.B(n_0),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_411),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_338),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_395),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_2),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_338),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_452),
.B(n_52),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_338),
.Y(n_539)
);

OAI22x1_ASAP7_75t_SL g540 ( 
.A1(n_396),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_479),
.Y(n_541)
);

NOR2x1_ASAP7_75t_L g542 ( 
.A(n_365),
.B(n_58),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_338),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_314),
.B(n_8),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_516),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_413),
.B(n_60),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_386),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_502),
.B(n_9),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_315),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_413),
.B(n_61),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_330),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_330),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_316),
.A2(n_10),
.B(n_11),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_404),
.B(n_10),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_319),
.A2(n_11),
.B(n_12),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_343),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_364),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g559 ( 
.A1(n_321),
.A2(n_13),
.B(n_15),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_339),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_502),
.B(n_13),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_371),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_323),
.B(n_18),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_388),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_386),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_408),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_339),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_326),
.B(n_332),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_322),
.A2(n_68),
.B(n_66),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_437),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_362),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_471),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_322),
.A2(n_70),
.B(n_69),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_357),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_373),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_386),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_362),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_386),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_481),
.Y(n_581)
);

AOI22x1_ASAP7_75t_SL g582 ( 
.A1(n_527),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_582)
);

OA21x2_ASAP7_75t_L g583 ( 
.A1(n_334),
.A2(n_19),
.B(n_23),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_387),
.Y(n_584)
);

BUFx12f_ASAP7_75t_L g585 ( 
.A(n_481),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_344),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_378),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_414),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_387),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_504),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_521),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_424),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_344),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_341),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_428),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_494),
.B(n_453),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_318),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_346),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_348),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_350),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_444),
.B(n_24),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_446),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_354),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_501),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_358),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_384),
.B(n_27),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_359),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_454),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_455),
.B(n_28),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_360),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_361),
.B(n_29),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_423),
.B(n_29),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_363),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_352),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_367),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_397),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_368),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_370),
.Y(n_623)
);

BUFx12f_ASAP7_75t_L g624 ( 
.A(n_477),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_372),
.Y(n_625)
);

CKINVDCx11_ASAP7_75t_R g626 ( 
.A(n_402),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_496),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_374),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_407),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_376),
.Y(n_631)
);

BUFx8_ASAP7_75t_L g632 ( 
.A(n_433),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_379),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_381),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_385),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_392),
.A2(n_38),
.B(n_39),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_394),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_507),
.B(n_39),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_513),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_398),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_406),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_409),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_418),
.Y(n_643)
);

BUFx8_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

OA21x2_ASAP7_75t_L g645 ( 
.A1(n_419),
.A2(n_40),
.B(n_41),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_440),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_515),
.Y(n_647)
);

BUFx8_ASAP7_75t_SL g648 ( 
.A(n_380),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_422),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_426),
.B(n_41),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_317),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_518),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_430),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_520),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_465),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_432),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_435),
.B(n_45),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_448),
.B(n_46),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_383),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_320),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_461),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_469),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_478),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_486),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_497),
.B(n_47),
.Y(n_667)
);

BUFx8_ASAP7_75t_SL g668 ( 
.A(n_484),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_517),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_485),
.A2(n_50),
.B1(n_51),
.B2(n_72),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_324),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_487),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_519),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_525),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_399),
.Y(n_675)
);

AO21x2_ASAP7_75t_L g676 ( 
.A1(n_531),
.A2(n_438),
.B(n_328),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_537),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_668),
.Y(n_678)
);

NOR2xp67_ASAP7_75t_L g679 ( 
.A(n_529),
.B(n_327),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_646),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_651),
.B(n_597),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_562),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_564),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_648),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_672),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_571),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_626),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_576),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_533),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_660),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_671),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_546),
.A2(n_498),
.B1(n_505),
.B2(n_491),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_575),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_659),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_552),
.B(n_336),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_537),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_596),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_612),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_537),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_624),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_552),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_550),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_567),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_585),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_553),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_577),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_665),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_614),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_665),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_651),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_588),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_627),
.B(n_526),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_614),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_652),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_539),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_654),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_552),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_535),
.A2(n_417),
.B1(n_468),
.B2(n_401),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_560),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_539),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_560),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_R g724 ( 
.A(n_579),
.B(n_329),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_593),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_572),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_543),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_606),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_627),
.B(n_331),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_622),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_622),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_572),
.B(n_579),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_622),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_572),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_616),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_634),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_634),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_581),
.B(n_500),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_639),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_647),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_634),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_R g743 ( 
.A(n_628),
.B(n_333),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_635),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_544),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_632),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_644),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_590),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_644),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_595),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_R g751 ( 
.A(n_628),
.B(n_581),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_607),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_533),
.B(n_335),
.Y(n_753)
);

AND2x6_ASAP7_75t_L g754 ( 
.A(n_610),
.B(n_349),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_635),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_SL g756 ( 
.A(n_555),
.B(n_337),
.Y(n_756)
);

CKINVDCx16_ASAP7_75t_R g757 ( 
.A(n_538),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_635),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_528),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_543),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_590),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_543),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_675),
.B(n_340),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_536),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_675),
.B(n_342),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_578),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_584),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_690),
.B(n_675),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_759),
.B(n_610),
.Y(n_769)
);

BUFx6f_ASAP7_75t_SL g770 ( 
.A(n_685),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_709),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_757),
.B(n_670),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_682),
.B(n_568),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_690),
.B(n_657),
.Y(n_774)
);

AO221x1_ASAP7_75t_L g775 ( 
.A1(n_693),
.A2(n_621),
.B1(n_655),
.B2(n_599),
.C(n_534),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_766),
.B(n_657),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_766),
.B(n_658),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_764),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_764),
.A2(n_615),
.B(n_667),
.C(n_658),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_754),
.B(n_667),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_754),
.B(n_578),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_712),
.B(n_750),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_763),
.B(n_618),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_754),
.B(n_617),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_754),
.B(n_617),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_SL g786 ( 
.A(n_761),
.B(n_545),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_754),
.B(n_625),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_733),
.B(n_629),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_752),
.B(n_528),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_703),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_765),
.B(n_633),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_748),
.B(n_642),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_751),
.B(n_605),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_681),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_760),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_696),
.B(n_643),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_739),
.B(n_666),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_683),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_707),
.B(n_650),
.C(n_563),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_713),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_707),
.B(n_601),
.Y(n_801)
);

AOI221xp5_ASAP7_75t_L g802 ( 
.A1(n_720),
.A2(n_532),
.B1(n_530),
.B2(n_561),
.C(n_549),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_760),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_767),
.B(n_603),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_684),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_715),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_702),
.B(n_604),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_719),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_714),
.B(n_631),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_687),
.B(n_547),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_689),
.B(n_547),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_745),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_731),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_732),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_734),
.Y(n_815)
);

BUFx6f_ASAP7_75t_SL g816 ( 
.A(n_678),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_756),
.A2(n_561),
.B1(n_549),
.B2(n_613),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_760),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_730),
.B(n_631),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_737),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_738),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_743),
.B(n_641),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_708),
.B(n_638),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_742),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_744),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_704),
.B(n_641),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_755),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_758),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_716),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_753),
.B(n_649),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_725),
.B(n_630),
.C(n_619),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_677),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_697),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_721),
.B(n_649),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_724),
.B(n_556),
.C(n_554),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_725),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_711),
.B(n_637),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_700),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_694),
.B(n_609),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_710),
.B(n_662),
.C(n_566),
.Y(n_840)
);

INVxp33_ASAP7_75t_L g841 ( 
.A(n_679),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_717),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_723),
.B(n_611),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_722),
.B(n_547),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_736),
.B(n_661),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_740),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_726),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_718),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_741),
.B(n_661),
.Y(n_849)
);

INVxp33_ASAP7_75t_L g850 ( 
.A(n_729),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_728),
.B(n_547),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_727),
.B(n_551),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_760),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_735),
.B(n_661),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_762),
.B(n_551),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_676),
.A2(n_551),
.B1(n_623),
.B2(n_620),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_775),
.A2(n_676),
.B1(n_551),
.B2(n_673),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_790),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_794),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_798),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_773),
.B(n_640),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_778),
.B(n_653),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_808),
.B(n_706),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_805),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_771),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_801),
.B(n_656),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_810),
.A2(n_574),
.B(n_569),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_806),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_804),
.B(n_686),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_846),
.Y(n_870)
);

BUFx8_ASAP7_75t_L g871 ( 
.A(n_770),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_814),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_800),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_831),
.A2(n_554),
.B1(n_559),
.B2(n_556),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_809),
.B(n_695),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_815),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_819),
.B(n_691),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_836),
.B(n_705),
.Y(n_878)
);

O2A1O1Ixp5_ASAP7_75t_L g879 ( 
.A1(n_810),
.A2(n_664),
.B(n_663),
.C(n_570),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_813),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_829),
.Y(n_881)
);

AND3x2_ASAP7_75t_SL g882 ( 
.A(n_772),
.B(n_582),
.C(n_680),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_822),
.B(n_793),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_783),
.B(n_559),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_811),
.A2(n_542),
.B(n_583),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_821),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_839),
.B(n_692),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_824),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_825),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_828),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_795),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_779),
.A2(n_636),
.B1(n_645),
.B2(n_583),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_799),
.B(n_698),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_826),
.B(n_699),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_827),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_791),
.B(n_636),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_835),
.A2(n_645),
.B(n_573),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_832),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_833),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_816),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_838),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_795),
.Y(n_903)
);

INVx5_ASAP7_75t_L g904 ( 
.A(n_808),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_797),
.B(n_586),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_780),
.A2(n_582),
.B1(n_540),
.B2(n_669),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_784),
.B(n_586),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_847),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_817),
.A2(n_785),
.B1(n_787),
.B2(n_840),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_795),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_792),
.A2(n_673),
.B1(n_674),
.B2(n_669),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_782),
.B(n_834),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_842),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_768),
.B(n_701),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_796),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_802),
.A2(n_673),
.B1(n_674),
.B2(n_669),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_812),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_774),
.B(n_674),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_853),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_776),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_803),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_777),
.B(n_594),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_788),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_769),
.B(n_746),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_843),
.B(n_747),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_856),
.A2(n_600),
.B1(n_594),
.B2(n_591),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_823),
.B(n_749),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_807),
.B(n_688),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_830),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_811),
.A2(n_351),
.B(n_347),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_835),
.A2(n_600),
.B1(n_592),
.B2(n_557),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_789),
.B(n_541),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_781),
.B(n_349),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_803),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_803),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_841),
.B(n_353),
.Y(n_936)
);

NOR2x1p5_ASAP7_75t_L g937 ( 
.A(n_816),
.B(n_355),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_818),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_837),
.B(n_786),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_818),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_818),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_844),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_844),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_850),
.B(n_848),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_855),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_855),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_845),
.B(n_51),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_852),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_852),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_849),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_904),
.B(n_854),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_861),
.B(n_851),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_861),
.B(n_356),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_883),
.B(n_920),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_943),
.A2(n_369),
.B(n_366),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_869),
.A2(n_866),
.B(n_859),
.C(n_864),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_SL g957 ( 
.A(n_873),
.B(n_375),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_867),
.A2(n_349),
.B(n_76),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_909),
.A2(n_377),
.B1(n_389),
.B2(n_382),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_871),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_860),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_888),
.B(n_390),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_909),
.A2(n_391),
.B(n_400),
.C(n_393),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_SL g964 ( 
.A(n_894),
.B(n_405),
.C(n_403),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_865),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_912),
.A2(n_412),
.B(n_410),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_863),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_866),
.A2(n_463),
.B(n_415),
.C(n_416),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_858),
.B(n_762),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_917),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_871),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_947),
.A2(n_466),
.B1(n_420),
.B2(n_421),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_923),
.A2(n_467),
.B1(n_425),
.B2(n_427),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_863),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_870),
.B(n_548),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_878),
.B(n_429),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_930),
.A2(n_349),
.B(n_79),
.C(n_81),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_933),
.A2(n_434),
.B(n_431),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_933),
.A2(n_439),
.B(n_436),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_901),
.Y(n_980)
);

AO21x2_ASAP7_75t_L g981 ( 
.A1(n_898),
.A2(n_349),
.B(n_548),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_922),
.A2(n_476),
.B(n_442),
.C(n_443),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_925),
.B(n_441),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_928),
.A2(n_881),
.B(n_918),
.C(n_876),
.Y(n_984)
);

OR2x6_ASAP7_75t_L g985 ( 
.A(n_944),
.B(n_548),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_858),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_915),
.B(n_447),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_872),
.A2(n_489),
.B(n_450),
.C(n_451),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_929),
.B(n_449),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_885),
.A2(n_493),
.B1(n_457),
.B2(n_458),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_947),
.B(n_762),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_886),
.A2(n_77),
.B(n_83),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_910),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_857),
.A2(n_506),
.B1(n_459),
.B2(n_460),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_875),
.A2(n_508),
.B1(n_462),
.B2(n_464),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_945),
.A2(n_470),
.B(n_456),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_932),
.A2(n_522),
.B1(n_475),
.B2(n_480),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_884),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_945),
.A2(n_942),
.B(n_897),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_924),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_897),
.A2(n_523),
.B1(n_482),
.B2(n_488),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_936),
.B(n_914),
.C(n_927),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_907),
.A2(n_905),
.B(n_948),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_950),
.B(n_473),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_879),
.A2(n_490),
.B(n_499),
.C(n_509),
.Y(n_1005)
);

BUFx8_ASAP7_75t_SL g1006 ( 
.A(n_910),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_907),
.A2(n_524),
.B(n_514),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_916),
.A2(n_602),
.B1(n_587),
.B2(n_580),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_939),
.A2(n_762),
.B1(n_608),
.B2(n_598),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_937),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_910),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_939),
.A2(n_608),
.B1(n_598),
.B2(n_602),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_887),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_905),
.B(n_598),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_889),
.A2(n_602),
.B(n_587),
.C(n_580),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_899),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_935),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_877),
.B(n_608),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_890),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_891),
.A2(n_587),
.B(n_580),
.C(n_565),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_895),
.B(n_84),
.C(n_85),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_862),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_949),
.A2(n_565),
.B(n_86),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_868),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_946),
.A2(n_565),
.B(n_87),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_1006),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_958),
.A2(n_898),
.B(n_893),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_992),
.A2(n_893),
.B(n_874),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_967),
.B(n_935),
.Y(n_1029)
);

AO21x2_ASAP7_75t_L g1030 ( 
.A1(n_981),
.A2(n_874),
.B(n_862),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_999),
.A2(n_931),
.B(n_903),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_993),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_993),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_993),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_1003),
.A2(n_911),
.B(n_934),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_965),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_961),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_1025),
.A2(n_1023),
.B(n_952),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_1011),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_980),
.Y(n_1040)
);

AO21x2_ASAP7_75t_L g1041 ( 
.A1(n_1005),
.A2(n_911),
.B(n_938),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_1009),
.A2(n_903),
.B(n_892),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_1011),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_954),
.A2(n_919),
.B(n_921),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_1011),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_986),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_963),
.A2(n_913),
.B(n_940),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_956),
.A2(n_941),
.B(n_892),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1022),
.B(n_926),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1024),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_1017),
.Y(n_1051)
);

AO21x2_ASAP7_75t_L g1052 ( 
.A1(n_1014),
.A2(n_880),
.B(n_896),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_960),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_998),
.Y(n_1054)
);

OA21x2_ASAP7_75t_L g1055 ( 
.A1(n_982),
.A2(n_908),
.B(n_902),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_1017),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_977),
.A2(n_900),
.B(n_906),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_1012),
.A2(n_941),
.B(n_88),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_962),
.B(n_970),
.Y(n_1059)
);

BUFx8_ASAP7_75t_L g1060 ( 
.A(n_971),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_974),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_1013),
.Y(n_1062)
);

AO21x2_ASAP7_75t_L g1063 ( 
.A1(n_978),
.A2(n_906),
.B(n_882),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1019),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_983),
.B(n_313),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_991),
.Y(n_1066)
);

AO21x2_ASAP7_75t_L g1067 ( 
.A1(n_979),
.A2(n_95),
.B(n_96),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_969),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_969),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_1007),
.A2(n_98),
.B(n_99),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_980),
.B(n_1000),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_976),
.B(n_105),
.Y(n_1072)
);

BUFx12f_ASAP7_75t_L g1073 ( 
.A(n_1010),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_1016),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_975),
.Y(n_1075)
);

INVx6_ASAP7_75t_L g1076 ( 
.A(n_985),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1004),
.B(n_312),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_953),
.A2(n_955),
.B(n_990),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_964),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_991),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_985),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_989),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_972),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_984),
.A2(n_1020),
.B(n_1015),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_951),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_SL g1086 ( 
.A(n_957),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_1001),
.A2(n_107),
.B(n_110),
.Y(n_1087)
);

AO21x2_ASAP7_75t_L g1088 ( 
.A1(n_968),
.A2(n_112),
.B(n_118),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_994),
.A2(n_120),
.B(n_121),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1062),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1059),
.B(n_1083),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1072),
.A2(n_1002),
.B1(n_959),
.B2(n_997),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1028),
.A2(n_996),
.B(n_988),
.Y(n_1093)
);

OA21x2_ASAP7_75t_L g1094 ( 
.A1(n_1028),
.A2(n_1021),
.B(n_966),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_SL g1095 ( 
.A1(n_1063),
.A2(n_987),
.B1(n_973),
.B2(n_1018),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1027),
.A2(n_1008),
.B(n_995),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1063),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1036),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_1033),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1036),
.Y(n_1100)
);

OA21x2_ASAP7_75t_L g1101 ( 
.A1(n_1027),
.A2(n_130),
.B(n_132),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1050),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1037),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1050),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1046),
.B(n_308),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1033),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_1033),
.Y(n_1107)
);

AO21x2_ASAP7_75t_L g1108 ( 
.A1(n_1052),
.A2(n_133),
.B(n_135),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_1052),
.A2(n_136),
.B(n_138),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1054),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1038),
.A2(n_147),
.B(n_149),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1040),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1064),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_1033),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1082),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1030),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1082),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_1026),
.Y(n_1118)
);

INVxp33_ASAP7_75t_L g1119 ( 
.A(n_1074),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1085),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1038),
.A2(n_1031),
.B(n_1058),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1085),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_1032),
.B(n_156),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1045),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1080),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1066),
.B(n_158),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1045),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1031),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1030),
.Y(n_1129)
);

BUFx10_ASAP7_75t_L g1130 ( 
.A(n_1086),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1044),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1045),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1061),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1077),
.A2(n_160),
.B1(n_162),
.B2(n_166),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1045),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1061),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1079),
.A2(n_169),
.B1(n_175),
.B2(n_176),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1039),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1032),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_SL g1140 ( 
.A1(n_1048),
.A2(n_177),
.B(n_181),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1055),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1026),
.B(n_299),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1035),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1060),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_1086),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1034),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1034),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1106),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1139),
.B(n_1081),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1092),
.A2(n_1068),
.B1(n_1069),
.B2(n_1065),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1091),
.B(n_1069),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_1144),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1119),
.B(n_1071),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1126),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1095),
.A2(n_1049),
.B1(n_1089),
.B2(n_1076),
.Y(n_1155)
);

AND2x2_ASAP7_75t_SL g1156 ( 
.A(n_1097),
.B(n_1089),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1095),
.A2(n_1089),
.B1(n_1076),
.B2(n_1057),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1119),
.B(n_1081),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1113),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_SL g1160 ( 
.A(n_1118),
.B(n_1051),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1139),
.B(n_1039),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1103),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1142),
.B(n_1053),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1112),
.B(n_1053),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1145),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1105),
.B(n_1029),
.Y(n_1166)
);

CKINVDCx16_ASAP7_75t_R g1167 ( 
.A(n_1112),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1106),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1110),
.B(n_1039),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1139),
.B(n_1043),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1098),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_1106),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1117),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1145),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1090),
.B(n_1043),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1120),
.A2(n_1057),
.B1(n_1075),
.B2(n_1047),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1133),
.B(n_1073),
.Y(n_1177)
);

INVx11_ASAP7_75t_L g1178 ( 
.A(n_1130),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1125),
.B(n_1043),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_1139),
.B(n_1073),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1122),
.B(n_1056),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_R g1182 ( 
.A(n_1130),
.B(n_1060),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1136),
.Y(n_1183)
);

INVxp33_ASAP7_75t_L g1184 ( 
.A(n_1106),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1143),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1127),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_R g1187 ( 
.A(n_1099),
.B(n_1056),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_R g1188 ( 
.A(n_1107),
.B(n_1056),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1127),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1100),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_1127),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1126),
.B(n_1051),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1102),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1137),
.B(n_1107),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1146),
.B(n_1078),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1138),
.B(n_1042),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1147),
.B(n_1055),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1114),
.B(n_1087),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1171),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1162),
.B(n_1143),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1196),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1158),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1196),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1190),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1159),
.B(n_1116),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1164),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_1195),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1185),
.B(n_1153),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1148),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1151),
.B(n_1131),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1175),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1173),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1192),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1192),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1154),
.B(n_1128),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1148),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1191),
.B(n_1127),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1193),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1194),
.A2(n_1134),
.B(n_1115),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1197),
.B(n_1129),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1180),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1168),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1181),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1198),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1169),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1179),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1156),
.B(n_1141),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1186),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1189),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1168),
.B(n_1121),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1149),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1180),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1167),
.B(n_1155),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1183),
.B(n_1114),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1177),
.B(n_1138),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1187),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1149),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1176),
.B(n_1102),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1160),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1172),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1163),
.B(n_1124),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1191),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1161),
.B(n_1124),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1157),
.B(n_1104),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1152),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1188),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1166),
.B(n_1132),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1202),
.B(n_1241),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1211),
.B(n_1174),
.Y(n_1249)
);

OAI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_1219),
.A2(n_1150),
.B(n_1184),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1208),
.B(n_1165),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1208),
.B(n_1182),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1212),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1247),
.B(n_1170),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1236),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1247),
.B(n_1135),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1207),
.B(n_1094),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1233),
.A2(n_1101),
.B1(n_1109),
.B2(n_1108),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1210),
.B(n_1094),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1200),
.Y(n_1260)
);

NAND2x1_ASAP7_75t_L g1261 ( 
.A(n_1239),
.B(n_1140),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1226),
.B(n_1123),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1224),
.B(n_1223),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1203),
.B(n_1108),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1229),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1229),
.B(n_1123),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1225),
.Y(n_1267)
);

NOR2x1_ASAP7_75t_L g1268 ( 
.A(n_1236),
.B(n_1070),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1228),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1214),
.B(n_1111),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1201),
.B(n_1093),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1205),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1227),
.B(n_1088),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1201),
.B(n_1093),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1199),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1233),
.A2(n_1088),
.B1(n_1041),
.B2(n_1070),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1201),
.B(n_1042),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1218),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1246),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1228),
.B(n_1096),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1248),
.B(n_1230),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1255),
.B(n_1214),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1263),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1260),
.B(n_1230),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1253),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1255),
.B(n_1269),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1272),
.B(n_1220),
.Y(n_1287)
);

NOR3xp33_ASAP7_75t_L g1288 ( 
.A(n_1261),
.B(n_1240),
.C(n_1234),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1279),
.B(n_1214),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1278),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1250),
.A2(n_1244),
.B1(n_1238),
.B2(n_1067),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1275),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_1249),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1267),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1256),
.B(n_1265),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1264),
.B(n_1206),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1277),
.B(n_1215),
.Y(n_1297)
);

AOI32xp33_ASAP7_75t_L g1298 ( 
.A1(n_1291),
.A2(n_1268),
.A3(n_1252),
.B1(n_1258),
.B2(n_1273),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1295),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_1286),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1283),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1295),
.B(n_1251),
.Y(n_1302)
);

OAI21xp33_ASAP7_75t_L g1303 ( 
.A1(n_1291),
.A2(n_1259),
.B(n_1257),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1292),
.Y(n_1304)
);

AND2x4_ASAP7_75t_SL g1305 ( 
.A(n_1296),
.B(n_1254),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1285),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1287),
.B(n_1271),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1281),
.B(n_1274),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1289),
.Y(n_1309)
);

NAND2x2_ASAP7_75t_L g1310 ( 
.A(n_1288),
.B(n_1221),
.Y(n_1310)
);

OAI21xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1282),
.A2(n_1245),
.B(n_1276),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1304),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1310),
.A2(n_1213),
.B1(n_1262),
.B2(n_1293),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1301),
.Y(n_1314)
);

AOI21xp33_ASAP7_75t_L g1315 ( 
.A1(n_1311),
.A2(n_1290),
.B(n_1294),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1307),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1311),
.A2(n_1296),
.B1(n_1264),
.B2(n_1266),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1305),
.B(n_1284),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1303),
.A2(n_1237),
.B1(n_1231),
.B2(n_1280),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1306),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1300),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1298),
.A2(n_1235),
.B(n_1270),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1309),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1323),
.B(n_1302),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1322),
.A2(n_1299),
.B1(n_1308),
.B2(n_1284),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1314),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1320),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1321),
.B(n_1297),
.Y(n_1328)
);

AOI21xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1315),
.A2(n_1222),
.B(n_1216),
.Y(n_1329)
);

OAI32xp33_ASAP7_75t_L g1330 ( 
.A1(n_1316),
.A2(n_1318),
.A3(n_1317),
.B1(n_1312),
.B2(n_1232),
.Y(n_1330)
);

AOI211xp5_ASAP7_75t_L g1331 ( 
.A1(n_1325),
.A2(n_1313),
.B(n_1319),
.C(n_1213),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1326),
.B(n_1329),
.C(n_1327),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1324),
.B(n_1178),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1328),
.B(n_1209),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1332),
.B(n_1330),
.Y(n_1335)
);

NOR2x1_ASAP7_75t_L g1336 ( 
.A(n_1333),
.B(n_1242),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1334),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1335),
.B(n_1331),
.Y(n_1338)
);

NAND4xp25_ASAP7_75t_L g1339 ( 
.A(n_1337),
.B(n_1243),
.C(n_1217),
.D(n_1215),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1336),
.B(n_1217),
.Y(n_1340)
);

NOR2x1_ASAP7_75t_L g1341 ( 
.A(n_1338),
.B(n_1204),
.Y(n_1341)
);

NOR2x1_ASAP7_75t_L g1342 ( 
.A(n_1340),
.B(n_192),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_L g1343 ( 
.A(n_1339),
.B(n_193),
.Y(n_1343)
);

NOR2x1_ASAP7_75t_L g1344 ( 
.A(n_1338),
.B(n_194),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1343),
.A2(n_1084),
.B1(n_199),
.B2(n_201),
.Y(n_1345)
);

NAND4xp25_ASAP7_75t_L g1346 ( 
.A(n_1344),
.B(n_196),
.C(n_203),
.D(n_208),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1342),
.B(n_210),
.C(n_217),
.Y(n_1347)
);

XOR2xp5_ASAP7_75t_L g1348 ( 
.A(n_1346),
.B(n_1341),
.Y(n_1348)
);

CKINVDCx6p67_ASAP7_75t_R g1349 ( 
.A(n_1347),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1349),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1348),
.Y(n_1351)
);

OAI31xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1350),
.A2(n_1345),
.A3(n_1084),
.B(n_222),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1351),
.A2(n_227),
.B1(n_229),
.B2(n_231),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1352),
.B(n_237),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1353),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_1355)
);

OAI211xp5_ASAP7_75t_L g1356 ( 
.A1(n_1354),
.A2(n_245),
.B(n_247),
.C(n_252),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1356),
.B(n_1355),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1357),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1358),
.B(n_279),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1359),
.A2(n_282),
.B1(n_285),
.B2(n_292),
.Y(n_1360)
);


endmodule