module fake_jpeg_30064_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_47),
.B1(n_35),
.B2(n_45),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_37),
.B1(n_45),
.B2(n_48),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_58),
.B1(n_69),
.B2(n_37),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_4),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_84),
.B1(n_8),
.B2(n_9),
.Y(n_89)
);

OAI22x1_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_93),
.B(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_10),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_29),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_12),
.C(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_11),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_107),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_109),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_90),
.B(n_88),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_101),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.Y(n_115)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_112),
.C(n_104),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_113),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_110),
.B(n_109),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_110),
.B(n_90),
.C(n_106),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_100),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_87),
.Y(n_122)
);


endmodule