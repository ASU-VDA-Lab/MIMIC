module fake_jpeg_16323_n_148 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_14),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_20),
.B1(n_18),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_28),
.B1(n_26),
.B2(n_14),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_66),
.B1(n_77),
.B2(n_44),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_22),
.B1(n_15),
.B2(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_78),
.B1(n_44),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_27),
.B1(n_21),
.B2(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_68),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_15),
.B(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_45),
.C(n_62),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_74),
.Y(n_91)
);

OR2x6_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_28),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_28),
.B(n_3),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_72),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_3),
.B(n_5),
.C(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_10),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_88),
.B1(n_94),
.B2(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_97),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_73),
.B(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_51),
.B1(n_78),
.B2(n_69),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_83),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_73),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_105),
.B1(n_51),
.B2(n_12),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_73),
.B(n_69),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_86),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_121),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_87),
.B(n_95),
.C(n_88),
.D(n_98),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_120),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_106),
.B1(n_105),
.B2(n_109),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_86),
.B1(n_110),
.B2(n_99),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_112),
.C(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_128),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_102),
.B(n_12),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_125),
.C(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_131),
.B1(n_135),
.B2(n_11),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_127),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_137),
.B(n_13),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_130),
.B1(n_136),
.B2(n_102),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_143),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_141),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_144),
.Y(n_148)
);


endmodule