module real_jpeg_31133_n_27 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_180, n_10, n_178, n_9, n_186, n_12, n_24, n_189, n_187, n_6, n_190, n_183, n_179, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_26, n_182, n_20, n_19, n_184, n_16, n_15, n_13, n_27);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_180;
input n_10;
input n_178;
input n_9;
input n_186;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_183;
input n_179;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_26;
input n_182;
input n_20;
input n_19;
input n_184;
input n_16;
input n_15;
input n_13;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AND2x2_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_100),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_4),
.B(n_106),
.Y(n_105)
);

HAxp5_ASAP7_75t_SL g151 ( 
.A(n_4),
.B(n_106),
.CON(n_151),
.SN(n_151)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_5),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_9),
.B(n_71),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_10),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_11),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_78),
.Y(n_170)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_14),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_15),
.A2(n_89),
.A3(n_91),
.B1(n_98),
.B2(n_154),
.C1(n_156),
.C2(n_188),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_28),
.CI(n_35),
.CON(n_27),
.SN(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_19),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_19),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_20),
.A2(n_38),
.B1(n_40),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

AOI221xp5_ASAP7_75t_L g117 ( 
.A1(n_22),
.A2(n_24),
.B1(n_118),
.B2(n_123),
.C(n_127),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_24),
.B(n_118),
.C(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_25),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_26),
.B(n_64),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_31),
.B(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_80),
.B(n_159),
.Y(n_36)
);

NAND4xp25_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_47),
.C(n_69),
.D(n_76),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_42),
.B(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_57),
.C(n_61),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_49),
.B(n_169),
.C(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_50),
.B(n_56),
.Y(n_163)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

OAI322xp33_ASAP7_75t_L g167 ( 
.A1(n_57),
.A2(n_66),
.A3(n_168),
.B1(n_171),
.B2(n_172),
.C1(n_173),
.C2(n_190),
.Y(n_167)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI321xp33_ASAP7_75t_L g161 ( 
.A1(n_62),
.A2(n_162),
.A3(n_163),
.B1(n_164),
.B2(n_167),
.C(n_189),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_70),
.A2(n_161),
.B(n_174),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI31xp67_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_111),
.A3(n_144),
.B(n_149),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_97),
.C(n_105),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_82),
.A2(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_84),
.B(n_105),
.C(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_179),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

OA21x2_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_138),
.C(n_139),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_131),
.B(n_137),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_129),
.B2(n_130),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_119),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_184),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_136),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_178),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_180),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_181),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_182),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_183),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_185),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_186),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_187),
.Y(n_147)
);


endmodule