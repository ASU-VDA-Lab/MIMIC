module fake_jpeg_12403_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_48),
.Y(n_83)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_58),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_15),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_19),
.Y(n_99)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_63),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_68),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_6),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_22),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_7),
.B1(n_12),
.B2(n_63),
.Y(n_114)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_75),
.Y(n_117)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_73),
.Y(n_110)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_79),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_19),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_40),
.B1(n_25),
.B2(n_28),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_93),
.B1(n_114),
.B2(n_86),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_40),
.B1(n_25),
.B2(n_33),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_86),
.A2(n_80),
.B1(n_56),
.B2(n_51),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_24),
.B1(n_38),
.B2(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_33),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_38),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_122),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_44),
.A2(n_39),
.B1(n_8),
.B2(n_7),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_107),
.C(n_84),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_140),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_58),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_138),
.B(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_83),
.B(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_160),
.Y(n_162)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_159),
.B1(n_84),
.B2(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_89),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_174),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_105),
.B1(n_96),
.B2(n_116),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_176),
.B1(n_161),
.B2(n_145),
.Y(n_193)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_105),
.B1(n_89),
.B2(n_119),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_169),
.A2(n_175),
.B(n_189),
.C(n_178),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_108),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_119),
.B(n_138),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_158),
.B1(n_126),
.B2(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_135),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_197),
.Y(n_214)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_183),
.B1(n_179),
.B2(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_142),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_160),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_125),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_134),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_170),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_208),
.B(n_181),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_183),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_186),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_172),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_171),
.B(n_169),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_187),
.B(n_181),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_217),
.B1(n_201),
.B2(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_203),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_169),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_205),
.C(n_209),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_222),
.B(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_195),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_232),
.C(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_203),
.C(n_192),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_192),
.C(n_208),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_212),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_235),
.B1(n_223),
.B2(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_216),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_235),
.A2(n_193),
.B1(n_219),
.B2(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_205),
.B1(n_216),
.B2(n_207),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_233),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_249),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_229),
.B1(n_205),
.B2(n_215),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_247),
.B1(n_238),
.B2(n_239),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_236),
.B1(n_238),
.B2(n_215),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_196),
.B(n_191),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_245),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_241),
.C(n_182),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_254),
.B(n_187),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

AOI31xp33_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_248),
.A3(n_246),
.B(n_184),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_188),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_188),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_258),
.A2(n_259),
.B(n_255),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_260),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_164),
.C(n_260),
.Y(n_262)
);


endmodule