module real_aes_7494_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_756;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g578 ( .A1(n_0), .A2(n_157), .B(n_579), .C(n_582), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_1), .B(n_523), .Y(n_583) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g191 ( .A(n_3), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_4), .B(n_149), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_5), .A2(n_492), .B(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_6), .A2(n_134), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_7), .A2(n_35), .B1(n_143), .B2(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_8), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_9), .B(n_134), .Y(n_160) );
AND2x6_ASAP7_75t_L g158 ( .A(n_10), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_11), .A2(n_158), .B(n_482), .C(n_484), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_36), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_12), .B(n_36), .Y(n_444) );
INVx1_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
INVx1_ASAP7_75t_L g184 ( .A(n_14), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_15), .B(n_147), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_16), .B(n_149), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_17), .B(n_135), .Y(n_196) );
AO32x2_ASAP7_75t_L g218 ( .A1(n_18), .A2(n_134), .A3(n_164), .B1(n_175), .B2(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_19), .B(n_143), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_20), .B(n_135), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_21), .A2(n_54), .B1(n_143), .B2(n_221), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g243 ( .A1(n_22), .A2(n_83), .B1(n_143), .B2(n_147), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_23), .B(n_143), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_24), .A2(n_175), .B(n_482), .C(n_543), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_25), .A2(n_175), .B(n_482), .C(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_26), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_27), .B(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_28), .A2(n_492), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_29), .B(n_177), .Y(n_215) );
INVx2_ASAP7_75t_L g145 ( .A(n_30), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_31), .A2(n_494), .B(n_502), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_32), .B(n_143), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_33), .B(n_177), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_34), .B(n_229), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_37), .B(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_38), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_39), .A2(n_79), .B1(n_459), .B2(n_460), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_39), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_40), .B(n_149), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_41), .B(n_492), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_42), .A2(n_80), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_42), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_43), .A2(n_494), .B(n_496), .C(n_502), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_44), .A2(n_458), .B1(n_461), .B2(n_462), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_44), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_45), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g580 ( .A(n_46), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_47), .A2(n_92), .B1(n_221), .B2(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g497 ( .A(n_48), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_49), .B(n_143), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_50), .B(n_143), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_51), .B(n_121), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_51), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_52), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_53), .B(n_155), .Y(n_154) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_55), .A2(n_59), .B1(n_143), .B2(n_147), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_56), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_57), .B(n_143), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_58), .B(n_143), .Y(n_226) );
INVx1_ASAP7_75t_L g159 ( .A(n_60), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_61), .B(n_492), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_62), .B(n_523), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_63), .A2(n_155), .B(n_187), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_64), .B(n_143), .Y(n_192) );
INVx1_ASAP7_75t_L g138 ( .A(n_65), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_67), .B(n_149), .Y(n_533) );
AO32x2_ASAP7_75t_L g239 ( .A1(n_68), .A2(n_134), .A3(n_175), .B1(n_240), .B2(n_244), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_69), .B(n_150), .Y(n_485) );
INVx1_ASAP7_75t_L g170 ( .A(n_70), .Y(n_170) );
INVx1_ASAP7_75t_L g210 ( .A(n_71), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g577 ( .A(n_72), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_73), .A2(n_105), .B1(n_113), .B2(n_765), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_74), .B(n_499), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_75), .A2(n_482), .B(n_502), .C(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_76), .B(n_147), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_77), .Y(n_518) );
INVx1_ASAP7_75t_L g112 ( .A(n_78), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_79), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_80), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_80), .A2(n_125), .B1(n_126), .B2(n_436), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_81), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_82), .B(n_498), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_84), .B(n_221), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_85), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_86), .B(n_147), .Y(n_214) );
INVx2_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_88), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_89), .B(n_174), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_90), .B(n_147), .Y(n_146) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_91), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g441 ( .A(n_91), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g468 ( .A(n_91), .B(n_443), .Y(n_468) );
INVx2_ASAP7_75t_L g756 ( .A(n_91), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_93), .A2(n_103), .B1(n_147), .B2(n_148), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_94), .B(n_492), .Y(n_529) );
INVx1_ASAP7_75t_L g532 ( .A(n_95), .Y(n_532) );
INVxp67_ASAP7_75t_L g521 ( .A(n_96), .Y(n_521) );
AOI222xp33_ASAP7_75t_SL g456 ( .A1(n_97), .A2(n_457), .B1(n_463), .B2(n_757), .C1(n_758), .C2(n_762), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_98), .B(n_147), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g478 ( .A(n_100), .Y(n_478) );
INVx1_ASAP7_75t_L g556 ( .A(n_101), .Y(n_556) );
AND2x2_ASAP7_75t_L g504 ( .A(n_102), .B(n_177), .Y(n_504) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g766 ( .A(n_106), .Y(n_766) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g443 ( .A(n_109), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B1(n_453), .B2(n_456), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g455 ( .A(n_117), .Y(n_455) );
AOI211xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_445), .B(n_446), .C(n_450), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_437), .C(n_440), .Y(n_119) );
INVxp67_ASAP7_75t_L g447 ( .A(n_120), .Y(n_447) );
INVx1_ASAP7_75t_L g439 ( .A(n_121), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_436), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g436 ( .A(n_126), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_360), .Y(n_126) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_128), .B(n_318), .Y(n_127) );
NOR4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_258), .C(n_294), .D(n_308), .Y(n_128) );
OAI221xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_202), .B1(n_234), .B2(n_245), .C(n_249), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_130), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_178), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_161), .Y(n_132) );
AND2x2_ASAP7_75t_L g255 ( .A(n_133), .B(n_162), .Y(n_255) );
INVx3_ASAP7_75t_L g263 ( .A(n_133), .Y(n_263) );
AND2x2_ASAP7_75t_L g317 ( .A(n_133), .B(n_181), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_133), .B(n_180), .Y(n_353) );
AND2x2_ASAP7_75t_L g411 ( .A(n_133), .B(n_273), .Y(n_411) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_160), .Y(n_133) );
INVx4_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_134), .A2(n_509), .B(n_510), .Y(n_508) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_134), .Y(n_515) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_136), .B(n_137), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_152), .B(n_158), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_149), .Y(n_141) );
INVx3_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_143), .Y(n_558) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g221 ( .A(n_144), .Y(n_221) );
BUFx3_ASAP7_75t_L g242 ( .A(n_144), .Y(n_242) );
AND2x6_ASAP7_75t_L g482 ( .A(n_144), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx2_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_149), .A2(n_167), .B(n_168), .Y(n_166) );
O2A1O1Ixp5_ASAP7_75t_SL g208 ( .A1(n_149), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_149), .B(n_521), .Y(n_520) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g240 ( .A1(n_150), .A2(n_174), .B1(n_241), .B2(n_243), .Y(n_240) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx1_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
AND2x2_ASAP7_75t_L g480 ( .A(n_151), .B(n_156), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_151), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .Y(n_152) );
INVx2_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_157), .A2(n_171), .B(n_191), .C(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_157), .A2(n_174), .B1(n_199), .B2(n_200), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_157), .A2(n_174), .B1(n_220), .B2(n_222), .Y(n_219) );
BUFx3_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_158), .A2(n_183), .B(n_190), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_158), .A2(n_208), .B(n_212), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_158), .A2(n_225), .B(n_230), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_158), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g492 ( .A(n_158), .B(n_480), .Y(n_492) );
INVx4_ASAP7_75t_SL g503 ( .A(n_158), .Y(n_503) );
AND2x2_ASAP7_75t_L g246 ( .A(n_161), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g260 ( .A(n_161), .B(n_181), .Y(n_260) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_162), .B(n_181), .Y(n_275) );
AND2x2_ASAP7_75t_L g287 ( .A(n_162), .B(n_263), .Y(n_287) );
OR2x2_ASAP7_75t_L g289 ( .A(n_162), .B(n_247), .Y(n_289) );
AND2x2_ASAP7_75t_L g324 ( .A(n_162), .B(n_247), .Y(n_324) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_162), .Y(n_369) );
INVx1_ASAP7_75t_L g377 ( .A(n_162), .Y(n_377) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_176), .Y(n_162) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_163), .A2(n_182), .B(n_193), .Y(n_181) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_164), .B(n_488), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_175), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .C(n_173), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_171), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_173), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g581 ( .A(n_174), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g197 ( .A(n_175), .B(n_198), .C(n_201), .Y(n_197) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_177), .A2(n_207), .B(n_215), .Y(n_206) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_177), .A2(n_224), .B(n_233), .Y(n_223) );
INVx2_ASAP7_75t_L g244 ( .A(n_177), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_177), .A2(n_491), .B(n_493), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_177), .A2(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g549 ( .A(n_177), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g294 ( .A1(n_178), .A2(n_295), .B1(n_299), .B2(n_303), .C(n_304), .Y(n_294) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g254 ( .A(n_179), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_194), .Y(n_179) );
INVx2_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
AND2x2_ASAP7_75t_L g306 ( .A(n_180), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g325 ( .A(n_180), .B(n_263), .Y(n_325) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g388 ( .A(n_181), .B(n_263), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .C(n_187), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_185), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_185), .A2(n_512), .B(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_187), .A2(n_556), .B(n_557), .C(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_188), .A2(n_213), .B(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g499 ( .A(n_189), .Y(n_499) );
AND2x2_ASAP7_75t_L g310 ( .A(n_194), .B(n_255), .Y(n_310) );
OAI322xp33_ASAP7_75t_L g378 ( .A1(n_194), .A2(n_334), .A3(n_379), .B1(n_381), .B2(n_384), .C1(n_386), .C2(n_390), .Y(n_378) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_195), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g274 ( .A(n_195), .Y(n_274) );
AND2x2_ASAP7_75t_L g383 ( .A(n_195), .B(n_263), .Y(n_383) );
AND2x2_ASAP7_75t_L g415 ( .A(n_195), .B(n_287), .Y(n_415) );
OR2x2_ASAP7_75t_L g418 ( .A(n_195), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
AO21x1_ASAP7_75t_L g247 ( .A1(n_198), .A2(n_201), .B(n_248), .Y(n_247) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_201), .A2(n_477), .B(n_487), .Y(n_476) );
INVx3_ASAP7_75t_L g523 ( .A(n_201), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_201), .B(n_535), .Y(n_534) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_201), .A2(n_553), .B(n_560), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_201), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_216), .Y(n_203) );
INVx1_ASAP7_75t_L g431 ( .A(n_204), .Y(n_431) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g236 ( .A(n_205), .B(n_223), .Y(n_236) );
INVx2_ASAP7_75t_L g271 ( .A(n_205), .Y(n_271) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g293 ( .A(n_206), .Y(n_293) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_206), .Y(n_301) );
OR2x2_ASAP7_75t_L g425 ( .A(n_206), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g250 ( .A(n_216), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g290 ( .A(n_216), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g342 ( .A(n_216), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
AND2x2_ASAP7_75t_L g237 ( .A(n_217), .B(n_238), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_217), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g351 ( .A(n_217), .B(n_239), .Y(n_351) );
OR2x2_ASAP7_75t_L g359 ( .A(n_217), .B(n_293), .Y(n_359) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g268 ( .A(n_218), .Y(n_268) );
AND2x2_ASAP7_75t_L g278 ( .A(n_218), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g302 ( .A(n_218), .B(n_223), .Y(n_302) );
AND2x2_ASAP7_75t_L g366 ( .A(n_218), .B(n_239), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_223), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_223), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
INVx1_ASAP7_75t_L g284 ( .A(n_223), .Y(n_284) );
AND2x2_ASAP7_75t_L g296 ( .A(n_223), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_223), .Y(n_374) );
INVx1_ASAP7_75t_L g426 ( .A(n_223), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g403 ( .A(n_235), .B(n_312), .Y(n_403) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g330 ( .A(n_237), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g429 ( .A(n_237), .B(n_364), .Y(n_429) );
INVx1_ASAP7_75t_L g251 ( .A(n_238), .Y(n_251) );
AND2x2_ASAP7_75t_L g277 ( .A(n_238), .B(n_271), .Y(n_277) );
BUFx2_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_239), .Y(n_257) );
INVx1_ASAP7_75t_L g267 ( .A(n_239), .Y(n_267) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_242), .Y(n_501) );
INVx2_ASAP7_75t_L g582 ( .A(n_242), .Y(n_582) );
INVx1_ASAP7_75t_L g546 ( .A(n_244), .Y(n_546) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_245), .B(n_252), .Y(n_405) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI32xp33_ASAP7_75t_L g249 ( .A1(n_246), .A2(n_250), .A3(n_252), .B1(n_254), .B2(n_256), .Y(n_249) );
AND2x2_ASAP7_75t_L g389 ( .A(n_246), .B(n_262), .Y(n_389) );
AND2x2_ASAP7_75t_L g427 ( .A(n_246), .B(n_325), .Y(n_427) );
INVx1_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_251), .B(n_313), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_252), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_252), .B(n_255), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_252), .B(n_324), .Y(n_406) );
OR2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_289), .Y(n_420) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g347 ( .A(n_253), .B(n_255), .Y(n_347) );
OR2x2_ASAP7_75t_L g356 ( .A(n_253), .B(n_343), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_255), .B(n_306), .Y(n_328) );
INVx2_ASAP7_75t_L g343 ( .A(n_257), .Y(n_343) );
OR2x2_ASAP7_75t_L g358 ( .A(n_257), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_374), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_257), .A2(n_350), .B(n_431), .C(n_432), .Y(n_430) );
OAI321xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .A3(n_269), .B1(n_272), .B2(n_276), .C(n_280), .Y(n_258) );
INVx1_ASAP7_75t_L g371 ( .A(n_259), .Y(n_371) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g382 ( .A(n_260), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_263), .B(n_377), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_264), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x2_ASAP7_75t_L g339 ( .A(n_266), .B(n_313), .Y(n_339) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_267), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_269), .A2(n_310), .B(n_355), .C(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g321 ( .A(n_271), .B(n_278), .Y(n_321) );
BUFx2_ASAP7_75t_L g331 ( .A(n_271), .Y(n_331) );
INVx1_ASAP7_75t_L g346 ( .A(n_271), .Y(n_346) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OR2x2_ASAP7_75t_L g352 ( .A(n_274), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g435 ( .A(n_274), .Y(n_435) );
INVx1_ASAP7_75t_L g428 ( .A(n_275), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_277), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g385 ( .A(n_277), .B(n_302), .Y(n_385) );
INVx1_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .B1(n_288), .B2(n_290), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_282), .B(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g350 ( .A(n_283), .B(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_284), .B(n_293), .Y(n_313) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_292), .A2(n_410), .B1(n_412), .B2(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g298 ( .A(n_293), .Y(n_298) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_293), .Y(n_364) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_296), .B(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_297), .A2(n_302), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_300), .B(n_310), .Y(n_407) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g376 ( .A(n_301), .Y(n_376) );
AND2x2_ASAP7_75t_L g335 ( .A(n_302), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
INVx1_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
INVx1_ASAP7_75t_L g395 ( .A(n_306), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B1(n_314), .B2(n_315), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_312), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g380 ( .A(n_313), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_313), .B(n_351), .Y(n_417) );
OR2x2_ASAP7_75t_L g390 ( .A(n_314), .B(n_343), .Y(n_390) );
INVx1_ASAP7_75t_L g329 ( .A(n_315), .Y(n_329) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_317), .B(n_368), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_337), .C(n_348), .Y(n_318) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_322), .B(n_326), .C(n_332), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_321), .A2(n_392), .B1(n_396), .B2(n_399), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g333 ( .A(n_324), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g387 ( .A(n_324), .B(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_325), .A2(n_373), .B(n_375), .C(n_377), .Y(n_372) );
INVx2_ASAP7_75t_L g419 ( .A(n_325), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_329), .B(n_330), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g398 ( .A(n_331), .B(n_351), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
OAI21xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_341), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI21xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_347), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_342), .B(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_347), .B(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B(n_354), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g375 ( .A(n_351), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND4x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_391), .C(n_408), .D(n_430), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_378), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_367), .B(n_370), .C(n_372), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_366), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_377), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g412 ( .A(n_387), .Y(n_412) );
INVx2_ASAP7_75t_SL g400 ( .A(n_388), .Y(n_400) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_416), .Y(n_408) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_421), .C(n_422), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g448 ( .A(n_437), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g449 ( .A(n_441), .Y(n_449) );
BUFx2_ASAP7_75t_L g451 ( .A(n_441), .Y(n_451) );
NOR2x2_ASAP7_75t_L g764 ( .A(n_442), .B(n_756), .Y(n_764) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g755 ( .A(n_443), .B(n_756), .Y(n_755) );
AOI211xp5_ASAP7_75t_L g446 ( .A1(n_445), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_450), .B(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g757 ( .A(n_457), .Y(n_757) );
INVx1_ASAP7_75t_L g461 ( .A(n_458), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_466), .B1(n_469), .B2(n_753), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_465), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g759 ( .A(n_467), .Y(n_759) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g760 ( .A(n_469), .Y(n_760) );
OR3x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_651), .C(n_716), .Y(n_469) );
NAND4xp25_ASAP7_75t_SL g470 ( .A(n_471), .B(n_592), .C(n_618), .D(n_641), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_524), .B1(n_562), .B2(n_569), .C(n_584), .Y(n_471) );
CKINVDCx14_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_473), .A2(n_585), .B1(n_609), .B2(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_505), .Y(n_473) );
INVx1_ASAP7_75t_SL g645 ( .A(n_474), .Y(n_645) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_489), .Y(n_474) );
OR2x2_ASAP7_75t_L g567 ( .A(n_475), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g587 ( .A(n_475), .B(n_506), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_475), .B(n_514), .Y(n_600) );
AND2x2_ASAP7_75t_L g617 ( .A(n_475), .B(n_489), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_475), .B(n_565), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_475), .B(n_616), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_475), .B(n_505), .Y(n_738) );
AOI211xp5_ASAP7_75t_SL g749 ( .A1(n_475), .A2(n_655), .B(n_750), .C(n_751), .Y(n_749) );
INVx5_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_476), .B(n_506), .Y(n_621) );
AND2x2_ASAP7_75t_L g624 ( .A(n_476), .B(n_507), .Y(n_624) );
OR2x2_ASAP7_75t_L g669 ( .A(n_476), .B(n_506), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_476), .B(n_514), .Y(n_678) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_481), .Y(n_477) );
INVx5_ASAP7_75t_L g495 ( .A(n_482), .Y(n_495) );
INVx5_ASAP7_75t_SL g568 ( .A(n_489), .Y(n_568) );
AND2x2_ASAP7_75t_L g586 ( .A(n_489), .B(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_489), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g672 ( .A(n_489), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g704 ( .A(n_489), .B(n_514), .Y(n_704) );
OR2x2_ASAP7_75t_L g710 ( .A(n_489), .B(n_600), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_489), .B(n_660), .Y(n_719) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_504), .Y(n_489) );
BUFx2_ASAP7_75t_L g541 ( .A(n_492), .Y(n_541) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_495), .A2(n_503), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g576 ( .A1(n_495), .A2(n_503), .B(n_577), .C(n_578), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_500), .C(n_501), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_498), .A2(n_501), .B(n_532), .C(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
AND2x2_ASAP7_75t_L g601 ( .A(n_506), .B(n_568), .Y(n_601) );
INVx1_ASAP7_75t_SL g614 ( .A(n_506), .Y(n_614) );
OR2x2_ASAP7_75t_L g649 ( .A(n_506), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g655 ( .A(n_506), .B(n_514), .Y(n_655) );
AND2x2_ASAP7_75t_L g713 ( .A(n_506), .B(n_565), .Y(n_713) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_507), .B(n_568), .Y(n_640) );
INVx3_ASAP7_75t_L g565 ( .A(n_514), .Y(n_565) );
OR2x2_ASAP7_75t_L g606 ( .A(n_514), .B(n_568), .Y(n_606) );
AND2x2_ASAP7_75t_L g616 ( .A(n_514), .B(n_614), .Y(n_616) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_514), .Y(n_664) );
AND2x2_ASAP7_75t_L g673 ( .A(n_514), .B(n_587), .Y(n_673) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_522), .Y(n_514) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_523), .A2(n_575), .B(n_583), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_524), .A2(n_690), .B1(n_692), .B2(n_694), .C(n_697), .Y(n_689) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_536), .Y(n_525) );
AND2x2_ASAP7_75t_L g663 ( .A(n_526), .B(n_644), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_526), .B(n_722), .Y(n_726) );
OR2x2_ASAP7_75t_L g747 ( .A(n_526), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_526), .B(n_752), .Y(n_751) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx5_ASAP7_75t_L g594 ( .A(n_527), .Y(n_594) );
AND2x2_ASAP7_75t_L g671 ( .A(n_527), .B(n_538), .Y(n_671) );
AND2x2_ASAP7_75t_L g732 ( .A(n_527), .B(n_611), .Y(n_732) );
AND2x2_ASAP7_75t_L g745 ( .A(n_527), .B(n_565), .Y(n_745) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_550), .Y(n_536) );
AND2x4_ASAP7_75t_L g572 ( .A(n_537), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g590 ( .A(n_537), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g597 ( .A(n_537), .Y(n_597) );
AND2x2_ASAP7_75t_L g666 ( .A(n_537), .B(n_644), .Y(n_666) );
AND2x2_ASAP7_75t_L g676 ( .A(n_537), .B(n_594), .Y(n_676) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_537), .Y(n_684) );
AND2x2_ASAP7_75t_L g696 ( .A(n_537), .B(n_574), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_537), .B(n_628), .Y(n_700) );
AND2x2_ASAP7_75t_L g737 ( .A(n_537), .B(n_732), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_537), .B(n_611), .Y(n_748) );
OR2x2_ASAP7_75t_L g750 ( .A(n_537), .B(n_686), .Y(n_750) );
INVx5_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g636 ( .A(n_538), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_538), .B(n_591), .Y(n_646) );
AND2x2_ASAP7_75t_L g658 ( .A(n_538), .B(n_574), .Y(n_658) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_538), .Y(n_688) );
AND2x4_ASAP7_75t_L g722 ( .A(n_538), .B(n_573), .Y(n_722) );
OR2x6_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .Y(n_538) );
AOI21xp5_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_542), .B(n_546), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
BUFx2_ASAP7_75t_L g571 ( .A(n_550), .Y(n_571) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
AND2x2_ASAP7_75t_L g644 ( .A(n_551), .B(n_574), .Y(n_644) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g591 ( .A(n_552), .B(n_574), .Y(n_591) );
BUFx2_ASAP7_75t_L g637 ( .A(n_552), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_564), .B(n_645), .Y(n_724) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_565), .B(n_587), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_565), .B(n_568), .Y(n_626) );
AND2x2_ASAP7_75t_L g681 ( .A(n_565), .B(n_617), .Y(n_681) );
AOI221xp5_ASAP7_75t_SL g618 ( .A1(n_566), .A2(n_619), .B1(n_627), .B2(n_629), .C(n_633), .Y(n_618) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g613 ( .A(n_567), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g654 ( .A(n_567), .B(n_655), .Y(n_654) );
OAI321xp33_ASAP7_75t_L g661 ( .A1(n_567), .A2(n_620), .A3(n_662), .B1(n_664), .B2(n_665), .C(n_667), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_568), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_571), .B(n_722), .Y(n_740) );
AND2x2_ASAP7_75t_L g627 ( .A(n_572), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_572), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_573), .Y(n_603) );
AND2x2_ASAP7_75t_L g610 ( .A(n_573), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_573), .B(n_685), .Y(n_715) );
INVx1_ASAP7_75t_L g752 ( .A(n_573), .Y(n_752) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B(n_589), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_586), .A2(n_696), .B(n_745), .C(n_746), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_587), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_587), .B(n_625), .Y(n_691) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g634 ( .A(n_591), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_591), .B(n_594), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_591), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_591), .B(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_607), .B2(n_612), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g608 ( .A(n_594), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g631 ( .A(n_594), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g643 ( .A(n_594), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_594), .B(n_637), .Y(n_679) );
OR2x2_ASAP7_75t_L g686 ( .A(n_594), .B(n_611), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_594), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g736 ( .A(n_594), .B(n_722), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B1(n_602), .B2(n_604), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g642 ( .A(n_597), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_600), .A2(n_615), .B1(n_683), .B2(n_687), .Y(n_682) );
INVx1_ASAP7_75t_L g730 ( .A(n_601), .Y(n_730) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_605), .A2(n_642), .B1(n_645), .B2(n_646), .C(n_647), .Y(n_641) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g620 ( .A(n_606), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_610), .B(n_676), .Y(n_708) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_611), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_611), .Y(n_632) );
NAND2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g650 ( .A(n_617), .Y(n_650) );
AND2x2_ASAP7_75t_L g659 ( .A(n_617), .B(n_660), .Y(n_659) );
NAND2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g703 ( .A(n_624), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_627), .A2(n_653), .B1(n_656), .B2(n_659), .C(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_631), .B(n_688), .Y(n_687) );
AOI21xp33_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_635), .B(n_638), .Y(n_633) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_638), .Y(n_735) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g677 ( .A(n_640), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g698 ( .A(n_643), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_643), .B(n_703), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_646), .B(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_670), .C(n_689), .D(n_702), .Y(n_651) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g660 ( .A(n_655), .Y(n_660) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g693 ( .A(n_664), .B(n_669), .Y(n_693) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_674), .C(n_682), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_672), .A2(n_714), .B(n_742), .C(n_749), .Y(n_741) );
INVx1_ASAP7_75t_SL g701 ( .A(n_673), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_674) );
INVx1_ASAP7_75t_L g705 ( .A(n_679), .Y(n_705) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_685), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_685), .B(n_696), .Y(n_729) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g706 ( .A(n_696), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B(n_701), .Y(n_697) );
INVxp33_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .A3(n_706), .B1(n_707), .B2(n_709), .C1(n_711), .C2(n_714), .Y(n_702) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND3xp33_ASAP7_75t_SL g716 ( .A(n_717), .B(n_734), .C(n_741), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g733 ( .A(n_722), .Y(n_733) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_737), .B2(n_738), .C(n_739), .Y(n_734) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVxp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g761 ( .A(n_754), .Y(n_761) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
endmodule