module fake_jpeg_17664_n_351 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_49),
.B1(n_30),
.B2(n_32),
.Y(n_87)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_22),
.B1(n_49),
.B2(n_48),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_16),
.C(n_18),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_16),
.C(n_18),
.Y(n_99)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_22),
.B1(n_34),
.B2(n_19),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_73),
.B1(n_31),
.B2(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_34),
.B1(n_31),
.B2(n_35),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_78),
.Y(n_118)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_97),
.B1(n_109),
.B2(n_55),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_27),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_27),
.B(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_79),
.B(n_86),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_87),
.B1(n_110),
.B2(n_55),
.Y(n_129)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_88),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_89),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_46),
.B1(n_50),
.B2(n_47),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_138)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_42),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_58),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_18),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_46),
.B1(n_50),
.B2(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_54),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_18),
.B(n_16),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_18),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_28),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_127),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_55),
.B(n_41),
.C(n_42),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_137),
.B(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_125),
.B(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_88),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_94),
.B1(n_106),
.B2(n_77),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_90),
.B(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_94),
.A3(n_80),
.B1(n_98),
.B2(n_102),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_151),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_149),
.B1(n_162),
.B2(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_84),
.B1(n_91),
.B2(n_81),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_150),
.B1(n_171),
.B2(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_81),
.B1(n_66),
.B2(n_104),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_74),
.B1(n_107),
.B2(n_96),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_33),
.C(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_92),
.C(n_103),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_164),
.C(n_167),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_119),
.B(n_37),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_117),
.B(n_28),
.Y(n_193)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_100),
.C(n_37),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_33),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_21),
.B(n_20),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_114),
.A2(n_75),
.B1(n_97),
.B2(n_89),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_44),
.C(n_41),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_173),
.C(n_28),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_37),
.C(n_76),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_147),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_127),
.B(n_141),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_193),
.B(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_120),
.B1(n_112),
.B2(n_133),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_136),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_120),
.B1(n_136),
.B2(n_123),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_112),
.B1(n_133),
.B2(n_111),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_131),
.B1(n_111),
.B2(n_125),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_194),
.B1(n_196),
.B2(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_17),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_173),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_111),
.B1(n_124),
.B2(n_126),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_184),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_126),
.B1(n_25),
.B2(n_33),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_25),
.B1(n_20),
.B2(n_17),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_25),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_148),
.B(n_21),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_151),
.B(n_15),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_3),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_150),
.A2(n_20),
.B1(n_17),
.B2(n_21),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_14),
.B1(n_13),
.B2(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_208),
.A2(n_215),
.B1(n_219),
.B2(n_224),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_162),
.C(n_171),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_214),
.C(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_152),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_229),
.Y(n_247)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_177),
.B(n_161),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_188),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_154),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_145),
.B1(n_163),
.B2(n_142),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_3),
.B(n_4),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_0),
.B(n_1),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_231),
.B(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_182),
.B(n_21),
.CI(n_13),
.CON(n_229),
.SN(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_146),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_186),
.C(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_SL g235 ( 
.A(n_178),
.B(n_1),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_207),
.B1(n_181),
.B2(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_241),
.B(n_256),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_195),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_243),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_185),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_245),
.C(n_248),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_212),
.C(n_233),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_194),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_251),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_196),
.C(n_198),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_193),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_204),
.C(n_179),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_258),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_260),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_205),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_204),
.C(n_187),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_235),
.C(n_237),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_262),
.A2(n_211),
.B1(n_227),
.B2(n_209),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_211),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_281),
.B1(n_200),
.B2(n_261),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_181),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_259),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_274),
.B(n_280),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_217),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_247),
.B(n_225),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_226),
.B1(n_209),
.B2(n_218),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_226),
.B1(n_220),
.B2(n_190),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_175),
.B1(n_187),
.B2(n_208),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_208),
.B1(n_229),
.B2(n_200),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_241),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_246),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_290),
.C(n_295),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_240),
.CI(n_238),
.CON(n_289),
.SN(n_289)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_245),
.C(n_239),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_239),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_297),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_292),
.A2(n_294),
.B1(n_281),
.B2(n_279),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_242),
.CI(n_229),
.CON(n_293),
.SN(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_206),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_200),
.C(n_6),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_302),
.C(n_267),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_5),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_5),
.C(n_6),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_311),
.B1(n_294),
.B2(n_302),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_314),
.C(n_316),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_268),
.B(n_271),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_308),
.A2(n_7),
.B(n_8),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_310),
.B(n_289),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_286),
.B(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_315),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_270),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_272),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_272),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_268),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_300),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_327),
.C(n_316),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_291),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_325),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_324),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_296),
.B1(n_299),
.B2(n_293),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_307),
.B1(n_303),
.B2(n_325),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_293),
.B1(n_289),
.B2(n_290),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_7),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_304),
.B(n_10),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_306),
.Y(n_331)
);

AOI211xp5_ASAP7_75t_L g340 ( 
.A1(n_331),
.A2(n_326),
.B(n_321),
.C(n_327),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_333),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_306),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_319),
.A2(n_314),
.B(n_10),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_8),
.B(n_10),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_318),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_329),
.Y(n_343)
);

OAI211xp5_ASAP7_75t_L g344 ( 
.A1(n_339),
.A2(n_340),
.B(n_334),
.C(n_332),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_344),
.B(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_333),
.Y(n_345)
);

NAND4xp25_ASAP7_75t_SL g347 ( 
.A(n_346),
.B(n_337),
.C(n_342),
.D(n_338),
.Y(n_347)
);

AOI21x1_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_336),
.B(n_320),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_336),
.B(n_10),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_8),
.B(n_11),
.Y(n_350)
);

AOI221xp5_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_11),
.B1(n_12),
.B2(n_330),
.C(n_256),
.Y(n_351)
);


endmodule