module real_aes_10718_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_917;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_922;
wire n_679;
wire n_926;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_0), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_1), .B(n_155), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_2), .A2(n_82), .B1(n_593), .B2(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_3), .B(n_171), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_4), .B(n_166), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_5), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_6), .A2(n_37), .B1(n_145), .B2(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g104 ( .A(n_7), .Y(n_104) );
NOR2xp67_ASAP7_75t_L g119 ( .A(n_7), .B(n_84), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_8), .B(n_147), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_9), .B(n_128), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_10), .A2(n_62), .B1(n_145), .B2(n_250), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_11), .B(n_145), .C(n_148), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_12), .B(n_128), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_13), .B(n_168), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_14), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_15), .B(n_567), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_16), .B(n_135), .Y(n_580) );
AND2x2_ASAP7_75t_L g249 ( .A(n_17), .B(n_250), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_18), .B(n_141), .C(n_147), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_19), .A2(n_27), .B1(n_147), .B2(n_610), .Y(n_631) );
INVx1_ASAP7_75t_L g931 ( .A(n_20), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_21), .B(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_22), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_23), .B(n_176), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_24), .B(n_154), .Y(n_239) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_25), .B(n_184), .Y(n_183) );
NAND2xp33_ASAP7_75t_L g207 ( .A(n_26), .B(n_184), .Y(n_207) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_29), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_30), .B(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_31), .A2(n_51), .B1(n_184), .B2(n_250), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_32), .B(n_141), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_33), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g109 ( .A(n_34), .Y(n_109) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_35), .A2(n_65), .B(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_36), .A2(n_140), .B(n_255), .C(n_256), .Y(n_254) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_38), .B(n_165), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_39), .B(n_145), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_40), .Y(n_279) );
AND2x6_ASAP7_75t_L g151 ( .A(n_41), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g647 ( .A(n_42), .B(n_176), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_43), .B(n_176), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_44), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_45), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_46), .B(n_206), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g238 ( .A(n_47), .B(n_165), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_48), .B(n_135), .Y(n_569) );
INVx1_ASAP7_75t_L g152 ( .A(n_49), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_50), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_52), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_53), .B(n_176), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_54), .B(n_147), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_55), .A2(n_552), .B1(n_916), .B2(n_917), .Y(n_551) );
INVx1_ASAP7_75t_L g916 ( .A(n_55), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_55), .A2(n_916), .B1(n_919), .B2(n_921), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_56), .Y(n_275) );
AND2x2_ASAP7_75t_L g107 ( .A(n_57), .B(n_108), .Y(n_107) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_58), .B(n_176), .Y(n_574) );
AND2x2_ASAP7_75t_L g258 ( .A(n_59), .B(n_154), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_60), .B(n_147), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_61), .B(n_148), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_63), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_64), .B(n_654), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_66), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_67), .Y(n_657) );
NAND2xp33_ASAP7_75t_L g134 ( .A(n_68), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_69), .B(n_148), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_70), .A2(n_74), .B1(n_147), .B2(n_610), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_71), .B(n_171), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_72), .Y(n_602) );
BUFx10_ASAP7_75t_L g542 ( .A(n_73), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_75), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_SL g635 ( .A(n_76), .Y(n_635) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_77), .B(n_147), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_78), .A2(n_121), .B1(n_531), .B2(n_532), .Y(n_120) );
INVx1_ASAP7_75t_L g531 ( .A(n_78), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_79), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_80), .B(n_184), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_81), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_83), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_84), .B(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_86), .B(n_148), .Y(n_625) );
INVx1_ASAP7_75t_L g110 ( .A(n_87), .Y(n_110) );
OR2x2_ASAP7_75t_L g116 ( .A(n_87), .B(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g550 ( .A(n_87), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_87), .B(n_118), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_88), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_89), .B(n_165), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_90), .B(n_190), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_91), .B(n_176), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_92), .Y(n_233) );
INVx1_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
INVx1_ASAP7_75t_L g248 ( .A(n_94), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_95), .Y(n_219) );
AND2x2_ASAP7_75t_L g228 ( .A(n_96), .B(n_128), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_97), .B(n_226), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_98), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_111), .B(n_930), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx6_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g933 ( .A(n_102), .Y(n_933) );
AND2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .C(n_110), .Y(n_105) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g118 ( .A(n_109), .B(n_119), .Y(n_118) );
OR2x6_ASAP7_75t_L g111 ( .A(n_112), .B(n_534), .Y(n_111) );
OAI21xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_537), .B(n_543), .Y(n_112) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_120), .B(n_533), .Y(n_113) );
INVx5_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_116), .Y(n_536) );
AND2x2_ASAP7_75t_L g549 ( .A(n_117), .B(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g923 ( .A(n_117), .B(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g532 ( .A(n_121), .Y(n_532) );
INVx2_ASAP7_75t_L g920 ( .A(n_121), .Y(n_920) );
AND3x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_390), .C(n_481), .Y(n_121) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_123), .B(n_343), .Y(n_122) );
NAND3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_301), .C(n_325), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_193), .B1(n_264), .B2(n_266), .Y(n_124) );
AND2x2_ASAP7_75t_L g447 ( .A(n_125), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_156), .Y(n_125) );
OR2x6_ASAP7_75t_SL g483 ( .A(n_126), .B(n_352), .Y(n_483) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_127), .Y(n_327) );
INVx2_ASAP7_75t_L g359 ( .A(n_127), .Y(n_359) );
AND2x2_ASAP7_75t_L g506 ( .A(n_127), .B(n_383), .Y(n_506) );
NAND2x1_ASAP7_75t_L g514 ( .A(n_127), .B(n_347), .Y(n_514) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_153), .Y(n_127) );
INVx3_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
INVx4_ASAP7_75t_L g213 ( .A(n_128), .Y(n_213) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_128), .A2(n_132), .B(n_153), .Y(n_285) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_128), .A2(n_132), .B(n_153), .Y(n_295) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_128), .Y(n_705) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_129), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g155 ( .A(n_130), .Y(n_155) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_142), .B(n_149), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B(n_139), .Y(n_133) );
INVx2_ASAP7_75t_L g138 ( .A(n_135), .Y(n_138) );
INVx2_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
INVx1_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
INVx1_ASAP7_75t_L g571 ( .A(n_135), .Y(n_571) );
INVx2_ASAP7_75t_L g593 ( .A(n_135), .Y(n_593) );
INVx2_ASAP7_75t_L g600 ( .A(n_135), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_135), .B(n_602), .Y(n_601) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_136), .Y(n_145) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
INVx2_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_136), .Y(n_226) );
INVx1_ASAP7_75t_L g252 ( .A(n_136), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_139), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_139), .A2(n_237), .B(n_238), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_139), .A2(n_203), .B1(n_609), .B2(n_611), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_139), .A2(n_191), .B1(n_631), .B2(n_632), .Y(n_630) );
OA22x2_ASAP7_75t_L g643 ( .A1(n_139), .A2(n_191), .B1(n_644), .B2(n_645), .Y(n_643) );
CKINVDCx6p67_ASAP7_75t_R g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_SL g220 ( .A(n_140), .Y(n_220) );
AOI21x1_ASAP7_75t_L g564 ( .A1(n_140), .A2(n_565), .B(n_566), .Y(n_564) );
AOI21x1_ASAP7_75t_L g579 ( .A1(n_140), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_140), .A2(n_596), .B(n_601), .Y(n_595) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
BUFx12f_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_141), .A2(n_275), .B(n_276), .C(n_277), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_141), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_582) );
OAI321xp33_ASAP7_75t_L g590 ( .A1(n_141), .A2(n_147), .A3(n_591), .B1(n_592), .B2(n_593), .C(n_594), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_148), .Y(n_142) );
NOR2xp67_ASAP7_75t_L g218 ( .A(n_144), .B(n_219), .Y(n_218) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
INVx2_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
INVx2_ASAP7_75t_SL g206 ( .A(n_147), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_147), .B(n_217), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_147), .A2(n_148), .B(n_657), .C(n_658), .Y(n_656) );
AOI21x1_ASAP7_75t_L g163 ( .A1(n_148), .A2(n_164), .B(n_167), .Y(n_163) );
INVx1_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
OAI21x1_ASAP7_75t_L g180 ( .A1(n_149), .A2(n_181), .B(n_185), .Y(n_180) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_149), .A2(n_199), .B(n_204), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_149), .A2(n_232), .B(n_236), .Y(n_231) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_149), .A2(n_274), .B(n_278), .Y(n_273) );
AND2x2_ASAP7_75t_L g607 ( .A(n_149), .B(n_161), .Y(n_607) );
AO31x2_ASAP7_75t_L g629 ( .A1(n_149), .A2(n_213), .A3(n_630), .B(n_634), .Y(n_629) );
INVx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_150), .A2(n_215), .B(n_221), .Y(n_214) );
NOR2xp67_ASAP7_75t_L g243 ( .A(n_150), .B(n_244), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_150), .A2(n_594), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g642 ( .A(n_150), .Y(n_642) );
INVx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx2_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_151), .A2(n_579), .B(n_582), .Y(n_578) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_151), .A2(n_620), .B(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g664 ( .A(n_151), .Y(n_664) );
INVx2_ASAP7_75t_L g641 ( .A(n_154), .Y(n_641) );
BUFx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_155), .Y(n_604) );
INVx1_ASAP7_75t_L g614 ( .A(n_155), .Y(n_614) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_178), .Y(n_156) );
INVx2_ASAP7_75t_L g300 ( .A(n_157), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_157), .B(n_315), .Y(n_384) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g329 ( .A(n_158), .B(n_317), .Y(n_329) );
AND2x2_ASAP7_75t_L g339 ( .A(n_158), .B(n_316), .Y(n_339) );
OR2x2_ASAP7_75t_L g352 ( .A(n_158), .B(n_305), .Y(n_352) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_175), .Y(n_159) );
OAI21x1_ASAP7_75t_L g197 ( .A1(n_160), .A2(n_198), .B(n_209), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_160), .A2(n_162), .B(n_175), .Y(n_306) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_160), .A2(n_619), .B(n_627), .Y(n_618) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_160), .A2(n_619), .B(n_627), .Y(n_693) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_169), .B(n_174), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_165), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
INVx1_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
INVx1_ASAP7_75t_L g234 ( .A(n_168), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_173), .Y(n_169) );
INVx3_ASAP7_75t_L g191 ( .A(n_173), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_173), .Y(n_203) );
BUFx2_ASAP7_75t_L g253 ( .A(n_173), .Y(n_253) );
AOI21x1_ASAP7_75t_L g568 ( .A1(n_173), .A2(n_569), .B(n_570), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_173), .A2(n_660), .B(n_661), .Y(n_659) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_174), .A2(n_564), .B(n_568), .Y(n_563) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g286 ( .A(n_178), .Y(n_286) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_192), .Y(n_178) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_179), .A2(n_231), .B(n_239), .Y(n_230) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_179), .A2(n_273), .B(n_281), .Y(n_272) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_179), .A2(n_273), .B(n_281), .Y(n_305) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_179), .A2(n_180), .B(n_192), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_184), .B(n_257), .Y(n_256) );
O2A1O1Ixp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .C(n_191), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_187), .A2(n_191), .B(n_279), .C(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_191), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_259), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_210), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_195), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_195), .B(n_260), .Y(n_511) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g389 ( .A(n_196), .B(n_290), .Y(n_389) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g263 ( .A(n_197), .B(n_229), .Y(n_263) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_197), .Y(n_291) );
INVx1_ASAP7_75t_L g297 ( .A(n_197), .Y(n_297) );
INVx1_ASAP7_75t_L g337 ( .A(n_197), .Y(n_337) );
AND2x2_ASAP7_75t_L g398 ( .A(n_197), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g474 ( .A(n_197), .B(n_261), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_203), .Y(n_199) );
INVx1_ASAP7_75t_L g276 ( .A(n_202), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g221 ( .A1(n_203), .A2(n_222), .B(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B(n_208), .Y(n_204) );
INVx2_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
INVx1_ASAP7_75t_L g475 ( .A(n_210), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_240), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_229), .Y(n_211) );
INVx2_ASAP7_75t_SL g311 ( .A(n_212), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_212), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g364 ( .A(n_212), .Y(n_364) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_228), .Y(n_212) );
INVx3_ASAP7_75t_L g244 ( .A(n_213), .Y(n_244) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_213), .A2(n_214), .B(n_228), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_218), .B(n_220), .Y(n_215) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_225), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g567 ( .A(n_226), .Y(n_567) );
INVx2_ASAP7_75t_L g610 ( .A(n_226), .Y(n_610) );
INVx2_ASAP7_75t_L g662 ( .A(n_226), .Y(n_662) );
OR2x2_ASAP7_75t_L g296 ( .A(n_229), .B(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g333 ( .A(n_229), .Y(n_333) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g290 ( .A(n_230), .Y(n_290) );
AND2x2_ASAP7_75t_L g499 ( .A(n_230), .B(n_261), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_240), .B(n_290), .Y(n_492) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g265 ( .A(n_241), .Y(n_265) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_241), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_241), .B(n_290), .Y(n_438) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B(n_258), .Y(n_242) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_244), .A2(n_563), .B(n_574), .Y(n_562) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_244), .A2(n_578), .B(n_586), .Y(n_577) );
OAI21x1_ASAP7_75t_L g676 ( .A1(n_244), .A2(n_563), .B(n_574), .Y(n_676) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_244), .A2(n_578), .B(n_586), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_253), .Y(n_246) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g633 ( .A(n_252), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_255), .A2(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx2_ASAP7_75t_L g407 ( .A(n_260), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_260), .B(n_333), .Y(n_427) );
AND2x2_ASAP7_75t_L g440 ( .A(n_260), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_L g331 ( .A(n_261), .B(n_324), .Y(n_331) );
INVx1_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
AND2x2_ASAP7_75t_L g375 ( .A(n_262), .B(n_311), .Y(n_375) );
INVx1_ASAP7_75t_L g399 ( .A(n_262), .Y(n_399) );
AND2x2_ASAP7_75t_L g307 ( .A(n_263), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_263), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g374 ( .A(n_263), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_263), .B(n_401), .Y(n_400) );
NAND2xp67_ASAP7_75t_L g419 ( .A(n_263), .B(n_331), .Y(n_419) );
OR2x2_ASAP7_75t_L g356 ( .A(n_264), .B(n_296), .Y(n_356) );
OR2x2_ASAP7_75t_L g468 ( .A(n_264), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g381 ( .A(n_265), .B(n_335), .Y(n_381) );
OR2x2_ASAP7_75t_L g473 ( .A(n_265), .B(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_287), .B1(n_292), .B2(n_298), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_282), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g299 ( .A(n_270), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g328 ( .A(n_270), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g360 ( .A(n_270), .B(n_339), .Y(n_360) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g342 ( .A(n_272), .Y(n_342) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_272), .Y(n_434) );
AND2x2_ASAP7_75t_L g430 ( .A(n_282), .B(n_341), .Y(n_430) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_283), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g314 ( .A(n_285), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g354 ( .A(n_285), .B(n_315), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_285), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_286), .B(n_342), .Y(n_372) );
INVx1_ASAP7_75t_L g464 ( .A(n_286), .Y(n_464) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g406 ( .A(n_289), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g414 ( .A(n_290), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_290), .B(n_364), .Y(n_522) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
OR2x2_ASAP7_75t_L g421 ( .A(n_293), .B(n_352), .Y(n_421) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g320 ( .A(n_294), .B(n_315), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_294), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g369 ( .A(n_295), .Y(n_369) );
INVx1_ASAP7_75t_L g424 ( .A(n_295), .Y(n_424) );
INVx1_ASAP7_75t_SL g496 ( .A(n_295), .Y(n_496) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_296), .Y(n_378) );
INVx1_ASAP7_75t_SL g449 ( .A(n_296), .Y(n_449) );
INVx1_ASAP7_75t_L g508 ( .A(n_296), .Y(n_508) );
OAI322xp33_ASAP7_75t_L g512 ( .A1(n_298), .A2(n_478), .A3(n_513), .B1(n_514), .B2(n_515), .C1(n_517), .C2(n_521), .Y(n_512) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
AND2x4_ASAP7_75t_SL g454 ( .A(n_300), .B(n_342), .Y(n_454) );
AOI32xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_307), .A3(n_312), .B1(n_318), .B2(n_321), .Y(n_301) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_302), .B(n_478), .C(n_480), .Y(n_477) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_303), .A2(n_417), .B(n_487), .C(n_490), .Y(n_486) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g319 ( .A(n_304), .Y(n_319) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g349 ( .A(n_305), .B(n_315), .Y(n_349) );
INVx1_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
BUFx2_ASAP7_75t_L g466 ( .A(n_306), .Y(n_466) );
INVx1_ASAP7_75t_L g501 ( .A(n_308), .Y(n_501) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g411 ( .A(n_314), .B(n_341), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_314), .A2(n_381), .B1(n_452), .B2(n_455), .Y(n_451) );
NOR2xp33_ASAP7_75t_R g476 ( .A(n_314), .B(n_352), .Y(n_476) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2x1_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g497 ( .A(n_319), .Y(n_497) );
OR2x2_ASAP7_75t_L g432 ( .A(n_320), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g513 ( .A(n_323), .B(n_474), .Y(n_513) );
AND2x2_ASAP7_75t_L g528 ( .A(n_323), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_330), .B1(n_334), .B2(n_338), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_329), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g520 ( .A(n_329), .Y(n_520) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g409 ( .A(n_333), .B(n_375), .Y(n_409) );
AND2x2_ASAP7_75t_L g479 ( .A(n_333), .B(n_359), .Y(n_479) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g437 ( .A(n_336), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g491 ( .A(n_336), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g442 ( .A(n_337), .Y(n_442) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g367 ( .A(n_339), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g426 ( .A(n_339), .Y(n_426) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g444 ( .A(n_342), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_376), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_355), .B(n_357), .C(n_365), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_346), .A2(n_380), .B1(n_382), .B2(n_388), .Y(n_379) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g405 ( .A(n_353), .Y(n_405) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g445 ( .A(n_354), .Y(n_445) );
INVx1_ASAP7_75t_L g505 ( .A(n_354), .Y(n_505) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_356), .B(n_396), .C(n_400), .Y(n_395) );
OAI311xp33_ASAP7_75t_L g500 ( .A1(n_356), .A2(n_460), .A3(n_501), .B1(n_502), .C1(n_509), .Y(n_500) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
AOI21xp33_ASAP7_75t_SL g376 ( .A1(n_358), .A2(n_377), .B(n_379), .Y(n_376) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_359), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_359), .B(n_519), .Y(n_526) );
INVx3_ASAP7_75t_L g525 ( .A(n_360), .Y(n_525) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g397 ( .A(n_364), .B(n_398), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B(n_373), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g423 ( .A(n_372), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g448 ( .A(n_375), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g457 ( .A(n_375), .B(n_442), .Y(n_457) );
INVx1_ASAP7_75t_L g480 ( .A(n_375), .Y(n_480) );
INVxp33_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_385), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g518 ( .A(n_385), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g394 ( .A(n_387), .Y(n_394) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g469 ( .A(n_389), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_428), .C(n_450), .Y(n_390) );
NAND3xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_403), .C(n_412), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_393), .A2(n_472), .B1(n_494), .B2(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g413 ( .A(n_397), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g489 ( .A(n_398), .Y(n_489) );
AND2x4_ASAP7_75t_L g498 ( .A(n_398), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g485 ( .A(n_400), .Y(n_485) );
AND2x2_ASAP7_75t_L g507 ( .A(n_401), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_408), .B2(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI221x1_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_418), .B2(n_420), .C(n_422), .Y(n_412) );
AND2x4_ASAP7_75t_L g529 ( .A(n_414), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_419), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B(n_427), .Y(n_422) );
OR2x2_ASAP7_75t_L g425 ( .A(n_424), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g471 ( .A(n_425), .Y(n_471) );
BUFx2_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_435), .B(n_439), .C(n_446), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_432), .A2(n_524), .B(n_527), .Y(n_523) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_434), .Y(n_504) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g461 ( .A(n_437), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_458), .C(n_470), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B1(n_462), .B2(n_467), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_475), .B2(n_476), .C(n_477), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_474), .Y(n_516) );
INVx2_ASAP7_75t_L g530 ( .A(n_474), .Y(n_530) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_500), .C(n_512), .D(n_523), .Y(n_481) );
OAI211xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_484), .B(n_486), .C(n_493), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_506), .B(n_507), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g921 ( .A(n_532), .Y(n_921) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g928 ( .A(n_541), .B(n_929), .Y(n_928) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
INVx6_ASAP7_75t_L g548 ( .A(n_542), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_551), .B1(n_918), .B2(n_922), .C(n_925), .Y(n_543) );
INVx4_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_SL g922 ( .A(n_547), .B(n_923), .Y(n_922) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_550), .Y(n_924) );
INVx1_ASAP7_75t_L g917 ( .A(n_552), .Y(n_917) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR3x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_793), .C(n_888), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_736), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_682), .C(n_715), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_615), .B1(n_636), .B2(n_665), .C(n_669), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_587), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_559), .B(n_792), .Y(n_849) );
INVx2_ASAP7_75t_SL g860 ( .A(n_559), .Y(n_860) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_575), .Y(n_559) );
INVx1_ASAP7_75t_L g718 ( .A(n_560), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_560), .B(n_575), .Y(n_768) );
AND2x2_ASAP7_75t_L g862 ( .A(n_560), .B(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g765 ( .A(n_561), .B(n_605), .Y(n_765) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_561), .Y(n_788) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g686 ( .A(n_562), .Y(n_686) );
INVxp67_ASAP7_75t_L g622 ( .A(n_567), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g584 ( .A(n_571), .Y(n_584) );
INVx4_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g754 ( .A(n_576), .Y(n_754) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g750 ( .A(n_577), .Y(n_750) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g713 ( .A(n_588), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g734 ( .A(n_588), .B(n_735), .Y(n_734) );
BUFx3_ASAP7_75t_L g757 ( .A(n_588), .Y(n_757) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_605), .Y(n_588) );
INVx2_ASAP7_75t_L g668 ( .A(n_589), .Y(n_668) );
INVx1_ASAP7_75t_L g678 ( .A(n_589), .Y(n_678) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .B(n_603), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g688 ( .A(n_605), .Y(n_688) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g667 ( .A(n_606), .Y(n_667) );
AOI21x1_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_612), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_614), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g654 ( .A(n_614), .Y(n_654) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_628), .Y(n_616) );
INVx2_ASAP7_75t_L g731 ( .A(n_617), .Y(n_731) );
NOR2xp67_ASAP7_75t_L g839 ( .A(n_617), .B(n_840), .Y(n_839) );
NAND2xp33_ASAP7_75t_SL g882 ( .A(n_617), .B(n_806), .Y(n_882) );
BUFx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g650 ( .A(n_618), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g725 ( .A(n_618), .B(n_652), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_623), .Y(n_620) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_628), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g872 ( .A(n_628), .Y(n_872) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_628), .Y(n_896) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g694 ( .A(n_629), .Y(n_694) );
INVx1_ASAP7_75t_L g722 ( .A(n_629), .Y(n_722) );
AND2x2_ASAP7_75t_L g730 ( .A(n_629), .B(n_704), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_629), .B(n_639), .Y(n_807) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_629), .Y(n_886) );
OAI22xp33_ASAP7_75t_SL g890 ( .A1(n_636), .A2(n_891), .B1(n_892), .B2(n_893), .Y(n_890) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_648), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_637), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g759 ( .A(n_637), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g870 ( .A(n_637), .Y(n_870) );
AND2x2_ASAP7_75t_L g915 ( .A(n_637), .B(n_769), .Y(n_915) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g778 ( .A(n_638), .B(n_769), .Y(n_778) );
AND2x2_ASAP7_75t_L g850 ( .A(n_638), .B(n_851), .Y(n_850) );
NOR2x1_ASAP7_75t_L g864 ( .A(n_638), .B(n_721), .Y(n_864) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g681 ( .A(n_639), .Y(n_681) );
INVx1_ASAP7_75t_L g712 ( .A(n_639), .Y(n_712) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_639), .Y(n_727) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_639), .Y(n_914) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_646), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
OA21x2_ASAP7_75t_L g704 ( .A1(n_643), .A2(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g706 ( .A(n_647), .Y(n_706) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g680 ( .A(n_650), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g771 ( .A(n_650), .Y(n_771) );
INVx2_ASAP7_75t_L g703 ( .A(n_651), .Y(n_703) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g711 ( .A(n_652), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
OAI21x1_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B(n_663), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_665), .B(n_870), .C(n_871), .Y(n_869) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g717 ( .A(n_666), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g747 ( .A(n_666), .B(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_666), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g842 ( .A(n_666), .B(n_674), .Y(n_842) );
OR2x2_ASAP7_75t_L g868 ( .A(n_666), .B(n_768), .Y(n_868) );
NOR2xp67_ASAP7_75t_L g887 ( .A(n_666), .B(n_735), .Y(n_887) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AND2x2_ASAP7_75t_L g677 ( .A(n_667), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_667), .B(n_714), .Y(n_775) );
AND2x2_ASAP7_75t_L g697 ( .A(n_668), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g814 ( .A(n_668), .B(n_699), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_679), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_672), .B(n_677), .Y(n_671) );
OR2x2_ASAP7_75t_L g881 ( .A(n_672), .B(n_775), .Y(n_881) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g818 ( .A(n_673), .B(n_754), .Y(n_818) );
AND2x2_ASAP7_75t_L g854 ( .A(n_673), .B(n_697), .Y(n_854) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g700 ( .A(n_674), .B(n_687), .Y(n_700) );
AND2x2_ASAP7_75t_L g826 ( .A(n_674), .B(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g834 ( .A(n_674), .B(n_761), .Y(n_834) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_674), .Y(n_847) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g753 ( .A(n_675), .B(n_688), .Y(n_753) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g800 ( .A(n_676), .B(n_678), .Y(n_800) );
AND2x2_ASAP7_75t_L g763 ( .A(n_677), .B(n_749), .Y(n_763) );
INVx2_ASAP7_75t_L g792 ( .A(n_677), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_677), .B(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g832 ( .A(n_678), .Y(n_832) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g742 ( .A(n_681), .Y(n_742) );
AND2x2_ASAP7_75t_L g905 ( .A(n_681), .B(n_710), .Y(n_905) );
AOI322xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_689), .A3(n_695), .B1(n_700), .B2(n_701), .C1(n_707), .C2(n_713), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_684), .A2(n_909), .B(n_911), .C(n_915), .Y(n_908) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI32xp33_ASAP7_75t_L g883 ( .A1(n_685), .A2(n_813), .A3(n_851), .B1(n_884), .B2(n_887), .Y(n_883) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
BUFx2_ASAP7_75t_L g733 ( .A(n_686), .Y(n_733) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_686), .Y(n_756) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_688), .Y(n_799) );
NOR2x1p5_ASAP7_75t_L g809 ( .A(n_690), .B(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g701 ( .A(n_691), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
AND2x2_ASAP7_75t_L g761 ( .A(n_692), .B(n_703), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_692), .B(n_711), .Y(n_824) );
INVx1_ASAP7_75t_L g863 ( .A(n_692), .Y(n_863) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g785 ( .A(n_693), .B(n_704), .Y(n_785) );
AND2x4_ASAP7_75t_L g710 ( .A(n_694), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g841 ( .A(n_694), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_695), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_696), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g714 ( .A(n_699), .Y(n_714) );
INVx1_ASAP7_75t_L g815 ( .A(n_700), .Y(n_815) );
AND2x4_ASAP7_75t_L g892 ( .A(n_700), .B(n_754), .Y(n_892) );
INVx2_ASAP7_75t_L g816 ( .A(n_702), .Y(n_816) );
AND2x4_ASAP7_75t_L g838 ( .A(n_702), .B(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g769 ( .A(n_703), .B(n_722), .Y(n_769) );
INVx2_ASAP7_75t_L g784 ( .A(n_703), .Y(n_784) );
INVx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_708), .A2(n_836), .B1(n_837), .B2(n_842), .Y(n_835) );
OR2x6_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g743 ( .A(n_710), .B(n_731), .Y(n_743) );
INVx1_ASAP7_75t_L g819 ( .A(n_710), .Y(n_819) );
AND2x2_ASAP7_75t_L g851 ( .A(n_711), .B(n_841), .Y(n_851) );
AND2x2_ASAP7_75t_L g811 ( .A(n_712), .B(n_784), .Y(n_811) );
AND2x2_ASAP7_75t_L g879 ( .A(n_712), .B(n_725), .Y(n_879) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_713), .Y(n_779) );
INVx2_ASAP7_75t_L g735 ( .A(n_714), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B1(n_728), .B2(n_732), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_718), .B(n_814), .Y(n_836) );
AOI221xp5_ASAP7_75t_SL g772 ( .A1(n_719), .A2(n_773), .B1(n_776), .B2(n_779), .C(n_780), .Y(n_772) );
AND2x4_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp67_ASAP7_75t_L g783 ( .A(n_722), .B(n_784), .Y(n_783) );
BUFx2_ASAP7_75t_L g853 ( .A(n_723), .Y(n_853) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g776 ( .A(n_724), .B(n_759), .C(n_777), .Y(n_776) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx2_ASAP7_75t_L g805 ( .A(n_725), .Y(n_805) );
AND2x2_ASAP7_75t_L g884 ( .A(n_725), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
AND2x4_ASAP7_75t_L g831 ( .A(n_735), .B(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_772), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_744), .B(n_758), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2x1p5_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_740), .A2(n_821), .B(n_835), .Y(n_820) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g790 ( .A(n_742), .B(n_761), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_751), .C(n_755), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_748), .Y(n_910) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g848 ( .A(n_750), .B(n_832), .Y(n_848) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g893 ( .A(n_752), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx2_ASAP7_75t_L g878 ( .A(n_753), .Y(n_878) );
AND2x2_ASAP7_75t_L g795 ( .A(n_754), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g901 ( .A(n_754), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B(n_766), .Y(n_758) );
INVx2_ASAP7_75t_L g875 ( .A(n_760), .Y(n_875) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_763), .A2(n_767), .B1(n_769), .B2(n_770), .Y(n_766) );
INVx2_ASAP7_75t_L g796 ( .A(n_765), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_765), .A2(n_898), .B1(n_903), .B2(n_906), .C(n_908), .Y(n_897) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g827 ( .A(n_775), .Y(n_827) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_786), .B1(n_789), .B2(n_791), .Y(n_780) );
INVx1_ASAP7_75t_L g891 ( .A(n_781), .Y(n_891) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_785), .Y(n_782) );
INVx1_ASAP7_75t_L g859 ( .A(n_784), .Y(n_859) );
AND2x4_ASAP7_75t_L g865 ( .A(n_785), .B(n_851), .Y(n_865) );
OR2x2_ASAP7_75t_L g791 ( .A(n_787), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g797 ( .A(n_789), .Y(n_797) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g895 ( .A(n_790), .B(n_896), .Y(n_895) );
NAND4xp75_ASAP7_75t_L g793 ( .A(n_794), .B(n_820), .C(n_843), .D(n_866), .Y(n_793) );
AOI221x1_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_797), .B1(n_798), .B2(n_801), .C(n_812), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_798), .B(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_808), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_806), .B(n_859), .Y(n_858) );
AND2x2_ASAP7_75t_L g899 ( .A(n_806), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_807), .B(n_824), .Y(n_902) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI32xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_815), .A3(n_816), .B1(n_817), .B2(n_819), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_L g861 ( .A1(n_814), .A2(n_862), .B(n_864), .C(n_865), .Y(n_861) );
AND2x2_ASAP7_75t_L g876 ( .A(n_814), .B(n_877), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_825), .B1(n_828), .B2(n_833), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx4_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_831), .Y(n_907) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVxp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_842), .A2(n_881), .B(n_882), .C(n_883), .Y(n_880) );
NOR2xp67_ASAP7_75t_L g843 ( .A(n_844), .B(n_855), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_852), .Y(n_844) );
OAI21xp33_ASAP7_75t_SL g845 ( .A1(n_846), .A2(n_849), .B(n_850), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_856), .B(n_861), .Y(n_855) );
NAND2x1_ASAP7_75t_SL g856 ( .A(n_857), .B(n_860), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g900 ( .A(n_859), .Y(n_900) );
AND2x2_ASAP7_75t_L g904 ( .A(n_862), .B(n_905), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_863), .B(n_914), .Y(n_913) );
AOI221x1_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_873), .B1(n_876), .B2(n_879), .C(n_880), .Y(n_866) );
NAND2xp5_ASAP7_75t_SL g867 ( .A(n_868), .B(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OR2x2_ASAP7_75t_L g912 ( .A(n_872), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OR2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_897), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_894), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_901), .B(n_902), .Y(n_898) );
INVxp67_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVxp67_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
BUFx12f_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
NOR2xp33_ASAP7_75t_SL g930 ( .A(n_931), .B(n_932), .Y(n_930) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
endmodule