module fake_netlist_6_3578_n_1919 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1919);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1919;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_166;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_37),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_38),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_40),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_1),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_31),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_85),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_26),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_21),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_28),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_77),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_95),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_70),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_29),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_26),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_63),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_42),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_15),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_49),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_81),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_4),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_28),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_100),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_48),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_33),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_102),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_29),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_69),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_37),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_10),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_78),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_33),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_123),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_17),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_115),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_134),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_1),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_66),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_147),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_18),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_68),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_46),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_11),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_11),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_133),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_31),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_21),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_34),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_49),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_74),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_24),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_22),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_67),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_35),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_16),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_104),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_62),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_86),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_34),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_108),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_79),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_65),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_57),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_150),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_30),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_8),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_148),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_46),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_130),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_110),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_20),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_64),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_41),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_59),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_54),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_45),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_141),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_103),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_6),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_106),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_44),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_20),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_87),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_76),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_136),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_105),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_139),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_38),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_90),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_35),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_89),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_60),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_113),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_30),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_52),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_109),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_75),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_127),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_72),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_56),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_94),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_39),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_220),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_197),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_194),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_197),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_197),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_201),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_197),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_197),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_159),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_197),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_162),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_162),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_170),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_294),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_177),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_312),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_220),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_181),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_165),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_302),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_171),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_178),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_244),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_161),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_244),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_171),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_264),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_188),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_188),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_183),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_193),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_193),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_214),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_214),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_218),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_235),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_264),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_235),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_243),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_185),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_243),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_249),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_171),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_186),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_198),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_249),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_205),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_184),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_286),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_286),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_184),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_288),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_315),
.A2(n_242),
.B(n_179),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_304),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_324),
.B(n_184),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_314),
.A2(n_349),
.B1(n_351),
.B2(n_355),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_329),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_351),
.A2(n_307),
.B1(n_180),
.B2(n_196),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_331),
.B(n_191),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_356),
.B(n_191),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_381),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_319),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_335),
.A2(n_158),
.B1(n_257),
.B2(n_281),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_357),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_358),
.A2(n_296),
.B1(n_217),
.B2(n_306),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_317),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_352),
.A2(n_236),
.B1(n_221),
.B2(n_223),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_353),
.B(n_191),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_361),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_R g419 ( 
.A(n_364),
.B(n_207),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_316),
.A2(n_237),
.B1(n_206),
.B2(n_204),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_321),
.B(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_325),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_242),
.B(n_179),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_378),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_325),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_282),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_320),
.B(n_160),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_326),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_283),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_326),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_338),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_327),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_282),
.Y(n_441)
);

BUFx12f_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_328),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_332),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_321),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_328),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_342),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_332),
.B(n_282),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_334),
.B(n_283),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_330),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_334),
.B(n_255),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_435),
.B(n_379),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_419),
.B(n_380),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_420),
.A2(n_232),
.B1(n_274),
.B2(n_273),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_421),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_396),
.B(n_343),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_418),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_398),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_402),
.B(n_304),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_457),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_417),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_445),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_413),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_399),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_336),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_337),
.C(n_336),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_421),
.B(n_187),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_426),
.B(n_337),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_420),
.A2(n_272),
.B1(n_271),
.B2(n_270),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_458),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_426),
.B(n_215),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_340),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_416),
.B(n_234),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_416),
.B(n_277),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_428),
.B(n_285),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_394),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_429),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_394),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_429),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_437),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_445),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_L g516 ( 
.A1(n_409),
.A2(n_163),
.B1(n_247),
.B2(n_246),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_429),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_429),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_428),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_433),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_404),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_433),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_453),
.B(n_340),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_SL g531 ( 
.A(n_414),
.B(n_405),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_404),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_403),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_409),
.B(n_187),
.Y(n_540)
);

AND3x2_ASAP7_75t_L g541 ( 
.A(n_447),
.B(n_295),
.C(n_255),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_407),
.A2(n_397),
.B1(n_400),
.B2(n_231),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_451),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_431),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_422),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_447),
.A2(n_241),
.B1(n_239),
.B2(n_238),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_403),
.B(n_453),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_452),
.B(n_304),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_R g554 ( 
.A(n_453),
.B(n_164),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_422),
.Y(n_555)
);

OAI21xp33_ASAP7_75t_SL g556 ( 
.A1(n_455),
.A2(n_344),
.B(n_341),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_403),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_431),
.B(n_161),
.Y(n_558)
);

AND3x4_ASAP7_75t_L g559 ( 
.A(n_453),
.B(n_295),
.C(n_173),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_403),
.B(n_341),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_392),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_430),
.B(n_345),
.C(n_344),
.Y(n_562)
);

INVxp33_ASAP7_75t_SL g563 ( 
.A(n_400),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_430),
.B(n_345),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_393),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_393),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_411),
.B(n_346),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_399),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_411),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_432),
.B(n_346),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_411),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_432),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_438),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_434),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_442),
.B(n_187),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_434),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_442),
.B(n_187),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_438),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_399),
.Y(n_581)
);

AND3x2_ASAP7_75t_L g582 ( 
.A(n_448),
.B(n_169),
.C(n_168),
.Y(n_582)
);

BUFx6f_ASAP7_75t_SL g583 ( 
.A(n_448),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_399),
.B(n_347),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_450),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_450),
.B(n_347),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_390),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_401),
.B(n_348),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_395),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_390),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_401),
.A2(n_169),
.B(n_168),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_454),
.A2(n_167),
.B1(n_260),
.B2(n_259),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_434),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_401),
.B(n_348),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_434),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_434),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_408),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_436),
.Y(n_601)
);

AND2x2_ASAP7_75t_SL g602 ( 
.A(n_436),
.B(n_304),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_395),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_436),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_436),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_408),
.B(n_210),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_436),
.B(n_211),
.Y(n_607)
);

BUFx6f_ASAP7_75t_SL g608 ( 
.A(n_391),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_465),
.B(n_363),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_480),
.B(n_436),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_475),
.B(n_363),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_511),
.Y(n_612)
);

AO22x2_ASAP7_75t_L g613 ( 
.A1(n_559),
.A2(n_203),
.B1(n_209),
.B2(n_212),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_557),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_515),
.B(n_365),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_525),
.B(n_535),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_365),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_551),
.A2(n_519),
.B1(n_539),
.B2(n_557),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_439),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_591),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_463),
.B(n_366),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_602),
.B(n_519),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_496),
.B(n_366),
.Y(n_625)
);

AO22x2_ASAP7_75t_L g626 ( 
.A1(n_559),
.A2(n_203),
.B1(n_209),
.B2(n_212),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_525),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_597),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_497),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_535),
.B(n_367),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_539),
.B(n_367),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_574),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_549),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_495),
.B(n_176),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_575),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_555),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_585),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_512),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_585),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_586),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_586),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_580),
.B(n_182),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_588),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_476),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_588),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_512),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_565),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_565),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_584),
.Y(n_652)
);

BUFx8_ASAP7_75t_L g653 ( 
.A(n_583),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_512),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_512),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

OAI221xp5_ASAP7_75t_L g657 ( 
.A1(n_556),
.A2(n_267),
.B1(n_189),
.B2(n_175),
.C(n_174),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_190),
.Y(n_658)
);

OR2x2_ASAP7_75t_SL g659 ( 
.A(n_498),
.B(n_172),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_496),
.A2(n_229),
.B1(n_213),
.B2(n_216),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_523),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_512),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_540),
.B(n_192),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_561),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_513),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_554),
.Y(n_667)
);

OAI221xp5_ASAP7_75t_L g668 ( 
.A1(n_556),
.A2(n_311),
.B1(n_174),
.B2(n_175),
.C(n_189),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_549),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_560),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_513),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_569),
.B(n_439),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_511),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_502),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_569),
.B(n_439),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_529),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_564),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_566),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_566),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_567),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_368),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_504),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_504),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_368),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_545),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

NAND3x1_ASAP7_75t_L g691 ( 
.A(n_544),
.B(n_240),
.C(n_172),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_513),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_513),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_509),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_592),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_536),
.B(n_219),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_549),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_590),
.B(n_304),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_545),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_532),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_572),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_514),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_514),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_520),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_483),
.B(n_544),
.C(n_490),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_568),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_571),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_550),
.B(n_369),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_483),
.B(n_369),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_520),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_571),
.B(n_439),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_573),
.B(n_439),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_522),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_589),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_549),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_522),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_524),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_549),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_524),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_592),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_573),
.B(n_439),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_602),
.A2(n_478),
.B1(n_460),
.B2(n_526),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_526),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_530),
.B(n_443),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_532),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_530),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_462),
.A2(n_219),
.B1(n_225),
.B2(n_240),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_583),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_534),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_534),
.B(n_443),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_538),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_570),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_471),
.Y(n_733)
);

AOI22x1_ASAP7_75t_L g734 ( 
.A1(n_590),
.A2(n_593),
.B1(n_547),
.B2(n_538),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_594),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_547),
.B(n_443),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_459),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_487),
.B(n_195),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_531),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_473),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_443),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_461),
.B(n_370),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_570),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_473),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_600),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_516),
.B(n_284),
.C(n_248),
.Y(n_746)
);

CKINVDCx8_ASAP7_75t_R g747 ( 
.A(n_546),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_563),
.A2(n_225),
.B1(n_250),
.B2(n_256),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_558),
.B(n_250),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_563),
.A2(n_256),
.B1(n_261),
.B2(n_262),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_558),
.B(n_370),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_600),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_SL g754 ( 
.A(n_583),
.B(n_261),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_594),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_562),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_546),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_536),
.Y(n_758)
);

OAI221xp5_ASAP7_75t_L g759 ( 
.A1(n_562),
.A2(n_262),
.B1(n_267),
.B2(n_290),
.C(n_297),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_473),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_459),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_558),
.B(n_371),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_606),
.B(n_443),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_466),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_558),
.B(n_290),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_466),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_558),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_570),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

NOR2x1p5_ASAP7_75t_L g770 ( 
.A(n_577),
.B(n_199),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_471),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_536),
.B(n_222),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_581),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_581),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_533),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_533),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_541),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_537),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_536),
.B(n_297),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_537),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_607),
.A2(n_226),
.B1(n_224),
.B2(n_230),
.Y(n_781)
);

AOI211xp5_ASAP7_75t_L g782 ( 
.A1(n_664),
.A2(n_527),
.B(n_521),
.C(n_595),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_667),
.B(n_579),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_703),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_647),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_647),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_747),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_703),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_630),
.A2(n_468),
.B1(n_482),
.B2(n_484),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_663),
.B(n_464),
.Y(n_790)
);

AND2x6_ASAP7_75t_SL g791 ( 
.A(n_664),
.B(n_749),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_611),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_630),
.B(n_464),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_710),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_615),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_641),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_667),
.B(n_470),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_616),
.B(n_582),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_641),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_609),
.B(n_471),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_705),
.A2(n_481),
.B1(n_503),
.B2(n_470),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_663),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_707),
.B(n_481),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_624),
.B(n_471),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_758),
.A2(n_593),
.B(n_471),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_707),
.B(n_482),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_710),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_701),
.B(n_714),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_624),
.B(n_471),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_621),
.B(n_484),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_719),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_756),
.A2(n_503),
.B1(n_501),
.B2(n_499),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_672),
.B(n_489),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_637),
.A2(n_499),
.B1(n_494),
.B2(n_493),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_757),
.B(n_303),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_719),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_637),
.A2(n_309),
.B(n_311),
.C(n_303),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_726),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_672),
.B(n_489),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_752),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_756),
.A2(n_552),
.B(n_309),
.C(n_543),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_R g822 ( 
.A(n_754),
.B(n_608),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_738),
.A2(n_658),
.B(n_645),
.C(n_628),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_726),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_612),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_616),
.B(n_603),
.Y(n_826)
);

NOR2x2_ASAP7_75t_L g827 ( 
.A(n_749),
.B(n_765),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_746),
.B(n_200),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_729),
.Y(n_829)
);

INVx5_ASAP7_75t_L g830 ( 
.A(n_641),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_758),
.B(n_245),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_758),
.B(n_251),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_652),
.A2(n_492),
.B1(n_494),
.B2(n_493),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_701),
.B(n_492),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_618),
.B(n_371),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_623),
.A2(n_501),
.B1(n_469),
.B2(n_510),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_722),
.A2(n_598),
.B1(n_605),
.B2(n_604),
.Y(n_837)
);

NOR2x1_ASAP7_75t_R g838 ( 
.A(n_675),
.B(n_202),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_641),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_729),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_627),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_619),
.A2(n_598),
.B1(n_605),
.B2(n_604),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_714),
.B(n_542),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_689),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_706),
.B(n_542),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_645),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_631),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_706),
.B(n_543),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_737),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_699),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_649),
.B(n_548),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_650),
.A2(n_576),
.B1(n_578),
.B2(n_601),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_657),
.A2(n_548),
.B(n_553),
.C(n_601),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_737),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_622),
.B(n_373),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_649),
.B(n_553),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_757),
.Y(n_857)
);

OR2x2_ASAP7_75t_SL g858 ( 
.A(n_728),
.B(n_373),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_649),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_649),
.B(n_576),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_629),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_631),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_658),
.B(n_625),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_654),
.B(n_578),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_676),
.A2(n_599),
.B1(n_596),
.B2(n_587),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_633),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_758),
.B(n_252),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_SL g868 ( 
.A1(n_738),
.A2(n_608),
.B1(n_292),
.B2(n_287),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_654),
.B(n_587),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_633),
.B(n_603),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_757),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_629),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_676),
.A2(n_614),
.B1(n_617),
.B2(n_742),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_639),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_708),
.B(n_208),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_639),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_775),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_654),
.B(n_596),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_654),
.B(n_599),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_655),
.B(n_666),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_655),
.B(n_469),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_739),
.B(n_228),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_745),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_753),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_651),
.B(n_233),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_656),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_775),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_627),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_653),
.Y(n_889)
);

INVx5_ASAP7_75t_L g890 ( 
.A(n_655),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_655),
.B(n_603),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_653),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_665),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_666),
.B(n_472),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_666),
.B(n_673),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_666),
.B(n_673),
.Y(n_896)
);

NAND2xp33_ASAP7_75t_SL g897 ( 
.A(n_770),
.B(n_608),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_671),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_673),
.B(n_472),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_754),
.B(n_266),
.C(n_258),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_673),
.B(n_254),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_683),
.B(n_474),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_683),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_776),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_679),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_777),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_683),
.B(n_269),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_SL g908 ( 
.A(n_657),
.B(n_268),
.C(n_265),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_749),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_683),
.B(n_474),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_692),
.B(n_477),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_765),
.Y(n_912)
);

NAND2x1_ASAP7_75t_L g913 ( 
.A(n_692),
.B(n_467),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_776),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_762),
.B(n_467),
.Y(n_915)
);

BUFx8_ASAP7_75t_L g916 ( 
.A(n_767),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_692),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_692),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_685),
.B(n_374),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_732),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_680),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_693),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_681),
.Y(n_923)
);

NOR2x2_ASAP7_75t_L g924 ( 
.A(n_765),
.B(n_454),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_682),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_632),
.A2(n_518),
.B(n_517),
.C(n_510),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_732),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_763),
.A2(n_485),
.B(n_473),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_661),
.B(n_467),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_685),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_688),
.B(n_374),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_623),
.A2(n_505),
.B1(n_507),
.B2(n_508),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_688),
.A2(n_505),
.B1(n_507),
.B2(n_508),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_659),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_693),
.B(n_275),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_693),
.B(n_279),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_693),
.B(n_634),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_695),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_740),
.Y(n_939)
);

NOR2x1_ASAP7_75t_R g940 ( 
.A(n_709),
.B(n_280),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_781),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_691),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_709),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_635),
.B(n_289),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_638),
.B(n_491),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_613),
.B(n_376),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_640),
.B(n_642),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_695),
.B(n_376),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_643),
.B(n_477),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_644),
.B(n_486),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_646),
.B(n_491),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_648),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_686),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_687),
.B(n_690),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_684),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_743),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_694),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_748),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_727),
.A2(n_518),
.B1(n_517),
.B2(n_506),
.Y(n_959)
);

BUFx4f_ASAP7_75t_SL g960 ( 
.A(n_720),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_702),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_704),
.B(n_291),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_613),
.B(n_377),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_720),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_713),
.B(n_491),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_716),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_717),
.B(n_500),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_620),
.A2(n_479),
.B(n_473),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_613),
.B(n_377),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_723),
.B(n_486),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_731),
.B(n_506),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_743),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_768),
.B(n_293),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_735),
.B(n_750),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_796),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_943),
.B(n_769),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_784),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_798),
.B(n_773),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_788),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_825),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_863),
.B(n_610),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_798),
.B(n_774),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_824),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_823),
.B(n_696),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_802),
.B(n_735),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_846),
.B(n_696),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_794),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_796),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_830),
.B(n_890),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_871),
.B(n_636),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_875),
.B(n_668),
.C(n_772),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_877),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_887),
.Y(n_993)
);

OR2x4_ASAP7_75t_L g994 ( 
.A(n_808),
.B(n_626),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_904),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_830),
.B(n_779),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_947),
.A2(n_668),
.B(n_698),
.C(n_759),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_844),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_807),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_796),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_903),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_793),
.B(n_835),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_787),
.B(n_759),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_850),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_914),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_841),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_930),
.B(n_761),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_960),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_841),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_903),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_855),
.B(n_750),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_845),
.A2(n_698),
.B(n_741),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_843),
.B(n_755),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_792),
.B(n_755),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_817),
.A2(n_730),
.B(n_724),
.C(n_736),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_786),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_843),
.B(n_727),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_785),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_888),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_834),
.B(n_727),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_903),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_811),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_849),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_816),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_834),
.B(n_626),
.Y(n_1025)
);

INVx3_ASAP7_75t_SL g1026 ( 
.A(n_857),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_917),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_964),
.B(n_974),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_974),
.B(n_626),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_797),
.B(n_764),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_947),
.B(n_954),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_889),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_880),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_820),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_917),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_954),
.B(n_766),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_818),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_795),
.B(n_778),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_906),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_958),
.B(n_780),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_917),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_919),
.B(n_748),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_942),
.B(n_660),
.Y(n_1043)
);

AND2x6_ASAP7_75t_SL g1044 ( 
.A(n_815),
.B(n_382),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_830),
.B(n_890),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_845),
.A2(n_712),
.B(n_721),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_813),
.B(n_748),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_946),
.A2(n_751),
.B1(n_734),
.B2(n_772),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_819),
.B(n_751),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_830),
.B(n_890),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_931),
.B(n_751),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_941),
.A2(n_388),
.B1(n_386),
.B2(n_385),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_886),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_854),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_861),
.Y(n_1055)
);

BUFx8_ASAP7_75t_L g1056 ( 
.A(n_892),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_882),
.B(n_382),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_885),
.B(n_948),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_948),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_938),
.B(n_847),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_888),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_893),
.Y(n_1062)
);

CKINVDCx11_ASAP7_75t_R g1063 ( 
.A(n_934),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_862),
.B(n_385),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_938),
.B(n_636),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_898),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_905),
.B(n_674),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_921),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_938),
.B(n_669),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_953),
.B(n_662),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_874),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_873),
.B(n_670),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_866),
.B(n_669),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_916),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_952),
.B(n_929),
.Y(n_1076)
);

AND2x6_ASAP7_75t_L g1077 ( 
.A(n_895),
.B(n_740),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_924),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_916),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_828),
.Y(n_1080)
);

AND3x2_ASAP7_75t_SL g1081 ( 
.A(n_829),
.B(n_678),
.C(n_700),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_783),
.B(n_725),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_791),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_840),
.B(n_677),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_925),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_876),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_955),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_964),
.B(n_697),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_858),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_957),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_961),
.B(n_711),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_779),
.B1(n_299),
.B2(n_310),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_782),
.B(n_300),
.C(n_308),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_966),
.B(n_740),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_946),
.A2(n_386),
.B1(n_388),
.B2(n_440),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_810),
.B(n_740),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_909),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_872),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_810),
.B(n_744),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_883),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_952),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_826),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_799),
.Y(n_1103)
);

AOI22x1_ASAP7_75t_L g1104 ( 
.A1(n_968),
.A2(n_715),
.B1(n_718),
.B2(n_697),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_799),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_946),
.A2(n_456),
.B1(n_446),
.B2(n_440),
.Y(n_1106)
);

AND2x6_ASAP7_75t_L g1107 ( 
.A(n_895),
.B(n_896),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_912),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_833),
.A2(n_812),
.B1(n_937),
.B2(n_890),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_868),
.A2(n_301),
.B1(n_305),
.B2(n_718),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_848),
.A2(n_733),
.B(n_771),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_815),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_884),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_900),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_937),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_963),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_848),
.B(n_760),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_920),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_927),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_826),
.B(n_715),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_956),
.B(n_760),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_949),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_870),
.A2(n_944),
.B1(n_962),
.B2(n_897),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_972),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_908),
.A2(n_456),
.B(n_440),
.C(n_446),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_880),
.Y(n_1126)
);

OR2x4_ASAP7_75t_L g1127 ( 
.A(n_838),
.B(n_744),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_801),
.B(n_96),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1029),
.B(n_963),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1053),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1062),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1066),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1032),
.Y(n_1133)
);

CKINVDCx11_ASAP7_75t_R g1134 ( 
.A(n_1063),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1068),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_980),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1034),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_991),
.A2(n_969),
.B1(n_963),
.B2(n_870),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1034),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1008),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_1016),
.B(n_969),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1008),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1126),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_984),
.A2(n_918),
.B(n_859),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1072),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1085),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1126),
.Y(n_1147)
);

INVx8_ASAP7_75t_L g1148 ( 
.A(n_1033),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1031),
.B(n_803),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1076),
.A2(n_969),
.B1(n_901),
.B2(n_935),
.Y(n_1150)
);

BUFx2_ASAP7_75t_SL g1151 ( 
.A(n_1004),
.Y(n_1151)
);

BUFx8_ASAP7_75t_L g1152 ( 
.A(n_998),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1052),
.A2(n_973),
.B1(n_821),
.B2(n_853),
.C(n_971),
.Y(n_1153)
);

BUFx8_ASAP7_75t_SL g1154 ( 
.A(n_1018),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1102),
.B(n_1101),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1087),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1016),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1126),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1057),
.B(n_1042),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_997),
.A2(n_803),
.B1(n_806),
.B2(n_790),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_L g1162 ( 
.A(n_1093),
.B(n_815),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1090),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_997),
.A2(n_1125),
.B(n_986),
.C(n_984),
.Y(n_1164)
);

NAND3x1_ASAP7_75t_L g1165 ( 
.A(n_990),
.B(n_827),
.C(n_940),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1026),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1100),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1113),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1012),
.A2(n_790),
.B(n_896),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1076),
.A2(n_907),
.B1(n_936),
.B2(n_800),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1002),
.B(n_806),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1058),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_981),
.B(n_949),
.Y(n_1173)
);

AOI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1047),
.A2(n_971),
.B(n_970),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_1063),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1003),
.B(n_950),
.Y(n_1176)
);

NAND2x2_ASAP7_75t_L g1177 ( 
.A(n_1075),
.B(n_1079),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1082),
.A2(n_814),
.B(n_967),
.C(n_965),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1122),
.B(n_950),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_975),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_959),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1011),
.A2(n_922),
.B1(n_918),
.B2(n_859),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_992),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1078),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1012),
.A2(n_928),
.B(n_839),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_975),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1013),
.B(n_970),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1046),
.A2(n_839),
.B(n_851),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1116),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1025),
.A2(n_852),
.B1(n_933),
.B2(n_789),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1126),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_994),
.A2(n_951),
.B1(n_945),
.B2(n_939),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1082),
.A2(n_865),
.B(n_837),
.C(n_842),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1127),
.A2(n_879),
.B1(n_878),
.B2(n_864),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1098),
.Y(n_1195)
);

AOI222xp33_ASAP7_75t_L g1196 ( 
.A1(n_1064),
.A2(n_809),
.B1(n_804),
.B2(n_446),
.C1(n_456),
.C2(n_836),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_994),
.A2(n_856),
.B1(n_851),
.B2(n_860),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_987),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1059),
.B(n_860),
.Y(n_1199)
);

AND3x1_ASAP7_75t_SL g1200 ( 
.A(n_1044),
.B(n_0),
.C(n_2),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1075),
.B(n_891),
.Y(n_1201)
);

AND3x2_ASAP7_75t_L g1202 ( 
.A(n_1089),
.B(n_822),
.C(n_879),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1102),
.B(n_1060),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1046),
.A2(n_856),
.B(n_864),
.Y(n_1204)
);

OAI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1049),
.A2(n_932),
.B1(n_869),
.B2(n_878),
.C1(n_910),
.C2(n_902),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1056),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_993),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_999),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1097),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1022),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1033),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1056),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_975),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1033),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1060),
.B(n_869),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1024),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1026),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1037),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1020),
.A2(n_894),
.B1(n_881),
.B2(n_911),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_995),
.Y(n_1220)
);

BUFx4f_ASAP7_75t_L g1221 ( 
.A(n_1112),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_975),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1115),
.B(n_880),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1005),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1023),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1033),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_988),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_988),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1054),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1127),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_978),
.B(n_880),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_988),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1055),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1108),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1073),
.B(n_926),
.C(n_831),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1071),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1086),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1079),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1083),
.A2(n_899),
.B1(n_911),
.B2(n_910),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1114),
.A2(n_1080),
.B1(n_1123),
.B2(n_1043),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1007),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_978),
.Y(n_1242)
);

AOI221xp5_ASAP7_75t_L g1243 ( 
.A1(n_1043),
.A2(n_832),
.B1(n_867),
.B2(n_899),
.C(n_894),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_996),
.A2(n_760),
.B(n_744),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1017),
.A2(n_902),
.B1(n_881),
.B2(n_891),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1014),
.A2(n_880),
.B1(n_744),
.B2(n_760),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_1110),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_977),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1128),
.A2(n_913),
.B1(n_507),
.B2(n_505),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_982),
.B(n_805),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_988),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1040),
.A2(n_500),
.B1(n_443),
.B2(n_479),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_982),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1000),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1095),
.A2(n_500),
.B1(n_479),
.B2(n_485),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1028),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1000),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1065),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_996),
.A2(n_771),
.B(n_733),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1115),
.B(n_485),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1125),
.A2(n_408),
.B(n_423),
.C(n_3),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1070),
.B(n_1014),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1070),
.B(n_0),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_979),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1038),
.B(n_2),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_983),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1118),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_976),
.A2(n_391),
.B1(n_485),
.B2(n_479),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1000),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1103),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1103),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1065),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1000),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1001),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1120),
.B(n_83),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1001),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1040),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1105),
.Y(n_1278)
);

AOI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1048),
.A2(n_7),
.B(n_10),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1069),
.B(n_485),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1038),
.B(n_13),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1001),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1117),
.A2(n_479),
.B(n_423),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1149),
.A2(n_986),
.B(n_1111),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1135),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1247),
.A2(n_1073),
.B1(n_1007),
.B2(n_976),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1145),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1168),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1130),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1209),
.Y(n_1290)
);

AOI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1204),
.A2(n_1188),
.B(n_1169),
.Y(n_1291)
);

AOI221xp5_ASAP7_75t_L g1292 ( 
.A1(n_1279),
.A2(n_1048),
.B1(n_1095),
.B2(n_1084),
.C(n_1109),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_SL g1293 ( 
.A1(n_1261),
.A2(n_1036),
.B(n_1096),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1185),
.A2(n_1104),
.B(n_1015),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1265),
.A2(n_1030),
.B1(n_1084),
.B2(n_1094),
.C(n_1106),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1131),
.Y(n_1296)
);

INVx4_ASAP7_75t_SL g1297 ( 
.A(n_1194),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1133),
.B(n_1088),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1172),
.B(n_1119),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1132),
.Y(n_1300)
);

INVx4_ASAP7_75t_SL g1301 ( 
.A(n_1231),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1174),
.A2(n_1099),
.B(n_1067),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1146),
.Y(n_1303)
);

BUFx4f_ASAP7_75t_SL g1304 ( 
.A(n_1175),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1149),
.A2(n_985),
.B(n_1015),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1148),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1215),
.B(n_1069),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1235),
.A2(n_1092),
.B(n_1091),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1240),
.A2(n_1074),
.B1(n_1027),
.B2(n_1088),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1172),
.B(n_1124),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1156),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1176),
.B(n_1006),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1279),
.A2(n_1106),
.B1(n_1107),
.B2(n_1074),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1137),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1281),
.B(n_1120),
.C(n_1009),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1160),
.B(n_1006),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1174),
.A2(n_1111),
.B(n_1121),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1163),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1262),
.B(n_1009),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1193),
.A2(n_1178),
.B(n_1171),
.C(n_1179),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1283),
.A2(n_1121),
.B(n_989),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1161),
.A2(n_1192),
.B(n_1197),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1226),
.B(n_989),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1138),
.B(n_1019),
.C(n_1061),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1164),
.A2(n_1045),
.B(n_1050),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1209),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1244),
.A2(n_1245),
.B(n_1161),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1245),
.A2(n_1019),
.B(n_1061),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1219),
.A2(n_1105),
.B(n_1027),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1239),
.A2(n_1081),
.B(n_1041),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1259),
.A2(n_1081),
.B(n_1107),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1167),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1277),
.A2(n_1107),
.B1(n_1077),
.B2(n_1041),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1139),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1215),
.B(n_1041),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1235),
.A2(n_1107),
.B(n_1077),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1153),
.A2(n_1107),
.B(n_1077),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1243),
.A2(n_1077),
.B(n_408),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1219),
.A2(n_1077),
.A3(n_1041),
.B(n_1035),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1195),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1152),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1198),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1192),
.A2(n_1035),
.A3(n_1021),
.B(n_1010),
.Y(n_1343)
);

BUFx2_ASAP7_75t_SL g1344 ( 
.A(n_1166),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1144),
.A2(n_423),
.B(n_1021),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1208),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1263),
.B(n_1035),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1148),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1197),
.A2(n_423),
.B(n_1021),
.Y(n_1350)
);

AOI21xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1234),
.A2(n_14),
.B(n_19),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1181),
.A2(n_1035),
.B1(n_1021),
.B2(n_1010),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1241),
.B(n_1010),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1223),
.A2(n_1010),
.B(n_1001),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_SL g1355 ( 
.A1(n_1179),
.A2(n_19),
.B(n_23),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1173),
.A2(n_84),
.B(n_116),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1173),
.A2(n_23),
.B(n_25),
.C(n_27),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1241),
.B(n_25),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1148),
.B(n_1141),
.Y(n_1359)
);

INVx5_ASAP7_75t_L g1360 ( 
.A(n_1226),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1187),
.A2(n_391),
.B(n_36),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1210),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1216),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1199),
.B(n_32),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1218),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1205),
.A2(n_1252),
.B(n_1223),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1190),
.A2(n_1260),
.B(n_1129),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1162),
.A2(n_32),
.B1(n_36),
.B2(n_42),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1141),
.B(n_43),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1190),
.A2(n_43),
.A3(n_47),
.B(n_50),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1141),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1260),
.A2(n_114),
.B(n_53),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1152),
.Y(n_1373)
);

O2A1O1Ixp5_ASAP7_75t_SL g1374 ( 
.A1(n_1182),
.A2(n_51),
.B(n_55),
.C(n_61),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1189),
.B(n_71),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1154),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1203),
.B(n_73),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1150),
.A2(n_395),
.B1(n_82),
.B2(n_92),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1224),
.A2(n_1236),
.B1(n_1248),
.B2(n_1225),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1231),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1229),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1211),
.A2(n_80),
.B(n_93),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1249),
.A2(n_1182),
.B(n_1255),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1211),
.B(n_97),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1214),
.A2(n_107),
.B(n_119),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1237),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1214),
.B(n_122),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1275),
.A2(n_126),
.B(n_138),
.C(n_140),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1136),
.Y(n_1389)
);

OAI222xp33_ASAP7_75t_L g1390 ( 
.A1(n_1184),
.A2(n_1230),
.B1(n_1264),
.B2(n_1266),
.C1(n_1170),
.C2(n_1201),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1183),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1203),
.B(n_142),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1255),
.A2(n_144),
.B(n_152),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1242),
.B(n_157),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1275),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1250),
.A2(n_391),
.B(n_1233),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1207),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1258),
.A2(n_391),
.B1(n_1272),
.B2(n_1246),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1220),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1256),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1253),
.B(n_391),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1143),
.A2(n_1158),
.B(n_1191),
.C(n_1147),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1250),
.A2(n_1274),
.B(n_1269),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1270),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1143),
.A2(n_1191),
.B(n_1158),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1267),
.A2(n_1184),
.B1(n_1157),
.B2(n_1201),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1159),
.Y(n_1407)
);

CKINVDCx8_ASAP7_75t_R g1408 ( 
.A(n_1151),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1196),
.A2(n_1165),
.B(n_1268),
.Y(n_1409)
);

NOR2x1_ASAP7_75t_L g1410 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1147),
.A2(n_1278),
.B(n_1271),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1278),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1196),
.A2(n_1202),
.B(n_1177),
.Y(n_1413)
);

BUFx4_ASAP7_75t_SL g1414 ( 
.A(n_1206),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1180),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1180),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1280),
.A2(n_1257),
.B(n_1228),
.Y(n_1417)
);

AND2x4_ASAP7_75t_SL g1418 ( 
.A(n_1155),
.B(n_1201),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1155),
.B(n_1140),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1280),
.A2(n_1257),
.B(n_1228),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1280),
.A2(n_1222),
.B(n_1276),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1282),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1200),
.A2(n_1212),
.B1(n_1221),
.B2(n_1217),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1186),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1186),
.A2(n_1232),
.B(n_1276),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1186),
.A2(n_1232),
.A3(n_1276),
.B(n_1213),
.Y(n_1426)
);

AOI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1238),
.A2(n_1221),
.B1(n_1142),
.B2(n_1213),
.C(n_1227),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1282),
.B(n_1232),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_SL g1429 ( 
.A1(n_1213),
.A2(n_1222),
.B(n_1227),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_R g1430 ( 
.A(n_1134),
.B(n_1222),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1371),
.A2(n_1227),
.B1(n_1251),
.B2(n_1254),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1319),
.B(n_1251),
.Y(n_1432)
);

AOI222xp33_ASAP7_75t_L g1433 ( 
.A1(n_1368),
.A2(n_1251),
.B1(n_1254),
.B2(n_1273),
.C1(n_1282),
.C2(n_1371),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1291),
.A2(n_1284),
.B(n_1403),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1314),
.B(n_1334),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1347),
.B(n_1254),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1409),
.A2(n_1273),
.B1(n_1361),
.B2(n_1337),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1400),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1368),
.A2(n_1273),
.B1(n_1315),
.B2(n_1292),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1313),
.A2(n_1286),
.B1(n_1423),
.B2(n_1406),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1300),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1308),
.A2(n_1295),
.B(n_1320),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1359),
.B(n_1418),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1348),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1320),
.B(n_1367),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1294),
.A2(n_1305),
.B(n_1336),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_R g1447 ( 
.A1(n_1378),
.A2(n_1398),
.B(n_1309),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1300),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1303),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_R g1450 ( 
.A(n_1376),
.B(n_1389),
.Y(n_1450)
);

OAI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1298),
.A2(n_1322),
.B1(n_1359),
.B2(n_1312),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1313),
.A2(n_1423),
.B1(n_1406),
.B2(n_1388),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1408),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1311),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1355),
.A2(n_1369),
.B1(n_1338),
.B2(n_1383),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1359),
.B(n_1418),
.Y(n_1456)
);

INVx5_ASAP7_75t_L g1457 ( 
.A(n_1360),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1346),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1351),
.A2(n_1326),
.B1(n_1290),
.B2(n_1395),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1312),
.A2(n_1387),
.B1(n_1384),
.B2(n_1364),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_SL g1461 ( 
.A1(n_1388),
.A2(n_1390),
.B(n_1330),
.C(n_1427),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1294),
.A2(n_1321),
.B(n_1327),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1395),
.A2(n_1324),
.B1(n_1297),
.B2(n_1377),
.Y(n_1463)
);

BUFx4f_ASAP7_75t_SL g1464 ( 
.A(n_1341),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_SL g1465 ( 
.A1(n_1358),
.A2(n_1373),
.B(n_1394),
.C(n_1400),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1346),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1362),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1297),
.A2(n_1307),
.B1(n_1344),
.B2(n_1377),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1349),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1391),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1301),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1383),
.A2(n_1393),
.B1(n_1413),
.B2(n_1327),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1289),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1297),
.A2(n_1307),
.B1(n_1377),
.B2(n_1293),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1317),
.A2(n_1402),
.B(n_1302),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1349),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1314),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1393),
.A2(n_1366),
.B1(n_1357),
.B2(n_1341),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1407),
.B(n_1316),
.Y(n_1479)
);

NOR3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1376),
.B(n_1419),
.C(n_1299),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1428),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1307),
.A2(n_1356),
.B1(n_1335),
.B2(n_1367),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1367),
.B(n_1302),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1484)
);

BUFx10_ASAP7_75t_L g1485 ( 
.A(n_1419),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1335),
.A2(n_1380),
.B1(n_1304),
.B2(n_1392),
.Y(n_1486)
);

OR2x6_ASAP7_75t_SL g1487 ( 
.A(n_1375),
.B(n_1430),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1304),
.A2(n_1380),
.B1(n_1384),
.B2(n_1387),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1317),
.A2(n_1402),
.B(n_1302),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1379),
.A2(n_1365),
.B1(n_1363),
.B2(n_1332),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1334),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1357),
.A2(n_1342),
.B1(n_1340),
.B2(n_1318),
.C(n_1296),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1301),
.B(n_1335),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1301),
.B(n_1420),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1386),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1379),
.B(n_1386),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1391),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1366),
.A2(n_1285),
.B1(n_1287),
.B2(n_1288),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1397),
.B(n_1353),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1352),
.B(n_1366),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1321),
.A2(n_1328),
.B(n_1350),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1325),
.A2(n_1399),
.B1(n_1397),
.B2(n_1381),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1370),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1370),
.Y(n_1504)
);

AOI21xp33_ASAP7_75t_L g1505 ( 
.A1(n_1352),
.A2(n_1325),
.B(n_1333),
.Y(n_1505)
);

NAND2xp33_ASAP7_75t_SL g1506 ( 
.A(n_1306),
.B(n_1333),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1412),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1329),
.A2(n_1331),
.B(n_1345),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1348),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1370),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1360),
.B(n_1329),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1424),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1360),
.B(n_1404),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_SL g1514 ( 
.A1(n_1323),
.A2(n_1415),
.B1(n_1422),
.B2(n_1416),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1404),
.A2(n_1410),
.B1(n_1401),
.B2(n_1306),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1348),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1424),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1360),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1425),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1414),
.B(n_1429),
.Y(n_1520)
);

AOI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1345),
.A2(n_1328),
.B(n_1372),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1426),
.Y(n_1522)
);

AOI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1411),
.A2(n_1354),
.B(n_1385),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1411),
.B(n_1417),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1370),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1396),
.A2(n_1382),
.B1(n_1323),
.B2(n_1417),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1343),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1343),
.B(n_1339),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1374),
.A2(n_1396),
.B1(n_1425),
.B2(n_1414),
.C(n_1343),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1405),
.A2(n_1421),
.B1(n_1343),
.B2(n_1339),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1426),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1339),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1339),
.A2(n_1247),
.B1(n_664),
.B2(n_437),
.Y(n_1533)
);

NAND2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1426),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1300),
.Y(n_1536)
);

BUFx4f_ASAP7_75t_L g1537 ( 
.A(n_1377),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1319),
.B(n_1347),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1409),
.A2(n_563),
.B1(n_1281),
.B2(n_1265),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1300),
.Y(n_1540)
);

NOR3xp33_ASAP7_75t_SL g1541 ( 
.A(n_1315),
.B(n_1114),
.C(n_1083),
.Y(n_1541)
);

NAND4xp25_ASAP7_75t_L g1542 ( 
.A(n_1371),
.B(n_544),
.C(n_400),
.D(n_782),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1300),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1368),
.A2(n_1247),
.B1(n_664),
.B2(n_705),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1300),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1300),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1319),
.B(n_1347),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1314),
.B(n_1334),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1359),
.B(n_1418),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1368),
.A2(n_1247),
.B1(n_664),
.B2(n_705),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1473),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1527),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_R g1553 ( 
.A(n_1541),
.B(n_1480),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1481),
.Y(n_1554)
);

BUFx2_ASAP7_75t_SL g1555 ( 
.A(n_1453),
.Y(n_1555)
);

AO31x2_ASAP7_75t_L g1556 ( 
.A1(n_1475),
.A2(n_1489),
.A3(n_1508),
.B(n_1525),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1539),
.A2(n_1550),
.B(n_1544),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_R g1558 ( 
.A(n_1450),
.B(n_1537),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1539),
.A2(n_1542),
.B1(n_1440),
.B2(n_1452),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1464),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1538),
.B(n_1547),
.Y(n_1561)
);

AND2x4_ASAP7_75t_SL g1562 ( 
.A(n_1485),
.B(n_1494),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1484),
.B(n_1436),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1448),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1477),
.Y(n_1565)
);

AND2x2_ASAP7_75t_SL g1566 ( 
.A(n_1537),
.B(n_1492),
.Y(n_1566)
);

AO31x2_ASAP7_75t_L g1567 ( 
.A1(n_1475),
.A2(n_1489),
.A3(n_1508),
.B(n_1504),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1432),
.B(n_1499),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1434),
.A2(n_1462),
.B(n_1521),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_R g1570 ( 
.A(n_1541),
.B(n_1494),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1442),
.A2(n_1452),
.B(n_1437),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1491),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1435),
.B(n_1548),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1501),
.A2(n_1523),
.B(n_1511),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1438),
.B(n_1533),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1447),
.A2(n_1440),
.B1(n_1474),
.B2(n_1437),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1441),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_SL g1578 ( 
.A(n_1433),
.B(n_1442),
.C(n_1492),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1511),
.B(n_1524),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1479),
.B(n_1454),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1458),
.Y(n_1581)
);

INVx4_ASAP7_75t_SL g1582 ( 
.A(n_1471),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1463),
.A2(n_1459),
.B1(n_1468),
.B2(n_1488),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1449),
.B(n_1543),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1443),
.B(n_1456),
.Y(n_1585)
);

INVx4_ASAP7_75t_SL g1586 ( 
.A(n_1471),
.Y(n_1586)
);

INVxp33_ASAP7_75t_SL g1587 ( 
.A(n_1520),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1466),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_R g1589 ( 
.A(n_1506),
.B(n_1471),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1439),
.A2(n_1431),
.B(n_1455),
.C(n_1478),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1503),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1467),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1546),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1431),
.A2(n_1455),
.B1(n_1447),
.B2(n_1478),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1529),
.B(n_1513),
.C(n_1490),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1485),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1536),
.B(n_1540),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_R g1599 ( 
.A(n_1469),
.B(n_1476),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_SL g1600 ( 
.A(n_1493),
.B(n_1443),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1510),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1532),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1456),
.B(n_1549),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1495),
.B(n_1490),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1507),
.Y(n_1605)
);

BUFx10_ASAP7_75t_L g1606 ( 
.A(n_1516),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1507),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1512),
.B(n_1517),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1470),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1524),
.B(n_1445),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1496),
.Y(n_1611)
);

AND2x2_ASAP7_75t_SL g1612 ( 
.A(n_1445),
.B(n_1500),
.Y(n_1612)
);

NAND2xp33_ASAP7_75t_R g1613 ( 
.A(n_1549),
.B(n_1476),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1497),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1487),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1534),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1483),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1460),
.A2(n_1486),
.B1(n_1498),
.B2(n_1451),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1534),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1535),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1493),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1517),
.B(n_1482),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1522),
.B(n_1531),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1515),
.A2(n_1472),
.B1(n_1502),
.B2(n_1526),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1617),
.B(n_1483),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1528),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1617),
.B(n_1528),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1556),
.B(n_1446),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1588),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1611),
.B(n_1578),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1610),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1612),
.B(n_1446),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1579),
.B(n_1530),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1566),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1591),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1612),
.B(n_1472),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1610),
.B(n_1519),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1559),
.A2(n_1505),
.B1(n_1529),
.B2(n_1514),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1519),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1579),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1556),
.B(n_1505),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1556),
.B(n_1517),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1579),
.B(n_1457),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1601),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1567),
.B(n_1516),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1567),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1577),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1623),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1581),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1567),
.B(n_1516),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1592),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1552),
.B(n_1457),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1559),
.A2(n_1461),
.B1(n_1465),
.B2(n_1469),
.C(n_1518),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1573),
.B(n_1444),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1565),
.B(n_1444),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1564),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1623),
.Y(n_1657)
);

INVx3_ASAP7_75t_SL g1658 ( 
.A(n_1566),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1616),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1574),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1552),
.B(n_1457),
.Y(n_1661)
);

AND2x4_ASAP7_75t_SL g1662 ( 
.A(n_1622),
.B(n_1518),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1636),
.B(n_1631),
.Y(n_1663)
);

OAI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1658),
.A2(n_1557),
.B1(n_1571),
.B2(n_1590),
.C(n_1576),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1630),
.A2(n_1590),
.B1(n_1575),
.B2(n_1624),
.C(n_1594),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1630),
.A2(n_1594),
.B(n_1596),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1634),
.B(n_1558),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1636),
.B(n_1619),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1654),
.B(n_1572),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1634),
.A2(n_1658),
.B1(n_1636),
.B2(n_1638),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1654),
.B(n_1580),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1646),
.A2(n_1569),
.B(n_1596),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1568),
.Y(n_1673)
);

NAND4xp25_ASAP7_75t_L g1674 ( 
.A(n_1638),
.B(n_1618),
.C(n_1583),
.D(n_1553),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1626),
.B(n_1554),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1626),
.B(n_1563),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1602),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_L g1678 ( 
.A(n_1653),
.B(n_1618),
.C(n_1553),
.D(n_1604),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1653),
.A2(n_1607),
.B1(n_1605),
.B2(n_1561),
.C(n_1551),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1626),
.B(n_1598),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1626),
.B(n_1614),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1631),
.B(n_1602),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1658),
.A2(n_1587),
.B1(n_1615),
.B2(n_1597),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1631),
.B(n_1621),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1625),
.B(n_1562),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1625),
.B(n_1608),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1646),
.A2(n_1620),
.B(n_1593),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1625),
.B(n_1609),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1625),
.B(n_1656),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.B(n_1562),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1632),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1632),
.A2(n_1584),
.B1(n_1570),
.B2(n_1589),
.C(n_1558),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1633),
.A2(n_1603),
.B(n_1585),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1656),
.B(n_1603),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1656),
.B(n_1585),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1589),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1658),
.A2(n_1555),
.B1(n_1457),
.B2(n_1509),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1599),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1634),
.B(n_1570),
.C(n_1613),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1633),
.A2(n_1600),
.B(n_1582),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1634),
.B(n_1613),
.C(n_1509),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1629),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1658),
.A2(n_1560),
.B1(n_1582),
.B2(n_1586),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1647),
.B(n_1599),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1634),
.A2(n_1582),
.B1(n_1586),
.B2(n_1606),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1684),
.B(n_1640),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1663),
.B(n_1684),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1663),
.B(n_1662),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1677),
.B(n_1662),
.Y(n_1710)
);

NAND2x1_ASAP7_75t_L g1711 ( 
.A(n_1702),
.B(n_1634),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1686),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1677),
.B(n_1662),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1668),
.B(n_1662),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1703),
.Y(n_1716)
);

NOR2xp67_ASAP7_75t_L g1717 ( 
.A(n_1700),
.B(n_1640),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1688),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1692),
.B(n_1627),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1690),
.B(n_1627),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1703),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1669),
.B(n_1647),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1682),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1681),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1688),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1675),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1668),
.B(n_1657),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1671),
.B(n_1649),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1676),
.B(n_1649),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1680),
.B(n_1627),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1689),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1673),
.B(n_1649),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1682),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1691),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1687),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1695),
.B(n_1627),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1696),
.Y(n_1739)
);

NAND2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1683),
.B(n_1640),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1685),
.B(n_1657),
.Y(n_1741)
);

AND2x2_ASAP7_75t_SL g1742 ( 
.A(n_1670),
.B(n_1643),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1702),
.B(n_1640),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1712),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1717),
.B(n_1685),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1712),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_1691),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1713),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1708),
.B(n_1694),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1733),
.B(n_1697),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1724),
.B(n_1665),
.Y(n_1752)
);

AND2x4_ASAP7_75t_SL g1753 ( 
.A(n_1709),
.B(n_1643),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1709),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1743),
.B(n_1657),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1707),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1743),
.B(n_1657),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1666),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1716),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1743),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1733),
.B(n_1705),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1723),
.B(n_1648),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1716),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1710),
.B(n_1714),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1726),
.B(n_1666),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1710),
.B(n_1648),
.Y(n_1766)
);

NAND2x1p5_ASAP7_75t_L g1767 ( 
.A(n_1711),
.B(n_1667),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1718),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1721),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1730),
.B(n_1699),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1718),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1737),
.B(n_1731),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1714),
.B(n_1648),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1651),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1721),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1715),
.B(n_1701),
.Y(n_1776)
);

NAND2x1_ASAP7_75t_L g1777 ( 
.A(n_1707),
.B(n_1700),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1707),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1715),
.B(n_1639),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1730),
.B(n_1672),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1742),
.B(n_1639),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1722),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1727),
.Y(n_1783)
);

NAND2xp33_ASAP7_75t_R g1784 ( 
.A(n_1741),
.B(n_1643),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1742),
.B(n_1639),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1744),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1752),
.A2(n_1664),
.B1(n_1674),
.B2(n_1678),
.C(n_1679),
.Y(n_1787)
);

NAND2x1p5_ASAP7_75t_L g1788 ( 
.A(n_1777),
.B(n_1711),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1777),
.B(n_1704),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1756),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1744),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1764),
.B(n_1736),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1756),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1764),
.B(n_1741),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1746),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1747),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1752),
.B(n_1731),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1767),
.A2(n_1706),
.B1(n_1698),
.B2(n_1739),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1758),
.B(n_1739),
.Y(n_1799)
);

NAND4xp75_ASAP7_75t_SL g1800 ( 
.A(n_1781),
.B(n_1672),
.C(n_1637),
.D(n_1639),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1746),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1765),
.B(n_1740),
.Y(n_1802)
);

OAI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1767),
.A2(n_1738),
.B1(n_1719),
.B2(n_1732),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1765),
.B(n_1728),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1751),
.B(n_1729),
.Y(n_1805)
);

INVxp33_ASAP7_75t_L g1806 ( 
.A(n_1776),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1767),
.A2(n_1693),
.B1(n_1719),
.B2(n_1738),
.C(n_1720),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1748),
.Y(n_1808)
);

OAI322xp33_ASAP7_75t_L g1809 ( 
.A1(n_1758),
.A2(n_1735),
.A3(n_1734),
.B1(n_1720),
.B2(n_1628),
.C1(n_1725),
.C2(n_1641),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1748),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1760),
.B(n_1641),
.C(n_1734),
.D(n_1735),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1750),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1750),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1747),
.B(n_1727),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1760),
.A2(n_1783),
.B1(n_1754),
.B2(n_1778),
.Y(n_1815)
);

OAI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1784),
.A2(n_1672),
.B1(n_1628),
.B2(n_1642),
.Y(n_1816)
);

OA222x2_ASAP7_75t_L g1817 ( 
.A1(n_1780),
.A2(n_1725),
.B1(n_1628),
.B2(n_1642),
.C1(n_1655),
.C2(n_1646),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1751),
.B(n_1655),
.Y(n_1818)
);

O2A1O1Ixp5_ASAP7_75t_R g1819 ( 
.A1(n_1772),
.A2(n_1672),
.B(n_1659),
.C(n_1655),
.Y(n_1819)
);

OA222x2_ASAP7_75t_L g1820 ( 
.A1(n_1780),
.A2(n_1628),
.B1(n_1642),
.B2(n_1646),
.C1(n_1651),
.C2(n_1660),
.Y(n_1820)
);

OR2x6_ASAP7_75t_L g1821 ( 
.A(n_1789),
.B(n_1778),
.Y(n_1821)
);

NAND2xp67_ASAP7_75t_SL g1822 ( 
.A(n_1787),
.B(n_1776),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1806),
.B(n_1749),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1790),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1793),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1789),
.Y(n_1827)
);

AOI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1789),
.A2(n_1745),
.B(n_1755),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1791),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1794),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1804),
.B(n_1749),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1802),
.B(n_1783),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1795),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1815),
.Y(n_1834)
);

OAI32xp33_ASAP7_75t_L g1835 ( 
.A1(n_1788),
.A2(n_1761),
.A3(n_1781),
.B1(n_1785),
.B2(n_1772),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1797),
.B(n_1785),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1792),
.B(n_1754),
.Y(n_1837)
);

NAND3xp33_ASAP7_75t_L g1838 ( 
.A(n_1815),
.B(n_1782),
.C(n_1761),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1788),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1797),
.B(n_1770),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1799),
.B(n_1782),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1799),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1796),
.B(n_1762),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1801),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1814),
.B(n_1745),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1827),
.B(n_1803),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1822),
.B(n_1807),
.C(n_1819),
.Y(n_1847)
);

OAI222xp33_ASAP7_75t_L g1848 ( 
.A1(n_1821),
.A2(n_1798),
.B1(n_1816),
.B2(n_1805),
.C1(n_1818),
.C2(n_1770),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1821),
.A2(n_1823),
.B(n_1835),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1825),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1821),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1834),
.B(n_1762),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1837),
.B(n_1755),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1834),
.A2(n_1811),
.B(n_1808),
.C(n_1813),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1824),
.B(n_1812),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1826),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1831),
.A2(n_1753),
.B1(n_1757),
.B2(n_1779),
.Y(n_1857)
);

OAI32xp33_ASAP7_75t_L g1858 ( 
.A1(n_1836),
.A2(n_1811),
.A3(n_1820),
.B1(n_1817),
.B2(n_1810),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1824),
.Y(n_1859)
);

NOR2x1_ASAP7_75t_L g1860 ( 
.A(n_1839),
.B(n_1800),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1829),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1837),
.A2(n_1757),
.B1(n_1753),
.B2(n_1766),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1845),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1839),
.B(n_1809),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1859),
.Y(n_1865)
);

XOR2x2_ASAP7_75t_L g1866 ( 
.A(n_1847),
.B(n_1832),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1855),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1847),
.A2(n_1840),
.B1(n_1836),
.B2(n_1838),
.C(n_1828),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1856),
.B(n_1842),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1853),
.B(n_1830),
.Y(n_1870)
);

AOI32xp33_ASAP7_75t_L g1871 ( 
.A1(n_1864),
.A2(n_1840),
.A3(n_1830),
.B1(n_1844),
.B2(n_1833),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1851),
.B(n_1843),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1848),
.A2(n_1841),
.B(n_1759),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1850),
.Y(n_1874)
);

AOI222xp33_ASAP7_75t_L g1875 ( 
.A1(n_1858),
.A2(n_1763),
.B1(n_1775),
.B2(n_1759),
.C1(n_1769),
.C2(n_1771),
.Y(n_1875)
);

OAI32xp33_ASAP7_75t_L g1876 ( 
.A1(n_1868),
.A2(n_1849),
.A3(n_1846),
.B1(n_1852),
.B2(n_1863),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1871),
.A2(n_1854),
.B1(n_1861),
.B2(n_1857),
.C(n_1862),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1865),
.A2(n_1860),
.B1(n_1854),
.B2(n_1753),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1870),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1872),
.B(n_1774),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1873),
.A2(n_1763),
.B1(n_1775),
.B2(n_1769),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1867),
.A2(n_1768),
.B1(n_1771),
.B2(n_1774),
.C(n_1641),
.Y(n_1882)
);

AOI211xp5_ASAP7_75t_L g1883 ( 
.A1(n_1869),
.A2(n_1771),
.B(n_1768),
.C(n_1773),
.Y(n_1883)
);

OAI211xp5_ASAP7_75t_L g1884 ( 
.A1(n_1875),
.A2(n_1768),
.B(n_1773),
.C(n_1766),
.Y(n_1884)
);

OA211x2_ASAP7_75t_L g1885 ( 
.A1(n_1866),
.A2(n_1586),
.B(n_1779),
.C(n_1606),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1881),
.A2(n_1875),
.B(n_1874),
.Y(n_1886)
);

OA22x2_ASAP7_75t_L g1887 ( 
.A1(n_1878),
.A2(n_1659),
.B1(n_1643),
.B2(n_1633),
.Y(n_1887)
);

INVx4_ASAP7_75t_SL g1888 ( 
.A(n_1879),
.Y(n_1888)
);

NOR2x1_ASAP7_75t_L g1889 ( 
.A(n_1880),
.B(n_1884),
.Y(n_1889)
);

NOR2x1_ASAP7_75t_L g1890 ( 
.A(n_1885),
.B(n_1660),
.Y(n_1890)
);

AOI321xp33_ASAP7_75t_L g1891 ( 
.A1(n_1889),
.A2(n_1876),
.A3(n_1877),
.B1(n_1883),
.B2(n_1882),
.C(n_1633),
.Y(n_1891)
);

NOR4xp75_ASAP7_75t_L g1892 ( 
.A(n_1888),
.B(n_1659),
.C(n_1637),
.D(n_1645),
.Y(n_1892)
);

O2A1O1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1886),
.A2(n_1890),
.B(n_1887),
.C(n_1641),
.Y(n_1893)
);

AND4x1_ASAP7_75t_L g1894 ( 
.A(n_1889),
.B(n_1637),
.C(n_1645),
.D(n_1650),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1888),
.B(n_1660),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1886),
.A2(n_1637),
.B(n_1660),
.C(n_1645),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1895),
.Y(n_1897)
);

OAI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1891),
.A2(n_1894),
.B1(n_1892),
.B2(n_1896),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1893),
.A2(n_1659),
.B1(n_1643),
.B2(n_1642),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1895),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1895),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1901),
.Y(n_1902)
);

NOR2x1_ASAP7_75t_L g1903 ( 
.A(n_1897),
.B(n_1900),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1898),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1903),
.Y(n_1905)
);

NAND2xp33_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1904),
.Y(n_1906)
);

XOR2xp5_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1902),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1906),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1907),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1908),
.Y(n_1910)
);

AND3x4_ASAP7_75t_L g1911 ( 
.A(n_1910),
.B(n_1909),
.C(n_1899),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1910),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_SL g1913 ( 
.A(n_1912),
.B(n_1661),
.C(n_1652),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1913),
.A2(n_1911),
.B1(n_1644),
.B2(n_1635),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1914),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1643),
.B(n_1644),
.Y(n_1916)
);

AOI22x1_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1651),
.B1(n_1633),
.B2(n_1635),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1650),
.B1(n_1645),
.B2(n_1633),
.Y(n_1918)
);

AOI211xp5_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1661),
.B(n_1652),
.C(n_1650),
.Y(n_1919)
);


endmodule