module fake_jpeg_32156_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_5),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_22),
.B(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_10),
.B1(n_21),
.B2(n_19),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_15),
.B(n_12),
.Y(n_31)
);

A2O1A1O1Ixp25_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_17),
.B(n_20),
.C(n_14),
.D(n_12),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_26),
.Y(n_37)
);

OAI22x1_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_28),
.B1(n_25),
.B2(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_27),
.C(n_26),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_41),
.B1(n_38),
.B2(n_42),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_38),
.Y(n_45)
);


endmodule