module fake_jpeg_20500_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_24),
.B1(n_32),
.B2(n_28),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_20),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_56),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_24),
.B1(n_31),
.B2(n_37),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_60),
.A2(n_70),
.B1(n_34),
.B2(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_27),
.Y(n_103)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_20),
.B1(n_31),
.B2(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_26),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_23),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_76),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_18),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_78),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_20),
.B1(n_30),
.B2(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_79),
.A2(n_87),
.B1(n_97),
.B2(n_36),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_42),
.Y(n_80)
);

MAJx3_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_16),
.C(n_1),
.Y(n_144)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_84),
.B(n_89),
.Y(n_146)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_30),
.B1(n_17),
.B2(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_30),
.B1(n_17),
.B2(n_59),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_39),
.C(n_27),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_102),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_17),
.A3(n_19),
.B1(n_35),
.B2(n_22),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_19),
.B(n_22),
.C(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_33),
.C(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_112),
.Y(n_139)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_54),
.B(n_35),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_19),
.B1(n_35),
.B2(n_22),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_116),
.A2(n_92),
.B1(n_88),
.B2(n_113),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_83),
.B1(n_113),
.B2(n_82),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_19),
.B1(n_36),
.B2(n_16),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_141),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_36),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_149),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_0),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_75),
.B(n_16),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_117),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_107),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_173),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_81),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_123),
.B1(n_119),
.B2(n_134),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_98),
.B1(n_105),
.B2(n_73),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_137),
.B1(n_128),
.B2(n_144),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_171),
.B1(n_126),
.B2(n_145),
.Y(n_197)
);

OAI22x1_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_80),
.B1(n_106),
.B2(n_74),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_180),
.B1(n_145),
.B2(n_126),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_167),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_80),
.C(n_111),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_130),
.C(n_114),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_3),
.C(n_4),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_85),
.B1(n_101),
.B2(n_94),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_116),
.B(n_9),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_12),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_182),
.B(n_153),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_9),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_3),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_3),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_136),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_188),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_130),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_177),
.B(n_152),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_136),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_115),
.C(n_135),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_204),
.C(n_210),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_211),
.B1(n_167),
.B2(n_153),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_174),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_170),
.C(n_6),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_115),
.C(n_149),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_122),
.C(n_120),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_120),
.B1(n_122),
.B2(n_138),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_227),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_151),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_236),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_226),
.A2(n_234),
.B1(n_193),
.B2(n_214),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_180),
.B1(n_172),
.B2(n_170),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_185),
.C(n_190),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_237),
.C(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_157),
.B1(n_176),
.B2(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_198),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_169),
.C(n_168),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_4),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_240),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_187),
.B1(n_194),
.B2(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_225),
.B1(n_220),
.B2(n_230),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_187),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_252),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_211),
.B(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_255),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_259),
.B1(n_217),
.B2(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_214),
.C(n_207),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_261),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_226),
.A2(n_205),
.B1(n_196),
.B2(n_183),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_202),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_274),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_221),
.B1(n_217),
.B2(n_230),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_265),
.A2(n_266),
.B1(n_281),
.B2(n_245),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_238),
.B1(n_219),
.B2(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_205),
.B1(n_241),
.B2(n_236),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_273),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_235),
.B1(n_233),
.B2(n_231),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_249),
.A2(n_237),
.B1(n_215),
.B2(n_239),
.Y(n_281)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_250),
.B(n_262),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_246),
.C(n_258),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_247),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_242),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_261),
.C(n_250),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_254),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_245),
.C(n_7),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_269),
.B(n_270),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_283),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_274),
.B1(n_273),
.B2(n_265),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_279),
.B1(n_276),
.B2(n_275),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_303),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_272),
.B(n_7),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_285),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_313),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_282),
.B(n_286),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_287),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_299),
.B(n_300),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_309),
.B(n_311),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_301),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_315),
.C(n_314),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_321),
.C(n_318),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_316),
.B1(n_304),
.B2(n_298),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_282),
.B(n_7),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_10),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_10),
.B(n_11),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_12),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_12),
.B(n_14),
.Y(n_330)
);


endmodule