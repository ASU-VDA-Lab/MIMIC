module real_jpeg_33470_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_150;
wire n_74;
wire n_41;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_240;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_295;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_0),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_0),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_1),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_1),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_2),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_2),
.B(n_27),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_2),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_3),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

AND2x4_ASAP7_75t_SL g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

NAND2x1_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_111),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_7),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_8),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_8),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_8),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_9),
.B(n_111),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_10),
.B(n_98),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_R g123 ( 
.A(n_10),
.B(n_124),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_10),
.A2(n_15),
.B1(n_124),
.B2(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_10),
.B(n_167),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g212 ( 
.A(n_10),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_10),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_10),
.B(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_13),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_13),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_13),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_13),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_14),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_15),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_15),
.B(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_179),
.B1(n_296),
.B2(n_297),
.Y(n_18)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_19),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_R g19 ( 
.A(n_20),
.B(n_176),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI221xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_104),
.B1(n_152),
.B2(n_153),
.C(n_154),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_23),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_23),
.B(n_104),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_65),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.C(n_51),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_25),
.B(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_26),
.B(n_35),
.C(n_39),
.Y(n_142)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_38),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_41),
.B(n_52),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_172)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_50),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_50),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_50),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.C(n_61),
.Y(n_52)
);

XNOR2x1_ASAP7_75t_SL g160 ( 
.A(n_53),
.B(n_57),
.Y(n_160)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_61),
.B(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_91),
.B2(n_92),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2x2_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_72),
.Y(n_276)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_86),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_89),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_90),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_138),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_122),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_122),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_115),
.C(n_118),
.Y(n_108)
);

XNOR2x2_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_188),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_112),
.Y(n_190)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_119),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_129),
.B(n_134),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_134),
.Y(n_140)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_173),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_182),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_172),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_172),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_168),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

AO21x2_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_200),
.B(n_295),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_181),
.B(n_183),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_185),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_187),
.B(n_189),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.C(n_196),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_196),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

AO22x1_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_199),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_289),
.B(n_294),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_240),
.B(n_288),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_232),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_203),
.B(n_232),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_218),
.B(n_231),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_205),
.B(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_215),
.C(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_234),
.B(n_238),
.C(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_253),
.B(n_287),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_251),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_251),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.C(n_249),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_244),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_244),
.B(n_268),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_249),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_270),
.B(n_284),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_267),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_261),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_278),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_277),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_292),
.Y(n_294)
);


endmodule