module fake_jpeg_15296_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_33),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_21),
.CI(n_26),
.CON(n_41),
.SN(n_41)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_18),
.B1(n_24),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_18),
.B1(n_27),
.B2(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_21),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_63),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_62),
.B1(n_48),
.B2(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_39),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_16),
.C(n_47),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_13),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_30),
.B1(n_29),
.B2(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_33),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_29),
.C(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_73),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_45),
.B1(n_48),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_72),
.B1(n_58),
.B2(n_59),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_14),
.C(n_39),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_23),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_46),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_22),
.B(n_19),
.C(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_89),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_74),
.B1(n_79),
.B2(n_73),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_55),
.C(n_33),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_88),
.Y(n_100)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_53),
.C(n_61),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_53),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_71),
.B1(n_77),
.B2(n_75),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_95),
.C(n_3),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_105),
.B1(n_103),
.B2(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_81),
.Y(n_101)
);

OR2x6_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_74),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_103),
.B(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_74),
.B1(n_91),
.B2(n_94),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_70),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_106),
.B(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_107),
.A2(n_8),
.B1(n_11),
.B2(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_98),
.C(n_102),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_104),
.Y(n_120)
);

BUFx12f_ASAP7_75t_SL g111 ( 
.A(n_102),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_102),
.B(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_88),
.B1(n_82),
.B2(n_17),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_9),
.C(n_7),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_3),
.B(n_4),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_100),
.C(n_23),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_125),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_128),
.B1(n_122),
.B2(n_17),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_4),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

OR2x6_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_5),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_124),
.B(n_17),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_131),
.B(n_23),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_134),
.C(n_23),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_137),
.Y(n_139)
);


endmodule