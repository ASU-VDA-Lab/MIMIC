module fake_netlist_1_8926_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_7), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
AOI21x1_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_9), .B(n_1), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_14), .B(n_0), .C(n_2), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_17), .B(n_2), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_14), .B(n_8), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_13), .B(n_8), .Y(n_22) );
NOR2xp33_ASAP7_75t_R g23 ( .A(n_18), .B(n_16), .Y(n_23) );
NAND2xp33_ASAP7_75t_R g24 ( .A(n_19), .B(n_15), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_21), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_22), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_11), .B1(n_17), .B2(n_23), .Y(n_29) );
AOI211xp5_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_28), .B(n_26), .C(n_6), .Y(n_30) );
A2O1A1Ixp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_17), .B(n_4), .C(n_5), .Y(n_31) );
AND2x4_ASAP7_75t_L g32 ( .A(n_31), .B(n_17), .Y(n_32) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
BUFx2_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_4), .B1(n_32), .B2(n_35), .Y(n_36) );
endmodule