module fake_jpeg_27915_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_59),
.Y(n_66)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_45),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_56),
.C(n_54),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_49),
.B1(n_56),
.B2(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_73),
.B1(n_74),
.B2(n_1),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_57),
.B1(n_46),
.B2(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_51),
.B1(n_47),
.B2(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_55),
.B1(n_53),
.B2(n_42),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_92),
.B1(n_96),
.B2(n_2),
.Y(n_104)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_88),
.B1(n_85),
.B2(n_81),
.Y(n_102)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_1),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_87),
.C(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_104),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_16),
.B(n_31),
.C(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_111),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_91),
.B(n_86),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_112),
.B(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_7),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_102),
.B1(n_105),
.B2(n_101),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_119),
.B1(n_8),
.B2(n_10),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_103),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_11),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.C(n_122),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_118),
.C(n_117),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_123),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_116),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_21),
.C(n_22),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_23),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_41),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_27),
.Y(n_134)
);


endmodule