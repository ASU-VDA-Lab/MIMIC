module fake_aes_10361_n_616 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_616);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_616;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_25), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_70), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_50), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_47), .Y(n_75) );
HB1xp67_ASAP7_75t_L g76 ( .A(n_3), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_71), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_26), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_57), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_59), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_66), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_19), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_24), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_11), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_28), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_40), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_36), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_69), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_10), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_4), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_33), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_38), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_9), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_68), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_39), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_29), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_49), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_18), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_62), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_42), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_61), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_48), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_13), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_54), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_13), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_16), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_87), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_102), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
NOR2xp33_ASAP7_75t_R g119 ( .A(n_102), .B(n_27), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_87), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_76), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_95), .B(n_1), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_108), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_86), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_112), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_73), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_97), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_99), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_73), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_74), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_74), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_113), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_75), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_106), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_85), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_115), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_75), .Y(n_147) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_78), .A2(n_30), .B(n_65), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_98), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_72), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_88), .B(n_2), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_78), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_79), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_79), .Y(n_154) );
AO22x2_ASAP7_75t_L g155 ( .A1(n_151), .A2(n_100), .B1(n_111), .B2(n_110), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_145), .B(n_107), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_150), .B(n_77), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_135), .B(n_94), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_117), .B(n_93), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_135), .B(n_107), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_143), .B(n_114), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_133), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_138), .B(n_81), .Y(n_168) );
NAND3xp33_ASAP7_75t_L g169 ( .A(n_121), .B(n_114), .C(n_88), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_121), .B(n_109), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_151), .B(n_111), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_151), .B(n_109), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_138), .B(n_90), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_139), .B(n_92), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_139), .B(n_104), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_116), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_142), .B(n_110), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_142), .B(n_105), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_152), .B(n_105), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_116), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_116), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_136), .B(n_96), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_152), .B(n_96), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_116), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_116), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_122), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_118), .Y(n_191) );
OAI22x1_ASAP7_75t_L g192 ( .A1(n_144), .A2(n_104), .B1(n_103), .B2(n_100), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_154), .B(n_103), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_118), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_154), .B(n_93), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_122), .B(n_91), .Y(n_198) );
BUFx4_ASAP7_75t_L g199 ( .A(n_125), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_129), .A2(n_132), .B1(n_149), .B2(n_146), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_118), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_190), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_190), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_187), .Y(n_206) );
OR2x6_ASAP7_75t_L g207 ( .A(n_200), .B(n_153), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_187), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_166), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_187), .Y(n_212) );
NOR3xp33_ASAP7_75t_SL g213 ( .A(n_200), .B(n_141), .C(n_137), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_172), .Y(n_214) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_174), .B(n_148), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_172), .A2(n_153), .B1(n_124), .B2(n_123), .Y(n_216) );
NOR2xp33_ASAP7_75t_R g217 ( .A(n_164), .B(n_123), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_190), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_197), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_168), .B(n_153), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_169), .B(n_134), .Y(n_221) );
AND3x2_ASAP7_75t_SL g222 ( .A(n_199), .B(n_119), .C(n_127), .Y(n_222) );
CKINVDCx8_ASAP7_75t_R g223 ( .A(n_174), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_179), .Y(n_224) );
NAND2xp33_ASAP7_75t_L g225 ( .A(n_197), .B(n_147), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_171), .B(n_134), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_156), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_197), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_156), .B(n_134), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g231 ( .A(n_163), .B(n_101), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_171), .B(n_134), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_164), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_163), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_158), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_176), .B(n_124), .Y(n_236) );
BUFx12f_ASAP7_75t_L g237 ( .A(n_174), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_174), .B(n_131), .Y(n_238) );
OR2x6_ASAP7_75t_L g239 ( .A(n_199), .B(n_83), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_159), .B(n_131), .Y(n_241) );
INVx6_ASAP7_75t_L g242 ( .A(n_177), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_155), .A2(n_120), .B1(n_127), .B2(n_126), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_161), .B(n_128), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_177), .B(n_128), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_155), .A2(n_126), .B1(n_120), .B2(n_83), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_175), .B(n_101), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_195), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_155), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_164), .B(n_2), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_180), .B(n_91), .Y(n_253) );
OR2x2_ASAP7_75t_SL g254 ( .A(n_192), .B(n_148), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_186), .B(n_84), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_160), .B(n_84), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_181), .B(n_130), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_182), .B(n_130), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_212), .B(n_192), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_209), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_237), .B(n_198), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_229), .B(n_148), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_205), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_209), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_214), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_219), .B(n_4), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_214), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_233), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_206), .B(n_148), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_233), .Y(n_274) );
INVx3_ASAP7_75t_SL g275 ( .A(n_239), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_219), .B(n_5), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_215), .A2(n_203), .B(n_157), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_237), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_214), .B(n_118), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_206), .B(n_118), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_215), .A2(n_203), .B(n_157), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_208), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_210), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_208), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_251), .A2(n_118), .B1(n_130), .B2(n_184), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_226), .A2(n_130), .B1(n_201), .B2(n_173), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_220), .A2(n_184), .B(n_201), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_234), .B(n_5), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_247), .A2(n_130), .B1(n_162), .B2(n_194), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_246), .B(n_130), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_204), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_204), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_243), .A2(n_162), .B1(n_165), .B2(n_194), .Y(n_296) );
BUFx4_ASAP7_75t_SL g297 ( .A(n_239), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_218), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_246), .B(n_6), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_218), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_248), .B(n_165), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_217), .Y(n_303) );
OR2x6_ASAP7_75t_L g304 ( .A(n_268), .B(n_239), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_275), .A2(n_231), .B1(n_223), .B2(n_211), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_268), .A2(n_228), .B1(n_207), .B2(n_242), .Y(n_306) );
NAND3x1_ASAP7_75t_L g307 ( .A(n_297), .B(n_222), .C(n_256), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_302), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_284), .B(n_250), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_268), .A2(n_207), .B1(n_242), .B2(n_243), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_268), .A2(n_207), .B1(n_255), .B2(n_256), .Y(n_312) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_276), .B(n_227), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_283), .B(n_227), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_265), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_297), .Y(n_316) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_290), .B(n_213), .C(n_252), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_283), .B(n_232), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_293), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_265), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_275), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g322 ( .A1(n_276), .A2(n_252), .B1(n_222), .B2(n_217), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_270), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_270), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_278), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_284), .B(n_232), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_282), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_299), .B(n_242), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_277), .A2(n_236), .B(n_225), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_309), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_313), .B(n_276), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_313), .B(n_276), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_313), .A2(n_303), .B1(n_290), .B2(n_299), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_331), .A2(n_264), .B(n_281), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_325), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_305), .A2(n_255), .B1(n_230), .B2(n_213), .C(n_221), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_310), .A2(n_221), .B1(n_259), .B2(n_287), .C(n_300), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_325), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_312), .B(n_304), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_304), .A2(n_275), .B1(n_263), .B2(n_303), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_329), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_312), .B(n_259), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_306), .B(n_287), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_304), .A2(n_263), .B1(n_291), .B2(n_261), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_304), .A2(n_263), .B1(n_295), .B2(n_249), .Y(n_349) );
AOI21x1_ASAP7_75t_L g350 ( .A1(n_332), .A2(n_295), .B(n_264), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_263), .B1(n_291), .B2(n_295), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_308), .B(n_263), .Y(n_353) );
AOI222xp33_ASAP7_75t_L g354 ( .A1(n_317), .A2(n_300), .B1(n_278), .B2(n_244), .C1(n_241), .C2(n_253), .Y(n_354) );
OAI211xp5_ASAP7_75t_L g355 ( .A1(n_322), .A2(n_249), .B(n_292), .C(n_280), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_311), .A2(n_292), .B1(n_285), .B2(n_272), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_315), .B(n_260), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_334), .A2(n_346), .B1(n_343), .B2(n_335), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_345), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_333), .B(n_328), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_343), .A2(n_318), .B1(n_328), .B2(n_327), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_352), .Y(n_363) );
AO31x2_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_277), .A3(n_281), .B(n_315), .Y(n_364) );
BUFx8_ASAP7_75t_SL g365 ( .A(n_335), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_350), .A2(n_273), .B(n_286), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_340), .A2(n_330), .B1(n_328), .B2(n_318), .C(n_327), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_333), .B(n_320), .Y(n_368) );
NAND3xp33_ASAP7_75t_L g369 ( .A(n_354), .B(n_273), .C(n_296), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_354), .A2(n_318), .B1(n_328), .B2(n_314), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_355), .A2(n_318), .A3(n_314), .B(n_216), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_352), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_337), .B(n_321), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_350), .A2(n_286), .B(n_280), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_346), .A2(n_316), .B1(n_272), .B2(n_274), .Y(n_377) );
AO21x2_ASAP7_75t_L g378 ( .A1(n_351), .A2(n_332), .B(n_289), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_339), .B(n_320), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_342), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_336), .A2(n_316), .B(n_321), .C(n_307), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_288), .B1(n_285), .B2(n_258), .C(n_274), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_342), .B(n_341), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_347), .A2(n_289), .B(n_258), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_352), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_356), .B(n_307), .C(n_257), .D(n_329), .Y(n_386) );
AOI31xp33_ASAP7_75t_L g387 ( .A1(n_334), .A2(n_326), .A3(n_324), .B(n_323), .Y(n_387) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_351), .A2(n_326), .B1(n_324), .B2(n_323), .C1(n_261), .C2(n_260), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_385), .B(n_357), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_385), .B(n_363), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_363), .B(n_357), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_363), .B(n_353), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_371), .B(n_353), .Y(n_394) );
OAI33xp33_ASAP7_75t_L g395 ( .A1(n_374), .A2(n_348), .A3(n_193), .B1(n_178), .B2(n_173), .B3(n_167), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_365), .Y(n_396) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_387), .B(n_319), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_373), .B(n_319), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
INVx4_ASAP7_75t_L g401 ( .A(n_387), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
OAI22xp5_ASAP7_75t_SL g403 ( .A1(n_361), .A2(n_344), .B1(n_235), .B2(n_319), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_279), .B1(n_271), .B2(n_269), .C(n_262), .Y(n_405) );
AOI221x1_ASAP7_75t_L g406 ( .A1(n_386), .A2(n_319), .B1(n_267), .B2(n_266), .C(n_262), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_319), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_386), .A2(n_167), .A3(n_178), .B1(n_193), .B2(n_9), .B3(n_10), .Y(n_408) );
NAND2xp33_ASAP7_75t_SL g409 ( .A(n_358), .B(n_293), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_373), .B(n_262), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_372), .B(n_293), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_371), .B(n_262), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_375), .B(n_266), .Y(n_413) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_388), .B(n_266), .Y(n_414) );
NAND2x1_ASAP7_75t_L g415 ( .A(n_375), .B(n_266), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_368), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_379), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_380), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_379), .Y(n_420) );
OAI31xp33_ASAP7_75t_L g421 ( .A1(n_381), .A2(n_282), .A3(n_269), .B(n_271), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_358), .B(n_383), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_360), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_378), .B(n_364), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_378), .B(n_267), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_364), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_369), .B(n_269), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_364), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_378), .B(n_267), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_364), .Y(n_432) );
AOI221x1_ASAP7_75t_L g433 ( .A1(n_369), .A2(n_267), .B1(n_269), .B2(n_271), .C(n_179), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_424), .B(n_364), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_424), .B(n_364), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_426), .B(n_366), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_402), .Y(n_439) );
NAND2x1_ASAP7_75t_SL g440 ( .A(n_401), .B(n_271), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_390), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_426), .B(n_366), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_430), .B(n_366), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_390), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_398), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_416), .B(n_370), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_417), .B(n_384), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_408), .B(n_367), .C(n_382), .Y(n_449) );
AND4x1_ASAP7_75t_L g450 ( .A(n_396), .B(n_377), .C(n_7), .D(n_8), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_420), .B(n_384), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_420), .B(n_366), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_425), .B(n_179), .C(n_183), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_400), .Y(n_454) );
NOR2xp33_ASAP7_75t_R g455 ( .A(n_396), .B(n_6), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
NOR2xp33_ASAP7_75t_SL g457 ( .A(n_401), .B(n_279), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_430), .B(n_376), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_432), .B(n_376), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_403), .A2(n_376), .B1(n_293), .B2(n_294), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_397), .B(n_53), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_389), .B(n_7), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_389), .B(n_11), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_422), .B(n_394), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_397), .B(n_55), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_404), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_404), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_418), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_418), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_419), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_403), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_422), .A2(n_293), .B1(n_294), .B2(n_298), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_419), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g474 ( .A1(n_425), .A2(n_12), .A3(n_14), .B1(n_15), .B2(n_17), .B3(n_18), .Y(n_474) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_401), .B(n_294), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_432), .B(n_12), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_394), .B(n_14), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_427), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_423), .B(n_15), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_401), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_392), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_392), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_423), .B(n_17), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_393), .B(n_191), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_432), .B(n_202), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_450), .B(n_395), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_453), .A2(n_409), .B(n_433), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_466), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_466), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_439), .B(n_393), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_471), .B(n_412), .Y(n_492) );
OAI21xp33_ASAP7_75t_SL g493 ( .A1(n_440), .A2(n_414), .B(n_421), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_482), .B(n_429), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_471), .A2(n_421), .B1(n_428), .B2(n_414), .C(n_429), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_440), .A2(n_415), .B(n_405), .C(n_411), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_474), .A2(n_429), .B1(n_427), .B2(n_431), .C(n_412), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_480), .A2(n_406), .B(n_433), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_449), .B(n_406), .C(n_413), .D(n_410), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_457), .A2(n_415), .B(n_428), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_446), .A2(n_428), .B1(n_410), .B2(n_407), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_483), .B(n_407), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_464), .B(n_399), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_460), .A2(n_399), .B(n_293), .Y(n_505) );
AOI21xp33_ASAP7_75t_SL g506 ( .A1(n_481), .A2(n_20), .B(n_21), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
OAI221xp5_ASAP7_75t_SL g508 ( .A1(n_480), .A2(n_282), .B1(n_298), .B2(n_301), .C(n_202), .Y(n_508) );
NAND3xp33_ASAP7_75t_SL g509 ( .A(n_455), .B(n_301), .C(n_298), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_484), .A2(n_202), .B(n_196), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_441), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_435), .B(n_188), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_475), .A2(n_301), .B(n_179), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_445), .Y(n_514) );
AND2x2_ASAP7_75t_SL g515 ( .A(n_461), .B(n_22), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_481), .A2(n_185), .B1(n_188), .B2(n_191), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_444), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_435), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_484), .A2(n_189), .B1(n_183), .B2(n_179), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_445), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_448), .A2(n_189), .B1(n_183), .B2(n_179), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_448), .A2(n_196), .B1(n_191), .B2(n_188), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_438), .B(n_196), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_454), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g526 ( .A1(n_478), .A2(n_185), .B(n_189), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_476), .B(n_189), .C(n_183), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
AOI21xp33_ASAP7_75t_SL g530 ( .A1(n_461), .A2(n_23), .B(n_31), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_438), .B(n_32), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_469), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_456), .Y(n_533) );
OAI211xp5_ASAP7_75t_L g534 ( .A1(n_462), .A2(n_185), .B(n_189), .C(n_183), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_509), .B(n_463), .Y(n_535) );
O2A1O1Ixp5_ASAP7_75t_L g536 ( .A1(n_487), .A2(n_461), .B(n_465), .C(n_476), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_503), .B(n_434), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_511), .Y(n_538) );
INVxp33_ASAP7_75t_L g539 ( .A(n_509), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_491), .B(n_434), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_492), .B(n_436), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_529), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_518), .B(n_436), .Y(n_543) );
XNOR2x2_ASAP7_75t_L g544 ( .A(n_495), .B(n_452), .Y(n_544) );
O2A1O1Ixp5_ASAP7_75t_L g545 ( .A1(n_508), .A2(n_465), .B(n_451), .C(n_473), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_517), .B(n_458), .Y(n_546) );
NAND2xp33_ASAP7_75t_SL g547 ( .A(n_494), .B(n_465), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_493), .A2(n_458), .B(n_459), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_521), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_515), .A2(n_486), .B(n_459), .Y(n_550) );
AOI221x1_ASAP7_75t_L g551 ( .A1(n_499), .A2(n_479), .B1(n_477), .B2(n_486), .C(n_473), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_529), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_525), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_502), .B(n_437), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_501), .A2(n_437), .B1(n_442), .B2(n_443), .Y(n_555) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_528), .B(n_443), .Y(n_556) );
AOI322xp5_ASAP7_75t_L g557 ( .A1(n_497), .A2(n_442), .A3(n_456), .B1(n_470), .B2(n_479), .C1(n_472), .C2(n_485), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_532), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_489), .B(n_470), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_490), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_504), .Y(n_561) );
NOR4xp25_ASAP7_75t_SL g562 ( .A(n_513), .B(n_485), .C(n_35), .D(n_37), .Y(n_562) );
NOR4xp75_ASAP7_75t_L g563 ( .A(n_498), .B(n_34), .C(n_41), .D(n_43), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_507), .B(n_189), .Y(n_564) );
AND2x6_ASAP7_75t_L g565 ( .A(n_531), .B(n_505), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_533), .B(n_44), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_514), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_541), .B(n_508), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_554), .B(n_520), .Y(n_569) );
AOI322xp5_ASAP7_75t_L g570 ( .A1(n_541), .A2(n_519), .A3(n_510), .B1(n_496), .B2(n_522), .C1(n_512), .C2(n_524), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g571 ( .A1(n_556), .A2(n_527), .B(n_534), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g572 ( .A1(n_536), .A2(n_530), .B(n_506), .C(n_526), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_552), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_548), .B(n_500), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_542), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_538), .Y(n_576) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_565), .B(n_500), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_549), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_557), .B(n_534), .C(n_488), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_567), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_555), .A2(n_516), .B(n_523), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_537), .B(n_488), .Y(n_582) );
NOR3xp33_ASAP7_75t_L g583 ( .A(n_536), .B(n_245), .C(n_240), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_553), .Y(n_584) );
AOI322xp5_ASAP7_75t_L g585 ( .A1(n_540), .A2(n_183), .A3(n_51), .B1(n_52), .B2(n_56), .C1(n_60), .C2(n_63), .Y(n_585) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_543), .Y(n_586) );
XNOR2x1_ASAP7_75t_L g587 ( .A(n_544), .B(n_46), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_587), .A2(n_565), .B1(n_535), .B2(n_547), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_582), .B(n_546), .Y(n_589) );
NOR4xp25_ASAP7_75t_L g590 ( .A(n_579), .B(n_535), .C(n_558), .D(n_550), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_587), .A2(n_539), .B1(n_560), .B2(n_561), .Y(n_591) );
NAND4xp75_ASAP7_75t_L g592 ( .A(n_574), .B(n_551), .C(n_545), .D(n_566), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_576), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_573), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_568), .A2(n_565), .B1(n_539), .B2(n_559), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_574), .B(n_565), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_577), .B(n_565), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_568), .A2(n_545), .B(n_564), .C(n_562), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_571), .A2(n_563), .B(n_67), .C(n_224), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_586), .A2(n_224), .B1(n_578), .B2(n_584), .C(n_581), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_572), .A2(n_224), .B(n_575), .Y(n_601) );
NOR4xp25_ASAP7_75t_L g602 ( .A(n_573), .B(n_575), .C(n_580), .D(n_569), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_580), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g604 ( .A(n_570), .B(n_583), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_585), .B(n_537), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_593), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_591), .A2(n_604), .B1(n_595), .B2(n_596), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_597), .B(n_589), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_597), .A2(n_601), .B1(n_605), .B2(n_594), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_606), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_608), .Y(n_611) );
OAI222xp33_ASAP7_75t_L g612 ( .A1(n_611), .A2(n_607), .B1(n_609), .B2(n_588), .C1(n_590), .C2(n_603), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_610), .Y(n_613) );
XNOR2xp5_ASAP7_75t_L g614 ( .A(n_613), .B(n_611), .Y(n_614) );
AOI222xp33_ASAP7_75t_L g615 ( .A1(n_614), .A2(n_613), .B1(n_612), .B2(n_600), .C1(n_602), .C2(n_592), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_615), .A2(n_598), .B(n_599), .Y(n_616) );
endmodule