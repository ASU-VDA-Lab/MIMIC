module real_aes_2350_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_0), .B(n_176), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_1), .A2(n_184), .B(n_206), .Y(n_205) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_2), .A2(n_55), .B1(n_90), .B2(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_3), .B(n_191), .Y(n_254) );
INVx1_ASAP7_75t_L g160 ( .A(n_4), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g143 ( .A1(n_5), .A2(n_144), .B1(n_145), .B2(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g146 ( .A(n_5), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_6), .B(n_191), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_7), .A2(n_26), .B1(n_136), .B2(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g145 ( .A(n_8), .Y(n_145) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_9), .A2(n_25), .B1(n_90), .B2(n_98), .Y(n_97) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_10), .A2(n_20), .B1(n_133), .B2(n_134), .Y(n_132) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_11), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g173 ( .A(n_12), .Y(n_173) );
AOI221x1_ASAP7_75t_L g270 ( .A1(n_13), .A2(n_21), .B1(n_176), .B2(n_184), .C(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_14), .B(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_15), .A2(n_171), .B(n_174), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_16), .B(n_209), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_17), .A2(n_60), .B1(n_125), .B2(n_126), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_18), .B(n_191), .Y(n_218) );
INVx1_ASAP7_75t_L g492 ( .A(n_18), .Y(n_492) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_19), .A2(n_176), .B(n_250), .Y(n_249) );
NAND2x1_ASAP7_75t_L g240 ( .A(n_22), .B(n_191), .Y(n_240) );
NAND2x1_ASAP7_75t_L g228 ( .A(n_23), .B(n_193), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_24), .A2(n_39), .B1(n_112), .B2(n_116), .Y(n_111) );
OAI221xp5_ASAP7_75t_L g152 ( .A1(n_25), .A2(n_55), .B1(n_59), .B2(n_153), .C(n_155), .Y(n_152) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_27), .A2(n_67), .B(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g196 ( .A(n_27), .B(n_67), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_28), .A2(n_66), .B1(n_119), .B2(n_120), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_29), .B(n_193), .Y(n_208) );
INVx3_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_31), .A2(n_81), .B1(n_82), .B2(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_31), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_32), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_33), .B(n_193), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_34), .A2(n_184), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_SL g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g162 ( .A(n_36), .Y(n_162) );
AND2x2_ASAP7_75t_L g182 ( .A(n_36), .B(n_160), .Y(n_182) );
AND2x2_ASAP7_75t_L g185 ( .A(n_36), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_37), .B(n_176), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_38), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_40), .B(n_193), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_41), .A2(n_64), .B1(n_103), .B2(n_108), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_42), .A2(n_63), .B1(n_129), .B2(n_130), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_43), .A2(n_184), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_44), .B(n_86), .Y(n_85) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_45), .A2(n_59), .B1(n_90), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_46), .B(n_193), .Y(n_241) );
INVx1_ASAP7_75t_L g179 ( .A(n_47), .Y(n_179) );
INVx1_ASAP7_75t_L g188 ( .A(n_47), .Y(n_188) );
INVx1_ASAP7_75t_L g92 ( .A(n_48), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_49), .B(n_191), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_50), .A2(n_184), .B(n_239), .Y(n_238) );
AO21x1_ASAP7_75t_L g251 ( .A1(n_51), .A2(n_184), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_52), .B(n_176), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_53), .B(n_176), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_54), .A2(n_141), .B1(n_142), .B2(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_54), .Y(n_141) );
INVxp33_ASAP7_75t_L g157 ( .A(n_55), .Y(n_157) );
AND2x2_ASAP7_75t_L g264 ( .A(n_56), .B(n_210), .Y(n_264) );
INVx1_ASAP7_75t_L g181 ( .A(n_57), .Y(n_181) );
INVx1_ASAP7_75t_L g186 ( .A(n_57), .Y(n_186) );
AND2x2_ASAP7_75t_L g232 ( .A(n_58), .B(n_201), .Y(n_232) );
INVxp67_ASAP7_75t_L g156 ( .A(n_59), .Y(n_156) );
AND2x2_ASAP7_75t_L g200 ( .A(n_61), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_62), .B(n_176), .Y(n_220) );
INVx1_ASAP7_75t_L g513 ( .A(n_62), .Y(n_513) );
AND2x2_ASAP7_75t_L g250 ( .A(n_65), .B(n_195), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_68), .B(n_193), .Y(n_219) );
AND2x2_ASAP7_75t_L g244 ( .A(n_69), .B(n_201), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_70), .B(n_191), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_71), .A2(n_184), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_72), .B(n_193), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_73), .A2(n_140), .B1(n_147), .B2(n_148), .Y(n_139) );
INVx1_ASAP7_75t_L g147 ( .A(n_73), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_73), .B(n_191), .Y(n_207) );
BUFx2_ASAP7_75t_L g80 ( .A(n_74), .Y(n_80) );
BUFx2_ASAP7_75t_SL g154 ( .A(n_75), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_76), .A2(n_184), .B(n_189), .Y(n_183) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_149), .B1(n_163), .B2(n_485), .C(n_489), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_139), .Y(n_78) );
AOI22xp33_ASAP7_75t_SL g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_138), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_80), .Y(n_138) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_81), .A2(n_82), .B1(n_491), .B2(n_492), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
OR2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_123), .Y(n_83) );
NAND4xp25_ASAP7_75t_SL g84 ( .A(n_85), .B(n_102), .C(n_111), .D(n_118), .Y(n_84) );
AND2x4_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x2_ASAP7_75t_L g108 ( .A(n_87), .B(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g116 ( .A(n_87), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g106 ( .A(n_88), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g114 ( .A(n_88), .Y(n_114) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_88), .Y(n_121) );
OAI22x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g98 ( .A(n_90), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_90), .Y(n_101) );
INVx2_ASAP7_75t_L g107 ( .A(n_93), .Y(n_107) );
AND2x2_ASAP7_75t_L g113 ( .A(n_93), .B(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
AND2x2_ASAP7_75t_L g129 ( .A(n_95), .B(n_106), .Y(n_129) );
AND2x6_ASAP7_75t_L g134 ( .A(n_95), .B(n_113), .Y(n_134) );
AND2x2_ASAP7_75t_L g136 ( .A(n_95), .B(n_131), .Y(n_136) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g105 ( .A(n_97), .Y(n_105) );
AND2x4_ASAP7_75t_L g115 ( .A(n_97), .B(n_99), .Y(n_115) );
AND2x2_ASAP7_75t_L g122 ( .A(n_97), .B(n_100), .Y(n_122) );
INVxp67_ASAP7_75t_L g117 ( .A(n_99), .Y(n_117) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g104 ( .A(n_100), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g125 ( .A(n_104), .B(n_113), .Y(n_125) );
AND2x6_ASAP7_75t_L g137 ( .A(n_104), .B(n_131), .Y(n_137) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_105), .Y(n_110) );
AND2x4_ASAP7_75t_L g119 ( .A(n_106), .B(n_115), .Y(n_119) );
AND2x4_ASAP7_75t_L g131 ( .A(n_107), .B(n_114), .Y(n_131) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g133 ( .A(n_115), .B(n_131), .Y(n_133) );
AND2x2_ASAP7_75t_SL g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x4_ASAP7_75t_L g126 ( .A(n_122), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g130 ( .A(n_122), .B(n_131), .Y(n_130) );
NAND4xp25_ASAP7_75t_SL g123 ( .A(n_124), .B(n_128), .C(n_132), .D(n_135), .Y(n_123) );
INVx1_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_150), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_151), .Y(n_150) );
AND3x1_ASAP7_75t_SL g151 ( .A(n_152), .B(n_158), .C(n_161), .Y(n_151) );
INVxp67_ASAP7_75t_L g498 ( .A(n_152), .Y(n_498) );
CKINVDCx8_ASAP7_75t_R g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_158), .Y(n_496) );
AO21x1_ASAP7_75t_SL g506 ( .A1(n_158), .A2(n_507), .B(n_511), .Y(n_506) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OR2x2_ASAP7_75t_SL g503 ( .A(n_159), .B(n_161), .Y(n_503) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g187 ( .A(n_160), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_161), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2x1p5_ASAP7_75t_L g508 ( .A(n_162), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_406), .Y(n_164) );
NOR3xp33_ASAP7_75t_SL g165 ( .A(n_166), .B(n_318), .C(n_358), .Y(n_165) );
OAI221xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_233), .B1(n_282), .B2(n_297), .C(n_300), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_197), .Y(n_168) );
INVx2_ASAP7_75t_L g315 ( .A(n_169), .Y(n_315) );
AND2x2_ASAP7_75t_L g345 ( .A(n_169), .B(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g283 ( .A(n_170), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g290 ( .A(n_170), .B(n_223), .Y(n_290) );
INVx2_ASAP7_75t_L g296 ( .A(n_170), .Y(n_296) );
AND2x2_ASAP7_75t_L g305 ( .A(n_170), .B(n_199), .Y(n_305) );
INVx1_ASAP7_75t_L g321 ( .A(n_170), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_170), .B(n_367), .Y(n_366) );
BUFx4f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
AND2x4_ASAP7_75t_L g195 ( .A(n_173), .B(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_173), .B(n_196), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_183), .B(n_195), .Y(n_174) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_176), .Y(n_488) );
AND2x4_ASAP7_75t_L g176 ( .A(n_177), .B(n_182), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
AND2x6_ASAP7_75t_L g193 ( .A(n_178), .B(n_186), .Y(n_193) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g191 ( .A(n_180), .B(n_188), .Y(n_191) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx5_ASAP7_75t_L g194 ( .A(n_182), .Y(n_194) );
AND2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_187), .Y(n_184) );
INVx2_ASAP7_75t_L g510 ( .A(n_186), .Y(n_510) );
INVx2_ASAP7_75t_L g512 ( .A(n_188), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B(n_194), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_194), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_194), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_194), .A2(n_253), .B(n_254), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_194), .A2(n_261), .B(n_262), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_194), .A2(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_SL g214 ( .A(n_195), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_195), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_198), .B(n_211), .Y(n_197) );
INVx4_ASAP7_75t_L g286 ( .A(n_198), .Y(n_286) );
AND2x2_ASAP7_75t_L g317 ( .A(n_198), .B(n_224), .Y(n_317) );
AND2x2_ASAP7_75t_L g393 ( .A(n_198), .B(n_367), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_198), .B(n_223), .Y(n_435) );
INVx5_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_199), .B(n_223), .Y(n_322) );
AND2x2_ASAP7_75t_L g346 ( .A(n_199), .B(n_224), .Y(n_346) );
BUFx2_ASAP7_75t_L g362 ( .A(n_199), .Y(n_362) );
NOR2x1_ASAP7_75t_SL g465 ( .A(n_199), .B(n_367), .Y(n_465) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_203), .Y(n_199) );
INVx3_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_209), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_209), .Y(n_231) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_209), .A2(n_270), .B(n_274), .Y(n_269) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_209), .A2(n_270), .B(n_274), .Y(n_332) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g342 ( .A(n_211), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_211), .A2(n_409), .B1(n_411), .B2(n_413), .C(n_418), .Y(n_408) );
AND2x2_ASAP7_75t_L g428 ( .A(n_211), .B(n_321), .Y(n_428) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
INVx1_ASAP7_75t_L g337 ( .A(n_213), .Y(n_337) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_214), .B(n_222), .Y(n_221) );
AO21x2_ASAP7_75t_L g367 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_223), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g306 ( .A(n_223), .B(n_294), .Y(n_306) );
INVx2_ASAP7_75t_L g348 ( .A(n_223), .Y(n_348) );
AND2x2_ASAP7_75t_L g481 ( .A(n_223), .B(n_296), .Y(n_481) );
INVx4_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_224), .Y(n_338) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_231), .B(n_232), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_230), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_265), .C(n_280), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_245), .Y(n_234) );
INVx2_ASAP7_75t_L g395 ( .A(n_235), .Y(n_395) );
AND2x2_ASAP7_75t_L g440 ( .A(n_235), .B(n_317), .Y(n_440) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g385 ( .A(n_236), .Y(n_385) );
AND2x4_ASAP7_75t_SL g400 ( .A(n_236), .B(n_312), .Y(n_400) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_243), .B(n_244), .Y(n_236) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_237), .A2(n_243), .B(n_244), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_243), .A2(n_258), .B(n_264), .Y(n_257) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_243), .A2(n_258), .B(n_264), .Y(n_277) );
INVx2_ASAP7_75t_L g354 ( .A(n_245), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_245), .B(n_384), .Y(n_410) );
AND2x4_ASAP7_75t_L g443 ( .A(n_245), .B(n_390), .Y(n_443) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_257), .Y(n_245) );
AND2x2_ASAP7_75t_L g281 ( .A(n_246), .B(n_276), .Y(n_281) );
OR2x2_ASAP7_75t_L g311 ( .A(n_246), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_246), .B(n_332), .Y(n_380) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx2_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g299 ( .A(n_248), .Y(n_299) );
OAI21x1_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_251), .B(n_255), .Y(n_248) );
INVx1_ASAP7_75t_L g256 ( .A(n_250), .Y(n_256) );
INVx2_ASAP7_75t_L g312 ( .A(n_257), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_259), .B(n_263), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_265), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_275), .Y(n_266) );
AND2x2_ASAP7_75t_L g280 ( .A(n_267), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g353 ( .A(n_267), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g438 ( .A(n_267), .Y(n_438) );
BUFx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g298 ( .A(n_268), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g417 ( .A(n_268), .B(n_277), .Y(n_417) );
AND2x2_ASAP7_75t_L g421 ( .A(n_268), .B(n_287), .Y(n_421) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g390 ( .A(n_269), .Y(n_390) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_269), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_275), .B(n_298), .Y(n_374) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_276), .B(n_299), .Y(n_484) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g288 ( .A(n_277), .B(n_279), .Y(n_288) );
AND2x2_ASAP7_75t_L g370 ( .A(n_277), .B(n_332), .Y(n_370) );
AND2x2_ASAP7_75t_L g389 ( .A(n_277), .B(n_278), .Y(n_389) );
BUFx2_ASAP7_75t_L g310 ( .A(n_278), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_278), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx3_ASAP7_75t_L g287 ( .A(n_279), .Y(n_287) );
INVxp67_ASAP7_75t_L g330 ( .A(n_279), .Y(n_330) );
INVx1_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
AND2x2_ASAP7_75t_L g339 ( .A(n_281), .B(n_310), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g420 ( .A(n_281), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g457 ( .A(n_281), .B(n_458), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B1(n_288), .B2(n_289), .C(n_291), .Y(n_282) );
AND2x2_ASAP7_75t_L g386 ( .A(n_283), .B(n_286), .Y(n_386) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_283), .B(n_346), .Y(n_405) );
AND2x2_ASAP7_75t_L g423 ( .A(n_283), .B(n_348), .Y(n_423) );
AND2x2_ASAP7_75t_L g478 ( .A(n_283), .B(n_317), .Y(n_478) );
INVx1_ASAP7_75t_L g294 ( .A(n_284), .Y(n_294) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_284), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_285), .Y(n_430) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_286), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_286), .B(n_337), .Y(n_412) );
AND2x2_ASAP7_75t_L g379 ( .A(n_287), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g415 ( .A(n_287), .Y(n_415) );
AND2x2_ASAP7_75t_L g324 ( .A(n_288), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_288), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g466 ( .A(n_288), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_288), .B(n_390), .Y(n_476) );
AND2x4_ASAP7_75t_L g392 ( .A(n_289), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g463 ( .A(n_290), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
OR2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g341 ( .A(n_296), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g372 ( .A(n_296), .B(n_346), .Y(n_372) );
AND2x2_ASAP7_75t_L g446 ( .A(n_296), .B(n_367), .Y(n_446) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g394 ( .A(n_298), .B(n_395), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g459 ( .A1(n_298), .A2(n_460), .A3(n_462), .B1(n_463), .B2(n_466), .Y(n_459) );
AND2x4_ASAP7_75t_L g331 ( .A(n_299), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g429 ( .A(n_299), .B(n_332), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B1(n_307), .B2(n_313), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_SL g418 ( .A1(n_302), .A2(n_316), .B(n_419), .C(n_420), .Y(n_418) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g402 ( .A(n_303), .B(n_330), .Y(n_402) );
INVx1_ASAP7_75t_SL g473 ( .A(n_304), .Y(n_473) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x4_ASAP7_75t_L g376 ( .A(n_306), .B(n_315), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_306), .A2(n_455), .B1(n_456), .B2(n_457), .C(n_459), .Y(n_454) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_311), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_314), .A2(n_344), .B1(n_397), .B2(n_398), .Y(n_396) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_315), .A2(n_433), .B(n_441), .C(n_454), .Y(n_432) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g352 ( .A(n_317), .B(n_321), .Y(n_352) );
OAI211xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_323), .B(n_326), .C(n_355), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g349 ( .A(n_321), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g469 ( .A(n_321), .B(n_465), .Y(n_469) );
OAI32xp33_ASAP7_75t_L g426 ( .A1(n_322), .A2(n_427), .A3(n_429), .B1(n_430), .B2(n_431), .Y(n_426) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_325), .B(n_417), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_333), .B1(n_339), .B2(n_340), .C(n_343), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g483 ( .A(n_330), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_331), .B(n_395), .Y(n_397) );
A2O1A1O1Ixp25_ASAP7_75t_L g468 ( .A1(n_331), .A2(n_400), .B(n_416), .C(n_462), .D(n_469), .Y(n_468) );
AOI31xp33_ASAP7_75t_L g470 ( .A1(n_331), .A2(n_352), .A3(n_462), .B(n_469), .Y(n_470) );
AND2x2_ASAP7_75t_L g384 ( .A(n_332), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_334), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx2_ASAP7_75t_L g461 ( .A(n_336), .Y(n_461) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g456 ( .A(n_337), .B(n_348), .Y(n_456) );
INVx1_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
AND2x2_ASAP7_75t_L g356 ( .A(n_340), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI31xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .A3(n_351), .B(n_353), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_346), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g479 ( .A(n_346), .B(n_425), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g424 ( .A(n_348), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g450 ( .A(n_348), .Y(n_450) );
INVxp67_ASAP7_75t_L g419 ( .A(n_349), .Y(n_419) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g357 ( .A(n_353), .Y(n_357) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g358 ( .A(n_359), .B(n_375), .C(n_391), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_368), .B1(n_372), .B2(n_373), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_L g445 ( .A(n_362), .Y(n_445) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_366), .Y(n_425) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_366), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_366), .B(n_435), .Y(n_452) );
NAND2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g403 ( .A(n_370), .Y(n_403) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_386), .B2(n_387), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_378), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_384), .A2(n_389), .B1(n_423), .B2(n_424), .C(n_426), .Y(n_422) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g462 ( .A(n_389), .Y(n_462) );
AND2x2_ASAP7_75t_L g399 ( .A(n_390), .B(n_400), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_SL g447 ( .A1(n_390), .A2(n_448), .B(n_452), .C(n_453), .Y(n_447) );
AOI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_396), .C(n_401), .Y(n_391) );
AND2x2_ASAP7_75t_L g442 ( .A(n_395), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
AOI21xp33_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_403), .B(n_404), .Y(n_401) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_432), .C(n_467), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_408), .B(n_422), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g431 ( .A(n_416), .Y(n_431) );
INVxp67_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g439 ( .A(n_429), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_439), .B2(n_440), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .B(n_447), .Y(n_441) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g480 ( .A(n_465), .B(n_481), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B1(n_471), .B2(n_474), .C(n_477), .Y(n_467) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI31xp33_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_479), .A3(n_480), .B(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI222xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B1(n_499), .B2(n_501), .C1(n_504), .C2(n_513), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
endmodule