module fake_netlist_6_3239_n_107 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_107);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;

output n_107;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_93;
wire n_40;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx2_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

AND3x1_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_4),
.C(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_6),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_25),
.B1(n_32),
.B2(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_30),
.Y(n_50)
);

OR2x6_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_25),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_27),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_41),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_52),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_51),
.B1(n_42),
.B2(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_57),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_48),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_48),
.B1(n_56),
.B2(n_52),
.Y(n_73)
);

AND2x6_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_70),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_64),
.B(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_73),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_82),
.Y(n_94)
);

NAND2x1_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_24),
.Y(n_97)
);

NOR4xp25_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_24),
.C(n_32),
.D(n_26),
.Y(n_98)
);

AOI221x1_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_26),
.B1(n_40),
.B2(n_39),
.C(n_51),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_40),
.Y(n_100)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_33),
.B1(n_68),
.B2(n_55),
.C(n_54),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_63),
.C(n_95),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_100),
.B(n_99),
.Y(n_103)
);

NAND3x1_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_101),
.C(n_51),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_51),
.B1(n_100),
.B2(n_63),
.Y(n_105)
);

OAI222xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_63),
.B1(n_10),
.B2(n_56),
.C1(n_55),
.C2(n_16),
.Y(n_106)
);

AOI31xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_10),
.A3(n_56),
.B(n_15),
.Y(n_107)
);


endmodule