module fake_jpeg_32195_n_456 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_456);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_456;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_90),
.Y(n_102)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_62),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_70),
.Y(n_98)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_78),
.Y(n_111)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_17),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_36),
.B(n_14),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_91),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_13),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_100),
.B(n_134),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_49),
.A2(n_19),
.B(n_23),
.C(n_38),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_29),
.C(n_38),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_44),
.B1(n_43),
.B2(n_39),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_66),
.B1(n_89),
.B2(n_83),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_77),
.A2(n_43),
.B1(n_44),
.B2(n_33),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_55),
.B1(n_81),
.B2(n_75),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_53),
.B(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_49),
.B(n_27),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_27),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_62),
.B(n_21),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_65),
.B(n_21),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_102),
.Y(n_150)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_23),
.B1(n_33),
.B2(n_38),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_170),
.B1(n_185),
.B2(n_187),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_150),
.B(n_151),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_69),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_157),
.Y(n_198)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_33),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_91),
.B1(n_74),
.B2(n_52),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_130),
.B1(n_125),
.B2(n_120),
.Y(n_190)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_159),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_166),
.B1(n_176),
.B2(n_107),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_40),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_163),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_40),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_169),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_123),
.A2(n_45),
.B1(n_50),
.B2(n_92),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_174),
.Y(n_202)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_57),
.B1(n_72),
.B2(n_79),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_178),
.Y(n_208)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_181),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_99),
.B(n_29),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_34),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_61),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_131),
.A2(n_92),
.B1(n_47),
.B2(n_51),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_119),
.A2(n_43),
.B1(n_44),
.B2(n_29),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_139),
.C(n_110),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_192),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_197),
.B1(n_205),
.B2(n_176),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_126),
.C(n_60),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_209),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_152),
.A2(n_158),
.B1(n_182),
.B2(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_180),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_158),
.A2(n_141),
.B1(n_107),
.B2(n_120),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_125),
.B1(n_118),
.B2(n_96),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_225),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_218),
.B(n_227),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_222),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_156),
.B1(n_164),
.B2(n_137),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_224),
.B(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_154),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_151),
.B(n_137),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_239),
.B(n_206),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_159),
.B1(n_121),
.B2(n_97),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_161),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_121),
.B1(n_97),
.B2(n_113),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_230),
.Y(n_253)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_167),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_199),
.B1(n_189),
.B2(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_197),
.A2(n_118),
.B1(n_155),
.B2(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_194),
.B1(n_192),
.B2(n_212),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_202),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_172),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_238),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_190),
.B1(n_206),
.B2(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_199),
.B(n_99),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_177),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_251),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_250),
.B1(n_263),
.B2(n_235),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_260),
.B(n_263),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_242),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_206),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_266),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_199),
.B1(n_216),
.B2(n_213),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_255),
.A2(n_256),
.B1(n_235),
.B2(n_234),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_213),
.B1(n_212),
.B2(n_195),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_259),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_208),
.B(n_201),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_195),
.B1(n_208),
.B2(n_193),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_262),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_207),
.C(n_211),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_227),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_271),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_285),
.B(n_287),
.Y(n_301)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_281),
.Y(n_303)
);

AO22x1_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_239),
.B1(n_229),
.B2(n_234),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_276),
.A2(n_296),
.B(n_224),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_278),
.B1(n_290),
.B2(n_255),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_279),
.A2(n_261),
.B1(n_253),
.B2(n_219),
.Y(n_318)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_222),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_284),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_244),
.B(n_220),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_283),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_241),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_259),
.A2(n_248),
.B1(n_250),
.B2(n_247),
.Y(n_285)
);

INVx5_ASAP7_75t_SL g286 ( 
.A(n_253),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_288),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_262),
.B(n_218),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_246),
.B1(n_243),
.B2(n_254),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_265),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_231),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_256),
.B(n_247),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_217),
.B(n_221),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_293),
.B(n_285),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_299),
.A2(n_306),
.B(n_323),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_316),
.B1(n_295),
.B2(n_276),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_252),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_281),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_252),
.C(n_266),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_287),
.C(n_283),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_314),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_272),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_266),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_275),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_284),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_315),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_278),
.A2(n_258),
.B1(n_228),
.B2(n_261),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_318),
.A2(n_321),
.B1(n_286),
.B2(n_315),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_232),
.Y(n_320)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_279),
.A2(n_253),
.B1(n_230),
.B2(n_201),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_322),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_230),
.B(n_215),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_328),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_327),
.A2(n_329),
.B1(n_341),
.B2(n_321),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_295),
.B1(n_283),
.B2(n_273),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_288),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_334),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_299),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_301),
.A2(n_280),
.B(n_291),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_319),
.B1(n_318),
.B2(n_303),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_207),
.C(n_215),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_305),
.C(n_333),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_310),
.B(n_214),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_343),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_230),
.B1(n_201),
.B2(n_193),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_SL g343 ( 
.A(n_311),
.B(n_138),
.C(n_214),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_301),
.A2(n_186),
.B(n_181),
.Y(n_345)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_309),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_325),
.A2(n_297),
.B1(n_304),
.B2(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_327),
.A2(n_304),
.B1(n_317),
.B2(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_359),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_324),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_363),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_337),
.A2(n_308),
.B1(n_306),
.B2(n_298),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_357),
.A2(n_369),
.B1(n_330),
.B2(n_303),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_364),
.C(n_312),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_331),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_362),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_314),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_138),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_326),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_332),
.B(n_324),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_322),
.C(n_320),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_323),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_339),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_385),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_370),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_377),
.Y(n_400)
);

A2O1A1O1Ixp25_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_347),
.B(n_365),
.C(n_368),
.D(n_359),
.Y(n_375)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_375),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_388),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_347),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_302),
.C(n_348),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_386),
.C(n_390),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_319),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_382),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_339),
.C(n_336),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_354),
.B(n_196),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_389),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_196),
.C(n_169),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_369),
.A2(n_43),
.B1(n_44),
.B2(n_148),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_143),
.B1(n_114),
.B2(n_108),
.Y(n_397)
);

NOR3xp33_ASAP7_75t_SL g389 ( 
.A(n_353),
.B(n_138),
.C(n_9),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_178),
.C(n_173),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_367),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_395),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_391),
.A2(n_366),
.B(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_355),
.C(n_165),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_397),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_355),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_398),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_103),
.B(n_143),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_389),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_390),
.A2(n_114),
.B(n_12),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_402),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_373),
.C(n_379),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_410),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_373),
.Y(n_409)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_379),
.C(n_386),
.Y(n_410)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_375),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_417),
.B(n_419),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_SL g415 ( 
.A(n_392),
.B(n_103),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_415),
.A2(n_394),
.B(n_395),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_71),
.C(n_56),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_99),
.C(n_146),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_413),
.B(n_405),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_421),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_422),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_414),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_424),
.A2(n_425),
.B1(n_1),
.B2(n_3),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_414),
.B1(n_408),
.B2(n_418),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_413),
.A2(n_398),
.B(n_146),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_426),
.A2(n_430),
.B(n_4),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_413),
.A2(n_146),
.B(n_54),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_4),
.Y(n_436)
);

AOI221xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_433),
.A2(n_440),
.B(n_4),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_436),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_34),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_41),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_438),
.B(n_439),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_427),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_34),
.C(n_41),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_5),
.C(n_6),
.Y(n_449)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_423),
.B(n_6),
.Y(n_442)
);

AOI31xp67_ASAP7_75t_SL g448 ( 
.A1(n_442),
.A2(n_444),
.A3(n_5),
.B(n_6),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_5),
.Y(n_444)
);

AOI322xp5_ASAP7_75t_L g450 ( 
.A1(n_446),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_34),
.C1(n_41),
.C2(n_445),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_443),
.A2(n_433),
.B(n_437),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_447),
.A2(n_448),
.B(n_449),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_450),
.A2(n_7),
.B(n_8),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_452),
.B(n_7),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_451),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_454),
.B(n_8),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_455),
.A2(n_8),
.B(n_34),
.Y(n_456)
);


endmodule