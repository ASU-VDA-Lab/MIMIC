module real_jpeg_3804_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g129 ( 
.A(n_0),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_1),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_1),
.Y(n_243)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_2),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_3),
.A2(n_82),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_3),
.A2(n_82),
.B1(n_186),
.B2(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_3),
.A2(n_82),
.B1(n_303),
.B2(n_336),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_4),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_4),
.A2(n_177),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_4),
.A2(n_177),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_6),
.Y(n_194)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_6),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_6),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_6),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_7),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_7),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_10),
.A2(n_45),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_10),
.B(n_293),
.C(n_295),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_10),
.B(n_126),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_10),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_10),
.B(n_179),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_10),
.B(n_222),
.Y(n_370)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_12),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_12),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_12),
.A2(n_80),
.B1(n_105),
.B2(n_137),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_12),
.A2(n_137),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_12),
.A2(n_137),
.B1(n_289),
.B2(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_14),
.A2(n_63),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_14),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_14),
.A2(n_73),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_15),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_15),
.A2(n_68),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_16),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_16),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_16),
.A2(n_101),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_16),
.A2(n_101),
.B1(n_161),
.B2(n_183),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_16),
.A2(n_101),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_249),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_248),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_212),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_21),
.B(n_212),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_145),
.C(n_195),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_22),
.B(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_23),
.B(n_77),
.C(n_114),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_24),
.A2(n_50),
.B1(n_51),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_24),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.A3(n_34),
.B1(n_37),
.B2(n_44),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_27),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_28),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_28),
.Y(n_223)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_29),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_29),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_29),
.Y(n_211)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_43),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g201 ( 
.A1(n_44),
.A2(n_45),
.B(n_102),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_45),
.B(n_86),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_45),
.A2(n_52),
.B(n_306),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_SL g365 ( 
.A1(n_45),
.A2(n_366),
.B(n_369),
.Y(n_365)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_69),
.B2(n_71),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_52),
.A2(n_189),
.B1(n_237),
.B2(n_242),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_52),
.A2(n_299),
.B(n_306),
.Y(n_298)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_53),
.A2(n_72),
.B1(n_188),
.B2(n_193),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_53),
.A2(n_62),
.B1(n_238),
.B2(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_53),
.B(n_309),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_53),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_58),
.Y(n_266)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_59),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_59),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_63),
.Y(n_244)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g312 ( 
.A(n_64),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_65),
.Y(n_265)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_66),
.Y(n_245)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_67),
.Y(n_296)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_74),
.Y(n_301)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_113),
.B2(n_114),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_86),
.B(n_99),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_79),
.A2(n_86),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_87),
.B(n_100),
.Y(n_203)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_94),
.B2(n_97),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_107),
.Y(n_99)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_107),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_107),
.Y(n_226)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_134),
.B(n_139),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g218 ( 
.A1(n_115),
.A2(n_126),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_115),
.B(n_219),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_115),
.A2(n_139),
.B(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_116),
.A2(n_135),
.B1(n_144),
.B2(n_205),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_122),
.Y(n_382)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_122),
.Y(n_389)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

AO22x2_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_126)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_129),
.Y(n_291)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_129),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_129),
.Y(n_362)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g376 ( 
.A1(n_138),
.A2(n_370),
.A3(n_377),
.B1(n_379),
.B2(n_383),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_144),
.A2(n_205),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_145),
.A2(n_146),
.B1(n_195),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_187),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_147),
.B(n_187),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_172),
.B1(n_178),
.B2(n_180),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_148),
.A2(n_278),
.B(n_285),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_148),
.A2(n_178),
.B1(n_316),
.B2(n_361),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_148),
.A2(n_285),
.B(n_361),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_149),
.A2(n_179),
.B1(n_181),
.B2(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_154),
.B1(n_157),
.B2(n_161),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_165),
.B1(n_167),
.B2(n_169),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_164),
.A2(n_197),
.B(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_171),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_178),
.B(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_179),
.B(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_204),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_196),
.B(n_204),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_199),
.A2(n_200),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_208),
.Y(n_368)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_230),
.B1(n_246),
.B2(n_247),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_241),
.Y(n_331)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_271),
.B(n_408),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_268),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_252),
.B(n_268),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_259),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_253),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_259),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.C(n_267),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_260),
.B(n_399),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_262),
.B(n_267),
.Y(n_399)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_263),
.Y(n_373)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_402),
.B(n_407),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_391),
.B(n_401),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_355),
.B(n_390),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_322),
.B(n_354),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_297),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_276),
.B(n_297),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_277),
.A2(n_286),
.B1(n_287),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_284),
.Y(n_386)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_313),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_298),
.B(n_314),
.C(n_321),
.Y(n_356)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_320),
.B2(n_321),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_345),
.B(n_353),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_333),
.B(n_344),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_343),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_343),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_339),
.B(n_342),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_342),
.A2(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_351),
.Y(n_353)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_357),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_371),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_363),
.B2(n_364),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_363),
.C(n_371),
.Y(n_392)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_376),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_376),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_392),
.B(n_393),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_398),
.B2(n_400),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_397),
.C(n_400),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_398),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_403),
.B(n_404),
.Y(n_407)
);


endmodule