module fake_netlist_1_12416_n_684 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_684);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_684;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g95 ( .A(n_65), .Y(n_95) );
BUFx2_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_48), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_63), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_62), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_56), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_15), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_61), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_18), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_60), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_86), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_82), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_88), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_42), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_17), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_68), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_5), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_87), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_53), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_49), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_83), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_6), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_47), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_9), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_12), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_6), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_8), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_37), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_39), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_57), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_17), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_23), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_44), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_22), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_93), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_8), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_136), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx2_ASAP7_75t_SL g143 ( .A(n_122), .Y(n_143) );
INVx5_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_96), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_98), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_103), .B(n_19), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_100), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_114), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_122), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_131), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_100), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_103), .B(n_0), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g158 ( .A(n_146), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_157), .B(n_99), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_154), .B(n_102), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_150), .B(n_118), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_139), .B(n_106), .Y(n_164) );
BUFx10_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_142), .B(n_101), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_142), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
CKINVDCx6p67_ASAP7_75t_R g170 ( .A(n_150), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_141), .B(n_95), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_142), .B(n_101), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_157), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_143), .B(n_110), .Y(n_177) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_140), .B(n_120), .Y(n_178) );
OR2x6_ASAP7_75t_L g179 ( .A(n_143), .B(n_108), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
NOR3xp33_ASAP7_75t_L g182 ( .A(n_152), .B(n_123), .C(n_124), .Y(n_182) );
INVxp33_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_173), .B(n_99), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_166), .B(n_153), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_173), .B(n_104), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_174), .B(n_152), .Y(n_187) );
NOR2x1p5_ASAP7_75t_L g188 ( .A(n_158), .B(n_124), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_180), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_178), .B(n_150), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_178), .B(n_150), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_178), .B(n_147), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_175), .B(n_148), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_168), .B(n_104), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_176), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_175), .A2(n_156), .B1(n_155), .B2(n_151), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_168), .B(n_105), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_160), .B(n_105), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_179), .A2(n_130), .B1(n_176), .B2(n_171), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_164), .B(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_179), .B(n_112), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_173), .B(n_112), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_179), .B(n_115), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_180), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g208 ( .A(n_182), .B(n_125), .C(n_109), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_179), .B(n_115), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_173), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_156), .B(n_155), .C(n_151), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_165), .B(n_117), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_170), .B(n_125), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_177), .B(n_117), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_202), .B(n_187), .Y(n_215) );
AO22x1_ASAP7_75t_L g216 ( .A1(n_201), .A2(n_196), .B1(n_213), .B2(n_208), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_190), .A2(n_167), .B(n_163), .Y(n_217) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_213), .B(n_177), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_201), .A2(n_177), .B1(n_165), .B2(n_170), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_197), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
O2A1O1Ixp5_ASAP7_75t_L g222 ( .A1(n_184), .A2(n_120), .B(n_137), .C(n_148), .Y(n_222) );
OAI21xp33_ASAP7_75t_L g223 ( .A1(n_192), .A2(n_149), .B(n_111), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_183), .B(n_165), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_188), .B(n_119), .Y(n_225) );
OAI22x1_ASAP7_75t_L g226 ( .A1(n_187), .A2(n_134), .B1(n_128), .B2(n_116), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_192), .A2(n_149), .B(n_113), .C(n_126), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_212), .B(n_165), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_203), .A2(n_167), .B1(n_134), .B2(n_128), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_214), .B(n_167), .Y(n_230) );
AND2x2_ASAP7_75t_SL g231 ( .A(n_206), .B(n_127), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_210), .B(n_167), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_209), .B(n_167), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_185), .B(n_167), .Y(n_234) );
INVx5_ASAP7_75t_L g235 ( .A(n_210), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_210), .B(n_129), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_190), .B(n_132), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_200), .B(n_107), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_197), .B(n_133), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g240 ( .A1(n_198), .A2(n_135), .B1(n_138), .B2(n_137), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_191), .A2(n_159), .B(n_169), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_191), .A2(n_159), .B(n_169), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_186), .A2(n_172), .B(n_161), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_220), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_215), .A2(n_211), .B(n_193), .C(n_207), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_235), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_227), .A2(n_193), .B(n_207), .C(n_204), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_234), .A2(n_205), .B(n_210), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_216), .B(n_195), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_219), .A2(n_204), .B(n_194), .C(n_189), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_226), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_231), .B(n_199), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_219), .B(n_189), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_189), .B(n_194), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_235), .Y(n_257) );
AO31x2_ASAP7_75t_L g258 ( .A1(n_217), .A2(n_194), .A3(n_172), .B(n_161), .Y(n_258) );
BUFx12f_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g262 ( .A1(n_233), .A2(n_172), .B(n_161), .C(n_121), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_235), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_181), .B(n_121), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_221), .B(n_0), .Y(n_265) );
AO31x2_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_145), .A3(n_121), .B(n_144), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
OAI21x1_ASAP7_75t_SL g269 ( .A1(n_244), .A2(n_242), .B(n_228), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_244), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_245), .Y(n_272) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_223), .B(n_222), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_267), .B(n_224), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_245), .A2(n_223), .B(n_237), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_260), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_251), .B(n_240), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_250), .B(n_237), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_257), .B(n_229), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_247), .A2(n_232), .B(n_238), .Y(n_280) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_247), .A2(n_237), .B(n_145), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_266), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_249), .B(n_237), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_261), .B(n_1), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_254), .A2(n_144), .B(n_181), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_254), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_263), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
INVxp33_ASAP7_75t_L g289 ( .A(n_288), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_282), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_271), .B(n_266), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_271), .B(n_266), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_272), .B(n_249), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_282), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_286), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_270), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_282), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_270), .Y(n_298) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_275), .A2(n_278), .B(n_269), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_283), .B(n_266), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_285), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_275), .A2(n_253), .B(n_248), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_272), .B(n_249), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
AOI31xp33_ASAP7_75t_L g306 ( .A1(n_277), .A2(n_252), .A3(n_265), .B(n_262), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_283), .B(n_258), .Y(n_309) );
BUFx4f_ASAP7_75t_SL g310 ( .A(n_287), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_287), .B(n_257), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_283), .B(n_258), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_283), .B(n_257), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_291), .B(n_281), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_311), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_281), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_311), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_291), .B(n_281), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_305), .B(n_274), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_292), .B(n_281), .Y(n_323) );
BUFx2_ASAP7_75t_SL g324 ( .A(n_310), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_296), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_290), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_312), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_290), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_281), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_305), .B(n_274), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_292), .B(n_280), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_294), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_304), .B(n_280), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_300), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_297), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_297), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_304), .B(n_280), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_300), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_304), .B(n_280), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_300), .B(n_283), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_296), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_300), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_296), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_316), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_316), .B(n_308), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_337), .B(n_309), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_337), .B(n_309), .Y(n_363) );
NOR2x1_ASAP7_75t_L g364 ( .A(n_324), .B(n_283), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_339), .B(n_309), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_354), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_329), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_339), .B(n_309), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_318), .B(n_313), .Y(n_369) );
NOR2x1_ASAP7_75t_L g370 ( .A(n_324), .B(n_308), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_313), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_322), .B(n_259), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_344), .B(n_313), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_332), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_354), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_345), .B(n_313), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_346), .B(n_317), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_346), .B(n_313), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_348), .B(n_299), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_317), .B(n_299), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_351), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_351), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_348), .B(n_299), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_345), .B(n_293), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_336), .B(n_289), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_319), .B(n_299), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_319), .B(n_299), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_321), .B(n_307), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_328), .B(n_289), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_353), .B(n_293), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_321), .B(n_307), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_341), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_332), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_338), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_338), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_323), .B(n_314), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_348), .B(n_314), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_342), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_323), .B(n_314), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_333), .B(n_303), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_351), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_333), .B(n_303), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_357), .B(n_312), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_342), .B(n_312), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_357), .B(n_308), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_349), .B(n_298), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_353), .B(n_308), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_355), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_341), .B(n_308), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_326), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_350), .B(n_280), .Y(n_417) );
HB1xp67_ASAP7_75t_SL g418 ( .A(n_348), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_326), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_355), .B(n_298), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_347), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_326), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_381), .B(n_350), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_366), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_359), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_381), .B(n_347), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_363), .B(n_352), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_359), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_391), .B(n_352), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_384), .A2(n_277), .B1(n_298), .B2(n_268), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_406), .B(n_356), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_363), .B(n_327), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_385), .B(n_327), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_385), .B(n_327), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_392), .B(n_331), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_392), .B(n_331), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_362), .B(n_356), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_362), .B(n_356), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_406), .B(n_325), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_361), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_369), .B(n_390), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_393), .B(n_331), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_361), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_369), .B(n_334), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_370), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_379), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_367), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_418), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_390), .B(n_334), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_379), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_408), .B(n_334), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_367), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_375), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_387), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_384), .B(n_335), .Y(n_458) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_398), .B(n_351), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_387), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_393), .B(n_335), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_365), .B(n_335), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_394), .B(n_343), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_408), .B(n_343), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_421), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_375), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_376), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_365), .B(n_343), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_377), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_378), .B(n_340), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_368), .B(n_351), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_399), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_368), .B(n_351), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_396), .B(n_340), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_401), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_373), .Y(n_478) );
AOI211xp5_ASAP7_75t_L g479 ( .A1(n_358), .A2(n_268), .B(n_284), .C(n_246), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_401), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_371), .B(n_285), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_360), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_371), .B(n_285), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_404), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_409), .B(n_306), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_374), .B(n_285), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_374), .B(n_278), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_416), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_382), .B(n_258), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_398), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_404), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_400), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_409), .B(n_306), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_382), .B(n_258), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_396), .B(n_284), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_410), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_412), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_402), .B(n_273), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_395), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_402), .B(n_276), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_403), .B(n_259), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_394), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_444), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_497), .B(n_405), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_423), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_503), .B(n_397), .Y(n_508) );
XNOR2xp5_ASAP7_75t_L g509 ( .A(n_451), .B(n_405), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_469), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_471), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_478), .B(n_403), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_482), .B(n_364), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_424), .B(n_403), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_474), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_493), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_427), .B(n_397), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_427), .B(n_380), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_441), .Y(n_519) );
NAND2x1_ASAP7_75t_L g520 ( .A(n_448), .B(n_386), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_431), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_424), .B(n_415), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_441), .B(n_380), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_426), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_465), .Y(n_525) );
NOR2x2_ASAP7_75t_L g526 ( .A(n_502), .B(n_360), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_440), .B(n_415), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_491), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_500), .B(n_417), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_436), .B(n_417), .Y(n_530) );
AND2x4_ASAP7_75t_SL g531 ( .A(n_502), .B(n_386), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_425), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_429), .B(n_384), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_430), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_442), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_432), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_434), .B(n_389), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_443), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_436), .B(n_411), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_446), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_459), .Y(n_541) );
NOR3xp33_ASAP7_75t_SL g542 ( .A(n_486), .B(n_420), .C(n_279), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_437), .B(n_411), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_429), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_450), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_437), .B(n_413), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_473), .B(n_389), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_455), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_459), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_456), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_498), .B(n_360), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_454), .B(n_389), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_468), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_438), .B(n_413), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_477), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_438), .B(n_419), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_462), .B(n_386), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_439), .B(n_419), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_479), .A2(n_422), .B1(n_388), .B2(n_407), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_473), .B(n_388), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_466), .B(n_422), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_492), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_494), .A2(n_388), .B1(n_407), .B2(n_269), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_476), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_425), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_439), .B(n_407), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_501), .B(n_1), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_433), .A2(n_264), .B(n_3), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_428), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_448), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_445), .B(n_2), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_475), .B(n_144), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_445), .B(n_2), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_461), .B(n_273), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_535), .A2(n_488), .B1(n_495), .B2(n_490), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_461), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_510), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_572), .A2(n_464), .B(n_435), .Y(n_581) );
AOI32xp33_ASAP7_75t_L g582 ( .A1(n_507), .A2(n_482), .A3(n_435), .B1(n_470), .B2(n_464), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_544), .B(n_470), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_520), .A2(n_472), .B(n_458), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_515), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_516), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_561), .B(n_549), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g588 ( .A1(n_521), .A2(n_496), .B(n_495), .C(n_490), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_575), .A2(n_496), .B(n_489), .C(n_485), .Y(n_589) );
OAI32xp33_ASAP7_75t_L g590 ( .A1(n_528), .A2(n_447), .A3(n_452), .B1(n_487), .B2(n_481), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_565), .B(n_489), .C(n_485), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_547), .B(n_481), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_531), .A2(n_487), .B1(n_483), .B2(n_488), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_517), .B(n_566), .Y(n_594) );
AOI21xp33_ASAP7_75t_L g595 ( .A1(n_569), .A2(n_447), .B(n_452), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_504), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_505), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_561), .A2(n_483), .B1(n_458), .B2(n_499), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_509), .A2(n_458), .B(n_499), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_524), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_570), .A2(n_467), .B(n_463), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_536), .B(n_463), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_534), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_542), .B(n_467), .C(n_460), .Y(n_604) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_573), .A2(n_460), .B(n_457), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_557), .B(n_449), .C(n_453), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_512), .A2(n_449), .B1(n_273), .B2(n_256), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_540), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_551), .A2(n_273), .B1(n_262), .B2(n_181), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_513), .A2(n_273), .B1(n_5), .B2(n_7), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
AOI31xp33_ASAP7_75t_SL g613 ( .A1(n_526), .A2(n_4), .A3(n_7), .B(n_9), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_530), .B(n_10), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_548), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_525), .Y(n_616) );
OAI31xp33_ASAP7_75t_L g617 ( .A1(n_513), .A2(n_10), .A3(n_11), .B(n_12), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_541), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_550), .Y(n_619) );
OAI321xp33_ASAP7_75t_L g620 ( .A1(n_570), .A2(n_13), .A3(n_16), .B1(n_181), .B2(n_21), .C(n_24), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_553), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_541), .B(n_16), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_602), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_599), .A2(n_518), .B1(n_523), .B2(n_506), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_599), .A2(n_506), .B1(n_529), .B2(n_537), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_590), .A2(n_555), .B1(n_558), .B2(n_559), .C(n_564), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_600), .Y(n_628) );
NOR2xp67_ASAP7_75t_SL g629 ( .A(n_622), .B(n_574), .Y(n_629) );
OAI322xp33_ASAP7_75t_SL g630 ( .A1(n_587), .A2(n_539), .A3(n_543), .B1(n_546), .B2(n_554), .C1(n_519), .C2(n_556), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_593), .A2(n_552), .B1(n_527), .B2(n_514), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_588), .A2(n_556), .B(n_560), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_603), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_617), .B(n_562), .C(n_560), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_582), .A2(n_533), .B1(n_563), .B2(n_522), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_607), .Y(n_636) );
OAI21xp33_ASAP7_75t_SL g637 ( .A1(n_583), .A2(n_568), .B(n_576), .Y(n_637) );
NAND4xp25_ASAP7_75t_SL g638 ( .A(n_589), .B(n_576), .C(n_571), .D(n_567), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_609), .Y(n_639) );
AOI221x1_ASAP7_75t_L g640 ( .A1(n_618), .A2(n_532), .B1(n_25), .B2(n_26), .C(n_28), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_595), .A2(n_20), .B1(n_29), .B2(n_30), .C(n_31), .Y(n_641) );
OAI222xp33_ASAP7_75t_L g642 ( .A1(n_598), .A2(n_32), .B1(n_34), .B2(n_35), .C1(n_36), .C2(n_38), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_584), .A2(n_40), .B(n_41), .Y(n_643) );
AOI211xp5_ASAP7_75t_SL g644 ( .A1(n_613), .A2(n_43), .B(n_45), .C(n_46), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_612), .Y(n_645) );
AOI21xp5_ASAP7_75t_R g646 ( .A1(n_613), .A2(n_50), .B(n_51), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
AO22x2_ASAP7_75t_L g648 ( .A1(n_591), .A2(n_52), .B1(n_54), .B2(n_55), .Y(n_648) );
NOR4xp25_ASAP7_75t_L g649 ( .A(n_614), .B(n_58), .C(n_59), .D(n_64), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_617), .A2(n_605), .B(n_611), .C(n_581), .Y(n_650) );
NOR2xp33_ASAP7_75t_SL g651 ( .A(n_616), .B(n_66), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_620), .A2(n_67), .B(n_69), .C(n_70), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_601), .A2(n_71), .B(n_72), .C(n_73), .Y(n_653) );
AOI21xp33_ASAP7_75t_SL g654 ( .A1(n_606), .A2(n_75), .B(n_78), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_604), .A2(n_79), .B(n_80), .C(n_81), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_596), .A2(n_90), .B1(n_91), .B2(n_92), .C(n_94), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_597), .B(n_586), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_579), .A2(n_585), .B(n_580), .C(n_577), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_619), .A2(n_621), .B1(n_592), .B2(n_608), .C(n_578), .Y(n_659) );
NAND4xp25_ASAP7_75t_SL g660 ( .A(n_610), .B(n_582), .C(n_588), .D(n_451), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_624), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g662 ( .A(n_634), .B(n_660), .C(n_642), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_644), .B(n_650), .C(n_652), .D(n_643), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_630), .A2(n_625), .B1(n_638), .B2(n_659), .C(n_626), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_658), .B(n_632), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_627), .A2(n_637), .B(n_646), .C(n_641), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_653), .B(n_656), .C(n_654), .Y(n_667) );
XNOR2x1_ASAP7_75t_L g668 ( .A(n_665), .B(n_648), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_661), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_666), .B(n_657), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_662), .B(n_640), .C(n_655), .D(n_651), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_669), .B(n_671), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_670), .B(n_663), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_668), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_672), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_674), .Y(n_676) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_675), .B(n_673), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_676), .A2(n_664), .B1(n_623), .B2(n_631), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_677), .Y(n_679) );
NAND2xp33_ASAP7_75t_SL g680 ( .A(n_678), .B(n_629), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_679), .A2(n_667), .B1(n_657), .B2(n_635), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_680), .B(n_649), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_682), .A2(n_648), .B(n_645), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_628), .B1(n_647), .B2(n_633), .C1(n_636), .C2(n_639), .Y(n_684) );
endmodule