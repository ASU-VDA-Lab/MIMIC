module real_aes_7313_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_385;
wire n_214;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g240 ( .A1(n_0), .A2(n_241), .B(n_242), .C(n_246), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_1), .B(n_182), .Y(n_247) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_92), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g464 ( .A(n_2), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_3), .B(n_154), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_4), .A2(n_140), .B(n_145), .C(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_5), .A2(n_135), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_6), .A2(n_135), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_7), .B(n_182), .Y(n_556) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_8), .A2(n_170), .B(n_186), .Y(n_185) );
AND2x6_ASAP7_75t_L g140 ( .A(n_9), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_10), .A2(n_140), .B(n_145), .C(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g494 ( .A(n_11), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_12), .B(n_41), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_13), .B(n_245), .Y(n_514) );
INVx1_ASAP7_75t_L g164 ( .A(n_14), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_15), .B(n_154), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_16), .A2(n_155), .B(n_502), .C(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_17), .B(n_182), .Y(n_505) );
AOI22xp5_ASAP7_75t_SL g468 ( .A1(n_18), .A2(n_462), .B1(n_469), .B2(n_751), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_19), .A2(n_47), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_19), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_19), .B(n_219), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_20), .A2(n_145), .B(n_196), .C(n_215), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_21), .A2(n_194), .B(n_244), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_22), .B(n_245), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_23), .B(n_245), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_24), .Y(n_541) );
INVx1_ASAP7_75t_L g533 ( .A(n_25), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_26), .A2(n_145), .B(n_189), .C(n_196), .Y(n_188) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_28), .Y(n_510) );
INVx1_ASAP7_75t_L g590 ( .A(n_29), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_30), .A2(n_135), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g138 ( .A(n_31), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_32), .A2(n_143), .B(n_158), .C(n_204), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_33), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_34), .A2(n_244), .B(n_553), .C(n_555), .Y(n_552) );
INVxp67_ASAP7_75t_L g591 ( .A(n_35), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_36), .A2(n_46), .B1(n_126), .B2(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_36), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_37), .B(n_191), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_38), .A2(n_145), .B(n_196), .C(n_532), .Y(n_531) );
CKINVDCx14_ASAP7_75t_R g551 ( .A(n_39), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_40), .A2(n_45), .B1(n_476), .B2(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_40), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_42), .A2(n_246), .B(n_492), .C(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_43), .B(n_213), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_44), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_45), .Y(n_476) );
INVx1_ASAP7_75t_L g127 ( .A(n_46), .Y(n_127) );
INVx1_ASAP7_75t_L g123 ( .A(n_47), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_48), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_49), .B(n_135), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_50), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_51), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_52), .A2(n_143), .B(n_148), .C(n_158), .Y(n_142) );
INVx1_ASAP7_75t_L g243 ( .A(n_53), .Y(n_243) );
INVx1_ASAP7_75t_L g149 ( .A(n_54), .Y(n_149) );
INVx1_ASAP7_75t_L g522 ( .A(n_55), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_56), .B(n_135), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_57), .Y(n_222) );
CKINVDCx14_ASAP7_75t_R g490 ( .A(n_58), .Y(n_490) );
INVx1_ASAP7_75t_L g141 ( .A(n_59), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_60), .B(n_135), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_61), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_62), .A2(n_176), .B(n_178), .C(n_180), .Y(n_175) );
INVx1_ASAP7_75t_L g163 ( .A(n_63), .Y(n_163) );
INVx1_ASAP7_75t_SL g554 ( .A(n_64), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_66), .B(n_154), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_67), .B(n_182), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_68), .B(n_155), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_69), .A2(n_105), .B1(n_113), .B2(n_756), .Y(n_104) );
INVx1_ASAP7_75t_L g544 ( .A(n_70), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_71), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_72), .B(n_151), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_73), .A2(n_145), .B(n_158), .C(n_228), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_74), .Y(n_174) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_76), .A2(n_135), .B(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_77), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_78), .A2(n_135), .B(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_79), .A2(n_471), .B1(n_472), .B2(n_478), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_79), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_80), .A2(n_213), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g500 ( .A(n_81), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_82), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_83), .B(n_150), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_84), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_84), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_85), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_86), .A2(n_135), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g503 ( .A(n_87), .Y(n_503) );
INVx2_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
INVx1_ASAP7_75t_L g513 ( .A(n_89), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_90), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_91), .B(n_245), .Y(n_258) );
OR2x2_ASAP7_75t_L g461 ( .A(n_92), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g481 ( .A(n_92), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_93), .A2(n_145), .B(n_158), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_94), .B(n_135), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_95), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g205 ( .A(n_96), .Y(n_205) );
INVxp67_ASAP7_75t_L g179 ( .A(n_97), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_98), .B(n_170), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g229 ( .A(n_100), .Y(n_229) );
INVx1_ASAP7_75t_L g253 ( .A(n_101), .Y(n_253) );
INVx2_ASAP7_75t_L g525 ( .A(n_102), .Y(n_525) );
AND2x2_ASAP7_75t_L g165 ( .A(n_103), .B(n_160), .Y(n_165) );
INVx1_ASAP7_75t_SL g756 ( .A(n_105), .Y(n_756) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g463 ( .A(n_107), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_467), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g755 ( .A(n_117), .Y(n_755) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_458), .B(n_465), .Y(n_119) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
XOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_128), .A2(n_480), .B1(n_482), .B2(n_749), .Y(n_479) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR5x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_331), .C(n_409), .D(n_433), .E(n_450), .Y(n_129) );
OAI211xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_197), .B(n_248), .C(n_308), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_166), .Y(n_131) );
AND2x2_ASAP7_75t_L g262 ( .A(n_132), .B(n_168), .Y(n_262) );
INVx5_ASAP7_75t_SL g290 ( .A(n_132), .Y(n_290) );
AND2x2_ASAP7_75t_L g326 ( .A(n_132), .B(n_311), .Y(n_326) );
OR2x2_ASAP7_75t_L g365 ( .A(n_132), .B(n_167), .Y(n_365) );
OR2x2_ASAP7_75t_L g396 ( .A(n_132), .B(n_287), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_132), .B(n_300), .Y(n_432) );
AND2x2_ASAP7_75t_L g444 ( .A(n_132), .B(n_287), .Y(n_444) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_165), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_142), .B(n_160), .Y(n_133) );
BUFx2_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g254 ( .A(n_136), .B(n_140), .Y(n_254) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
INVx1_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_139), .Y(n_245) );
INVx4_ASAP7_75t_SL g159 ( .A(n_140), .Y(n_159) );
BUFx3_ASAP7_75t_L g196 ( .A(n_140), .Y(n_196) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_144), .A2(n_159), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_144), .A2(n_159), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_144), .A2(n_159), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_144), .A2(n_159), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_144), .A2(n_159), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_144), .A2(n_159), .B(n_551), .C(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_SL g586 ( .A1(n_144), .A2(n_159), .B(n_587), .C(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_153), .C(n_156), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_150), .A2(n_156), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_L g512 ( .A1(n_150), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_150), .A2(n_515), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_154), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g241 ( .A(n_154), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_154), .A2(n_218), .B(n_533), .C(n_534), .Y(n_532) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_154), .A2(n_177), .B1(n_590), .B2(n_591), .Y(n_589) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_155), .B(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g246 ( .A(n_157), .Y(n_246) );
INVx1_ASAP7_75t_L g504 ( .A(n_157), .Y(n_504) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_160), .A2(n_202), .B(n_203), .Y(n_201) );
INVx2_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_160), .Y(n_223) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_160), .A2(n_488), .B(n_495), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_160), .A2(n_254), .B(n_530), .C(n_531), .Y(n_529) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g171 ( .A(n_161), .B(n_162), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
AND2x2_ASAP7_75t_L g443 ( .A(n_166), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g306 ( .A(n_167), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_168), .B(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_168), .Y(n_299) );
INVx3_ASAP7_75t_L g314 ( .A(n_168), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_168), .B(n_184), .Y(n_338) );
OR2x2_ASAP7_75t_L g347 ( .A(n_168), .B(n_290), .Y(n_347) );
AND2x2_ASAP7_75t_L g351 ( .A(n_168), .B(n_311), .Y(n_351) );
AND2x2_ASAP7_75t_L g357 ( .A(n_168), .B(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g394 ( .A(n_168), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_168), .B(n_251), .Y(n_408) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_181), .Y(n_168) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_169), .A2(n_498), .B(n_505), .Y(n_497) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_169), .A2(n_520), .B(n_526), .Y(n_519) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_169), .A2(n_549), .B(n_556), .Y(n_548) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g183 ( .A(n_170), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_170), .A2(n_187), .B(n_188), .Y(n_186) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g261 ( .A(n_171), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_176), .A2(n_229), .B(n_230), .C(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_177), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_177), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g218 ( .A(n_180), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_180), .B(n_589), .Y(n_588) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_182), .A2(n_237), .B(n_247), .Y(n_236) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_183), .B(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_183), .A2(n_226), .B(n_234), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_183), .B(n_235), .Y(n_234) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_183), .A2(n_252), .B(n_259), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_183), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_183), .B(n_536), .Y(n_535) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_183), .A2(n_540), .B(n_546), .Y(n_539) );
OR2x2_ASAP7_75t_L g300 ( .A(n_184), .B(n_251), .Y(n_300) );
AND2x2_ASAP7_75t_L g311 ( .A(n_184), .B(n_287), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_184), .B(n_314), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_184), .B(n_251), .Y(n_346) );
INVx1_ASAP7_75t_SL g358 ( .A(n_184), .Y(n_358) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g250 ( .A(n_185), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_185), .B(n_290), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B(n_193), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_193), .A2(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_209), .Y(n_198) );
AND2x2_ASAP7_75t_L g271 ( .A(n_199), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_199), .B(n_224), .Y(n_275) );
AND2x2_ASAP7_75t_L g278 ( .A(n_199), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_199), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g303 ( .A(n_199), .B(n_294), .Y(n_303) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_199), .Y(n_322) );
AND2x2_ASAP7_75t_L g343 ( .A(n_199), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g353 ( .A(n_199), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g399 ( .A(n_199), .B(n_282), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_199), .B(n_305), .Y(n_426) );
INVx5_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g296 ( .A(n_200), .Y(n_296) );
AND2x2_ASAP7_75t_L g362 ( .A(n_200), .B(n_294), .Y(n_362) );
AND2x2_ASAP7_75t_L g446 ( .A(n_200), .B(n_314), .Y(n_446) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_207), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_209), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_209), .Y(n_435) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_224), .Y(n_209) );
AND2x2_ASAP7_75t_L g265 ( .A(n_210), .B(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g274 ( .A(n_210), .B(n_272), .Y(n_274) );
INVx5_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
AND2x2_ASAP7_75t_L g305 ( .A(n_210), .B(n_236), .Y(n_305) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_210), .Y(n_342) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
AOI21xp5_ASAP7_75t_SL g211 ( .A1(n_212), .A2(n_214), .B(n_219), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_220), .B(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_223), .A2(n_509), .B(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g383 ( .A(n_224), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_224), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g416 ( .A(n_224), .B(n_282), .Y(n_416) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_224), .A2(n_339), .B(n_446), .C(n_447), .Y(n_445) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_236), .Y(n_224) );
BUFx2_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
INVx2_ASAP7_75t_L g270 ( .A(n_225), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g555 ( .A(n_232), .Y(n_555) );
INVx2_ASAP7_75t_L g272 ( .A(n_236), .Y(n_272) );
AND2x2_ASAP7_75t_L g279 ( .A(n_236), .B(n_270), .Y(n_279) );
AND2x2_ASAP7_75t_L g370 ( .A(n_236), .B(n_282), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_244), .B(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g492 ( .A(n_245), .Y(n_492) );
INVx2_ASAP7_75t_L g515 ( .A(n_246), .Y(n_515) );
AOI211x1_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_263), .B(n_276), .C(n_301), .Y(n_248) );
INVx1_ASAP7_75t_L g367 ( .A(n_249), .Y(n_367) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_262), .Y(n_249) );
INVx5_ASAP7_75t_SL g287 ( .A(n_251), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_251), .B(n_357), .Y(n_356) );
AOI311xp33_ASAP7_75t_L g375 ( .A1(n_251), .A2(n_376), .A3(n_378), .B(n_379), .C(n_385), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_251), .A2(n_323), .B(n_411), .C(n_414), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_255), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_254), .A2(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_254), .A2(n_541), .B(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g583 ( .A(n_261), .Y(n_583) );
INVxp67_ASAP7_75t_L g330 ( .A(n_262), .Y(n_330) );
NAND4xp25_ASAP7_75t_SL g263 ( .A(n_264), .B(n_267), .C(n_273), .D(n_275), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_264), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g321 ( .A(n_265), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_268), .B(n_274), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_268), .B(n_281), .Y(n_401) );
BUFx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_269), .B(n_282), .Y(n_419) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g294 ( .A(n_270), .Y(n_294) );
INVxp67_ASAP7_75t_L g329 ( .A(n_271), .Y(n_329) );
AND2x4_ASAP7_75t_L g281 ( .A(n_272), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g355 ( .A(n_272), .B(n_294), .Y(n_355) );
INVx1_ASAP7_75t_L g382 ( .A(n_272), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_272), .B(n_369), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_273), .B(n_343), .Y(n_363) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_274), .B(n_296), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_274), .B(n_343), .Y(n_442) );
INVx1_ASAP7_75t_L g453 ( .A(n_275), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_283), .C(n_291), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g333 ( .A(n_279), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g315 ( .A(n_280), .Y(n_315) );
AND2x2_ASAP7_75t_L g292 ( .A(n_281), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_281), .B(n_343), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_281), .B(n_362), .Y(n_386) );
OR2x2_ASAP7_75t_L g302 ( .A(n_282), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g334 ( .A(n_282), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_282), .B(n_294), .Y(n_349) );
AND2x2_ASAP7_75t_L g406 ( .A(n_282), .B(n_362), .Y(n_406) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_282), .Y(n_413) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_284), .A2(n_296), .B1(n_418), .B2(n_420), .C(n_423), .Y(n_417) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_290), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_287), .B(n_357), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_287), .B(n_314), .Y(n_422) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g407 ( .A(n_289), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g421 ( .A(n_289), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_290), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g318 ( .A(n_290), .B(n_311), .Y(n_318) );
AND2x2_ASAP7_75t_L g388 ( .A(n_290), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_290), .B(n_337), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_290), .B(n_438), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_295), .B(n_297), .Y(n_291) );
INVx2_ASAP7_75t_L g324 ( .A(n_292), .Y(n_324) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g344 ( .A(n_294), .Y(n_344) );
OR2x2_ASAP7_75t_L g348 ( .A(n_296), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g451 ( .A(n_296), .B(n_419), .Y(n_451) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AOI21xp33_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_304), .B(n_306), .Y(n_301) );
INVx1_ASAP7_75t_L g455 ( .A(n_302), .Y(n_455) );
INVx2_ASAP7_75t_SL g369 ( .A(n_303), .Y(n_369) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_306), .A2(n_387), .B(n_451), .C(n_452), .Y(n_450) );
OAI322xp33_ASAP7_75t_SL g319 ( .A1(n_307), .A2(n_320), .A3(n_323), .B1(n_324), .B2(n_325), .C1(n_327), .C2(n_330), .Y(n_319) );
INVx2_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_315), .B1(n_316), .B2(n_318), .C(n_319), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI22xp33_ASAP7_75t_SL g385 ( .A1(n_310), .A2(n_386), .B1(n_387), .B2(n_390), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_311), .B(n_314), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_311), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g384 ( .A(n_313), .B(n_346), .Y(n_384) );
INVx1_ASAP7_75t_L g374 ( .A(n_314), .Y(n_374) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_318), .A2(n_428), .B(n_430), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g352 ( .A1(n_320), .A2(n_353), .B(n_356), .Y(n_352) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp67_ASAP7_75t_SL g381 ( .A(n_322), .B(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_322), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g438 ( .A(n_323), .Y(n_438) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND4xp25_ASAP7_75t_L g331 ( .A(n_332), .B(n_359), .C(n_375), .D(n_391), .Y(n_331) );
AOI211xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_340), .C(n_352), .Y(n_332) );
INVx1_ASAP7_75t_L g424 ( .A(n_333), .Y(n_424) );
AND2x2_ASAP7_75t_L g372 ( .A(n_334), .B(n_355), .Y(n_372) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_339), .B(n_374), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B1(n_348), .B2(n_350), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_342), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g404 ( .A1(n_343), .A2(n_382), .B(n_405), .C(n_407), .Y(n_404) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g389 ( .A(n_346), .Y(n_389) );
INVx1_ASAP7_75t_L g449 ( .A(n_347), .Y(n_449) );
NAND2xp33_ASAP7_75t_SL g439 ( .A(n_348), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g378 ( .A(n_357), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B(n_364), .C(n_366), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_371), .B2(n_373), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_369), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_374), .B(n_395), .Y(n_457) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_383), .B(n_384), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_397), .B1(n_400), .B2(n_402), .C(n_404), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_407), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
NAND3xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_417), .C(n_427), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_436), .C(n_445), .Y(n_433) );
INVx1_ASAP7_75t_L g454 ( .A(n_434), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_441), .B2(n_443), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g466 ( .A(n_461), .Y(n_466) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_462), .B(n_481), .Y(n_753) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_465), .B(n_468), .C(n_754), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g750 ( .A(n_481), .Y(n_750) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_679), .Y(n_482) );
NAND5xp2_ASAP7_75t_L g483 ( .A(n_484), .B(n_594), .C(n_626), .D(n_643), .E(n_666), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_527), .B1(n_557), .B2(n_561), .C(n_565), .Y(n_484) );
INVx1_ASAP7_75t_L g706 ( .A(n_485), .Y(n_706) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_506), .Y(n_485) );
AND3x2_ASAP7_75t_L g681 ( .A(n_486), .B(n_508), .C(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_487), .B(n_563), .Y(n_562) );
BUFx3_ASAP7_75t_L g572 ( .A(n_487), .Y(n_572) );
AND2x2_ASAP7_75t_L g576 ( .A(n_487), .B(n_518), .Y(n_576) );
INVx2_ASAP7_75t_L g603 ( .A(n_487), .Y(n_603) );
OR2x2_ASAP7_75t_L g614 ( .A(n_487), .B(n_519), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_487), .B(n_507), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_487), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g693 ( .A(n_487), .B(n_519), .Y(n_693) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_496), .Y(n_575) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_496), .B(n_507), .Y(n_653) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g564 ( .A(n_497), .B(n_507), .Y(n_564) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
AND2x2_ASAP7_75t_L g620 ( .A(n_497), .B(n_519), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_497), .B(n_506), .C(n_603), .Y(n_645) );
AND2x2_ASAP7_75t_L g710 ( .A(n_497), .B(n_508), .Y(n_710) );
AND2x2_ASAP7_75t_L g744 ( .A(n_497), .B(n_507), .Y(n_744) );
INVxp67_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_507), .B(n_603), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_507), .B(n_634), .Y(n_642) );
AND2x2_ASAP7_75t_L g692 ( .A(n_507), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g720 ( .A(n_507), .Y(n_720) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g627 ( .A(n_508), .B(n_620), .Y(n_627) );
BUFx3_ASAP7_75t_L g659 ( .A(n_508), .Y(n_659) );
INVx2_ASAP7_75t_L g635 ( .A(n_518), .Y(n_635) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_527), .A2(n_695), .B1(n_697), .B2(n_698), .Y(n_694) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_537), .Y(n_527) );
AND2x2_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
INVx3_ASAP7_75t_SL g568 ( .A(n_528), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_528), .B(n_598), .Y(n_630) );
OR2x2_ASAP7_75t_L g649 ( .A(n_528), .B(n_538), .Y(n_649) );
AND2x2_ASAP7_75t_L g654 ( .A(n_528), .B(n_606), .Y(n_654) );
AND2x2_ASAP7_75t_L g657 ( .A(n_528), .B(n_599), .Y(n_657) );
AND2x2_ASAP7_75t_L g669 ( .A(n_528), .B(n_548), .Y(n_669) );
AND2x2_ASAP7_75t_L g685 ( .A(n_528), .B(n_539), .Y(n_685) );
AND2x4_ASAP7_75t_L g688 ( .A(n_528), .B(n_559), .Y(n_688) );
OR2x2_ASAP7_75t_L g705 ( .A(n_528), .B(n_641), .Y(n_705) );
OR2x2_ASAP7_75t_L g736 ( .A(n_528), .B(n_581), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_528), .B(n_664), .Y(n_738) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_535), .Y(n_528) );
AND2x2_ASAP7_75t_L g612 ( .A(n_537), .B(n_579), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_537), .B(n_599), .Y(n_731) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_548), .Y(n_537) );
AND2x2_ASAP7_75t_L g567 ( .A(n_538), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g598 ( .A(n_538), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g606 ( .A(n_538), .B(n_581), .Y(n_606) );
AND2x2_ASAP7_75t_L g624 ( .A(n_538), .B(n_559), .Y(n_624) );
OR2x2_ASAP7_75t_L g641 ( .A(n_538), .B(n_599), .Y(n_641) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g560 ( .A(n_539), .Y(n_560) );
AND2x2_ASAP7_75t_L g664 ( .A(n_539), .B(n_548), .Y(n_664) );
INVx2_ASAP7_75t_L g559 ( .A(n_548), .Y(n_559) );
INVx1_ASAP7_75t_L g676 ( .A(n_548), .Y(n_676) );
AND2x2_ASAP7_75t_L g726 ( .A(n_548), .B(n_568), .Y(n_726) );
AND2x2_ASAP7_75t_L g578 ( .A(n_558), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g610 ( .A(n_558), .B(n_568), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_558), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g597 ( .A(n_559), .B(n_568), .Y(n_597) );
OR2x2_ASAP7_75t_L g713 ( .A(n_560), .B(n_687), .Y(n_713) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_563), .B(n_693), .Y(n_699) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
OAI32xp33_ASAP7_75t_L g655 ( .A1(n_564), .A2(n_656), .A3(n_658), .B1(n_660), .B2(n_661), .Y(n_655) );
OR2x2_ASAP7_75t_L g672 ( .A(n_564), .B(n_614), .Y(n_672) );
OAI21xp33_ASAP7_75t_SL g697 ( .A1(n_564), .A2(n_574), .B(n_602), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_574), .B2(n_577), .Y(n_565) );
INVxp33_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_567), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_568), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g623 ( .A(n_568), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g723 ( .A(n_568), .B(n_664), .Y(n_723) );
OR2x2_ASAP7_75t_L g747 ( .A(n_568), .B(n_641), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g730 ( .A1(n_569), .A2(n_629), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g607 ( .A(n_571), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_571), .B(n_576), .Y(n_625) );
AND2x2_ASAP7_75t_L g647 ( .A(n_572), .B(n_620), .Y(n_647) );
INVx1_ASAP7_75t_L g660 ( .A(n_572), .Y(n_660) );
OR2x2_ASAP7_75t_L g665 ( .A(n_572), .B(n_599), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_575), .B(n_614), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_576), .A2(n_596), .B1(n_601), .B2(n_605), .Y(n_595) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_579), .A2(n_638), .B1(n_645), .B2(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g722 ( .A(n_579), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_581), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g741 ( .A(n_581), .B(n_624), .Y(n_741) );
AO21x2_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B(n_592), .Y(n_581) );
INVx1_ASAP7_75t_L g600 ( .A(n_582), .Y(n_600) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OA21x2_ASAP7_75t_L g599 ( .A1(n_585), .A2(n_593), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_607), .B1(n_608), .B2(n_613), .C(n_615), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_597), .B(n_599), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_597), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g616 ( .A(n_598), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g703 ( .A1(n_598), .A2(n_704), .B(n_705), .C(n_706), .Y(n_703) );
AND2x2_ASAP7_75t_L g708 ( .A(n_598), .B(n_688), .Y(n_708) );
O2A1O1Ixp33_ASAP7_75t_SL g746 ( .A1(n_598), .A2(n_687), .B(n_747), .C(n_748), .Y(n_746) );
BUFx3_ASAP7_75t_L g638 ( .A(n_599), .Y(n_638) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_602), .B(n_659), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g721 ( .A1(n_602), .A2(n_722), .B(n_724), .C(n_730), .Y(n_721) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVxp67_ASAP7_75t_L g682 ( .A(n_604), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_606), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_610), .A2(n_627), .B(n_628), .C(n_636), .Y(n_626) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g711 ( .A(n_614), .Y(n_711) );
OR2x2_ASAP7_75t_L g728 ( .A(n_614), .B(n_658), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_622), .B2(n_625), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_617), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
OR2x2_ASAP7_75t_L g715 ( .A(n_619), .B(n_659), .Y(n_715) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g670 ( .A(n_620), .B(n_660), .Y(n_670) );
INVx1_ASAP7_75t_L g678 ( .A(n_621), .Y(n_678) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_624), .B(n_638), .Y(n_686) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_634), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g743 ( .A(n_635), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_642), .Y(n_636) );
INVx1_ASAP7_75t_L g673 ( .A(n_637), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_638), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_638), .B(n_669), .Y(n_668) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_638), .B(n_664), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_638), .B(n_685), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_638), .A2(n_648), .B(n_688), .C(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AOI221xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_648), .B1(n_650), .B2(n_654), .C(n_655), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_652), .B(n_660), .Y(n_734) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_654), .A2(n_669), .B(n_671), .C(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_657), .B(n_664), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_658), .B(n_711), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
INVxp33_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AOI21xp33_ASAP7_75t_SL g674 ( .A1(n_663), .A2(n_675), .B(n_677), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_663), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_664), .B(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B1(n_671), .B2(n_673), .C(n_674), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_670), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g704 ( .A(n_676), .Y(n_704) );
NAND5xp2_ASAP7_75t_L g679 ( .A(n_680), .B(n_707), .C(n_721), .D(n_732), .E(n_745), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B(n_690), .C(n_703), .Y(n_680) );
INVx2_ASAP7_75t_SL g727 ( .A(n_681), .Y(n_727) );
NAND4xp25_ASAP7_75t_SL g683 ( .A(n_684), .B(n_686), .C(n_687), .D(n_689), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_689), .A2(n_691), .B(n_694), .C(n_700), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_692), .A2(n_733), .B1(n_735), .B2(n_737), .C(n_739), .Y(n_732) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI221xp5_ASAP7_75t_SL g707 ( .A1(n_708), .A2(n_709), .B1(n_712), .B2(n_714), .C(n_716), .Y(n_707) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_715), .A2(n_738), .B1(n_740), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_724) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
endmodule