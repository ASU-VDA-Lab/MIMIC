module fake_netlist_1_7423_n_695 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_695);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_695;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g80 ( .A(n_74), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_78), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_62), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_19), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_42), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_16), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_15), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_23), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_69), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_32), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_37), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_36), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_34), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_70), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_51), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_1), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_20), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_2), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_68), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_5), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_13), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_76), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_53), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_64), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_12), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_10), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_55), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_46), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_14), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_21), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_52), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_60), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_41), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_21), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_29), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_38), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_49), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_43), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_45), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_15), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_77), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_95), .Y(n_130) );
NOR2xp33_ASAP7_75t_R g131 ( .A(n_80), .B(n_27), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_128), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_104), .B(n_0), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_104), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_109), .A2(n_26), .B(n_75), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_120), .B(n_0), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_108), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_121), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_111), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_112), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_123), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_115), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_109), .A2(n_28), .B(n_73), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_83), .B(n_2), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_86), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_129), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_93), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_87), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_84), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_97), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_122), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_89), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_97), .B(n_3), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_107), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_98), .B(n_4), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_94), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_85), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_94), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_85), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_88), .Y(n_171) );
NAND2xp33_ASAP7_75t_SL g172 ( .A(n_98), .B(n_6), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_88), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_114), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_134), .B(n_127), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_166), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_159), .B(n_105), .C(n_99), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_163), .B(n_90), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_134), .B(n_105), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_163), .B(n_90), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_170), .B(n_127), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_163), .B(n_126), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_170), .A2(n_106), .B1(n_99), .B2(n_100), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_146), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_158), .B(n_119), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_153), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_158), .B(n_106), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_153), .B(n_126), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_159), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_164), .B(n_174), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_153), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_141), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_155), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g212 ( .A(n_172), .B(n_101), .C(n_102), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_139), .B(n_116), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_130), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_173), .B(n_116), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_139), .B(n_125), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_169), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_169), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_132), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_168), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_169), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_140), .B(n_119), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_168), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_132), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_138), .B(n_125), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_154), .B(n_124), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_132), .Y(n_229) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_140), .A2(n_110), .B1(n_118), .B2(n_92), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_166), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_143), .B(n_103), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_143), .B(n_124), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_130), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_132), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_166), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_166), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_148), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_148), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_238), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_234), .B(n_142), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
NAND2x1p5_ASAP7_75t_L g244 ( .A(n_190), .B(n_133), .Y(n_244) );
AND2x6_ASAP7_75t_L g245 ( .A(n_217), .B(n_96), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_199), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_183), .B(n_156), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_238), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_203), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_215), .Y(n_250) );
INVxp33_ASAP7_75t_L g251 ( .A(n_186), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_215), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_190), .A2(n_138), .B1(n_161), .B2(n_173), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_227), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_230), .A2(n_171), .B1(n_167), .B2(n_160), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_227), .B(n_151), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_183), .B(n_142), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_202), .B(n_171), .Y(n_261) );
OAI221xp5_ASAP7_75t_L g262 ( .A1(n_191), .A2(n_165), .B1(n_151), .B2(n_167), .C(n_160), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_202), .B(n_157), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_180), .Y(n_265) );
INVx6_ASAP7_75t_L g266 ( .A(n_221), .Y(n_266) );
NOR2x1_ASAP7_75t_L g267 ( .A(n_178), .B(n_165), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_187), .B(n_157), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_203), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_227), .B(n_197), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_227), .B(n_149), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_176), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_199), .B(n_149), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_182), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_179), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_182), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_179), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_214), .B(n_150), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_185), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_228), .B(n_148), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_185), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_212), .A2(n_161), .B1(n_91), .B2(n_117), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_217), .B(n_131), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_214), .B(n_150), .Y(n_288) );
NOR3xp33_ASAP7_75t_SL g289 ( .A(n_209), .B(n_118), .C(n_113), .Y(n_289) );
NOR3xp33_ASAP7_75t_SL g290 ( .A(n_209), .B(n_113), .C(n_110), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_189), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_175), .B(n_92), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_199), .B(n_96), .Y(n_293) );
NOR3xp33_ASAP7_75t_SL g294 ( .A(n_205), .B(n_103), .C(n_152), .Y(n_294) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_208), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_203), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_180), .Y(n_297) );
OR2x4_ASAP7_75t_L g298 ( .A(n_188), .B(n_94), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_189), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_180), .B(n_150), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
INVx3_ASAP7_75t_SL g302 ( .A(n_203), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_207), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_195), .Y(n_304) );
BUFx12f_ASAP7_75t_L g305 ( .A(n_184), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_184), .B(n_137), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_213), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_184), .B(n_137), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_232), .B(n_137), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_305), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_265), .B(n_192), .Y(n_311) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_257), .B(n_204), .C(n_233), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_295), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_259), .B(n_230), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_297), .B(n_200), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_255), .A2(n_224), .B1(n_218), .B2(n_223), .C(n_220), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_268), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_295), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_297), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_250), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_286), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_302), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_249), .Y(n_328) );
NOR2x1_ASAP7_75t_SL g329 ( .A(n_271), .B(n_218), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_297), .B(n_230), .Y(n_331) );
CKINVDCx14_ASAP7_75t_R g332 ( .A(n_241), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_260), .Y(n_333) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_256), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_259), .B(n_230), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_251), .B(n_194), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_308), .A2(n_194), .B(n_213), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_254), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_271), .B(n_203), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_240), .Y(n_345) );
OAI21x1_ASAP7_75t_SL g346 ( .A1(n_257), .A2(n_220), .B(n_223), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_275), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_259), .B(n_201), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_270), .B(n_200), .Y(n_349) );
CKINVDCx6p67_ASAP7_75t_R g350 ( .A(n_245), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_278), .Y(n_351) );
HAxp5_ASAP7_75t_L g352 ( .A(n_262), .B(n_6), .CON(n_352), .SN(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_280), .Y(n_353) );
O2A1O1Ixp5_ASAP7_75t_L g354 ( .A1(n_300), .A2(n_229), .B(n_235), .C(n_198), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_253), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_249), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_242), .B(n_235), .Y(n_357) );
BUFx12f_ASAP7_75t_L g358 ( .A(n_253), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_240), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_298), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_251), .B(n_239), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_270), .B(n_239), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_282), .Y(n_363) );
BUFx8_ASAP7_75t_SL g364 ( .A(n_247), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
NAND2xp33_ASAP7_75t_R g366 ( .A(n_331), .B(n_300), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_317), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_342), .A2(n_306), .B(n_276), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_331), .A2(n_245), .B1(n_252), .B2(n_243), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_333), .A2(n_294), .B1(n_274), .B2(n_285), .C(n_261), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_331), .A2(n_245), .B1(n_281), .B2(n_288), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_317), .B(n_264), .Y(n_374) );
NAND2xp33_ASAP7_75t_R g375 ( .A(n_331), .B(n_306), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_276), .B(n_273), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_331), .A2(n_272), .B1(n_281), .B2(n_288), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_310), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_315), .B(n_245), .Y(n_382) );
AO31x2_ASAP7_75t_L g383 ( .A1(n_321), .A2(n_283), .A3(n_293), .B(n_301), .Y(n_383) );
AOI21xp5_ASAP7_75t_SL g384 ( .A1(n_326), .A2(n_281), .B(n_288), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_333), .A2(n_245), .B1(n_287), .B2(n_267), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_312), .A2(n_291), .B1(n_304), .B2(n_299), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_311), .B(n_249), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_321), .A2(n_309), .B(n_283), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_350), .A2(n_292), .B1(n_244), .B2(n_284), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_324), .A2(n_289), .B1(n_290), .B2(n_244), .C(n_246), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_310), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_311), .A2(n_246), .B1(n_298), .B2(n_296), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_315), .B(n_246), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_312), .A2(n_229), .B1(n_279), .B2(n_277), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_328), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_311), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_389), .A2(n_354), .B(n_346), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_372), .A2(n_332), .B1(n_355), .B2(n_358), .Y(n_402) );
NOR2xp33_ASAP7_75t_SL g403 ( .A(n_379), .B(n_350), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_385), .B(n_352), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_338), .B1(n_311), .B2(n_319), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_374), .A2(n_358), .B1(n_364), .B2(n_339), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_391), .A2(n_371), .B1(n_382), .B2(n_373), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_335), .B1(n_336), .B2(n_319), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_367), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_365), .B(n_352), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_376), .A2(n_352), .B1(n_363), .B2(n_353), .C1(n_334), .C2(n_320), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_378), .Y(n_414) );
INVx4_ASAP7_75t_R g415 ( .A(n_369), .Y(n_415) );
OAI21x1_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_346), .B(n_309), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_390), .A2(n_361), .B1(n_363), .B2(n_360), .Y(n_417) );
OAI221xp5_ASAP7_75t_SL g418 ( .A1(n_386), .A2(n_348), .B1(n_360), .B2(n_325), .C(n_336), .Y(n_418) );
OAI21xp33_ASAP7_75t_SL g419 ( .A1(n_384), .A2(n_325), .B(n_335), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_369), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_392), .B(n_337), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_366), .A2(n_362), .B1(n_337), .B2(n_316), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_368), .Y(n_424) );
OR2x6_ASAP7_75t_L g425 ( .A(n_388), .B(n_318), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_396), .Y(n_426) );
OAI33xp33_ASAP7_75t_L g427 ( .A1(n_399), .A2(n_314), .A3(n_322), .B1(n_337), .B2(n_330), .B3(n_340), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_387), .A2(n_318), .B1(n_340), .B2(n_313), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_412), .B(n_383), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_402), .A2(n_393), .B1(n_380), .B2(n_394), .C(n_387), .Y(n_432) );
AOI31xp33_ASAP7_75t_L g433 ( .A1(n_407), .A2(n_375), .A3(n_366), .B(n_318), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_403), .A2(n_375), .B1(n_329), .B2(n_323), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_405), .Y(n_435) );
INVxp33_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_424), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_415), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_412), .A2(n_395), .B1(n_377), .B2(n_357), .C(n_397), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_403), .A2(n_329), .B1(n_323), .B2(n_326), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_420), .B(n_313), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_404), .B(n_383), .Y(n_442) );
OA222x2_ASAP7_75t_L g443 ( .A1(n_425), .A2(n_419), .B1(n_415), .B2(n_413), .C1(n_418), .C2(n_414), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_414), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_421), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_413), .A2(n_397), .B1(n_357), .B2(n_330), .Y(n_446) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_423), .A2(n_326), .B1(n_327), .B2(n_316), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_422), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_421), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_427), .A2(n_357), .B1(n_279), .B2(n_277), .Y(n_451) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_428), .A2(n_359), .B(n_345), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_426), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_404), .B(n_357), .Y(n_455) );
NOR4xp25_ASAP7_75t_SL g456 ( .A(n_419), .B(n_383), .C(n_8), .D(n_9), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_417), .B(n_94), .C(n_221), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_406), .A2(n_344), .B1(n_327), .B2(n_341), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_409), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_408), .A2(n_359), .B1(n_345), .B2(n_341), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_428), .A2(n_341), .B1(n_327), .B2(n_344), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_410), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_445), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_442), .B(n_411), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_432), .A2(n_423), .B1(n_425), .B2(n_401), .C(n_94), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_437), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_430), .B(n_383), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_430), .B(n_401), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_445), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_464), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_442), .B(n_401), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_449), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_441), .Y(n_477) );
AOI31xp33_ASAP7_75t_L g478 ( .A1(n_434), .A2(n_411), .A3(n_344), .B(n_10), .Y(n_478) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_435), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_444), .B(n_454), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_464), .Y(n_481) );
AOI33xp33_ASAP7_75t_L g482 ( .A1(n_449), .A2(n_181), .A3(n_198), .B1(n_210), .B2(n_219), .B3(n_222), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_448), .B(n_401), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_431), .B(n_411), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_436), .A2(n_425), .B1(n_416), .B2(n_398), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_453), .A2(n_425), .B1(n_248), .B2(n_211), .C(n_221), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_448), .B(n_416), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_431), .Y(n_489) );
OAI33xp33_ASAP7_75t_L g490 ( .A1(n_450), .A2(n_7), .A3(n_9), .B1(n_11), .B2(n_13), .B3(n_14), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_429), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_429), .B(n_425), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_458), .B(n_7), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_458), .B(n_11), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_431), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_443), .B(n_16), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_431), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_460), .B(n_17), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_436), .A2(n_398), .B1(n_367), .B2(n_344), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_463), .B(n_17), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_433), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_446), .A2(n_248), .B1(n_211), .B2(n_226), .C(n_221), .Y(n_504) );
OAI31xp33_ASAP7_75t_L g505 ( .A1(n_447), .A2(n_18), .A3(n_19), .B(n_20), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_455), .B(n_18), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_439), .A2(n_398), .B1(n_367), .B2(n_341), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_463), .Y(n_509) );
AO31x2_ASAP7_75t_L g510 ( .A1(n_452), .A2(n_222), .A3(n_210), .B(n_219), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_463), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_452), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_452), .B(n_398), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_457), .B(n_225), .C(n_181), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g515 ( .A1(n_440), .A2(n_22), .B1(n_356), .B2(n_328), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_470), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_465), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_494), .B(n_461), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_479), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_472), .B(n_456), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_494), .B(n_462), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_474), .Y(n_522) );
INVx5_ASAP7_75t_L g523 ( .A(n_467), .Y(n_523) );
NOR2xp33_ASAP7_75t_R g524 ( .A(n_467), .B(n_468), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_471), .B(n_22), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_499), .B(n_459), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_471), .B(n_451), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_493), .Y(n_529) );
INVx3_ASAP7_75t_SL g530 ( .A(n_467), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_472), .B(n_24), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_499), .B(n_25), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_496), .B(n_177), .C(n_193), .Y(n_533) );
AND3x1_ASAP7_75t_L g534 ( .A(n_496), .B(n_30), .C(n_31), .Y(n_534) );
OR2x6_ASAP7_75t_L g535 ( .A(n_503), .B(n_356), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_466), .B(n_33), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_467), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_468), .B(n_328), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_466), .B(n_35), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_466), .B(n_39), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_476), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_466), .B(n_40), .Y(n_542) );
NOR2xp33_ASAP7_75t_R g543 ( .A(n_468), .B(n_44), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_502), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_513), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_476), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_515), .A2(n_356), .B1(n_328), .B2(n_221), .Y(n_547) );
AND2x4_ASAP7_75t_SL g548 ( .A(n_502), .B(n_356), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_475), .B(n_47), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_475), .B(n_50), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_513), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_474), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_488), .B(n_54), .Y(n_553) );
OAI211xp5_ASAP7_75t_L g554 ( .A1(n_505), .A2(n_221), .B(n_226), .C(n_225), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_493), .Y(n_556) );
BUFx12f_ASAP7_75t_L g557 ( .A(n_492), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_480), .B(n_56), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_481), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_491), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_492), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_483), .B(n_58), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_481), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_477), .B(n_61), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g566 ( .A1(n_478), .A2(n_296), .B(n_269), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_507), .B(n_63), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_512), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_533), .B(n_490), .C(n_554), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_566), .A2(n_505), .B(n_469), .C(n_486), .Y(n_570) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_519), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_534), .A2(n_515), .B1(n_485), .B2(n_508), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_530), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_532), .A2(n_504), .B(n_512), .C(n_509), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_516), .B(n_500), .C(n_511), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_530), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_529), .B(n_489), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_526), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_556), .B(n_506), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_527), .B(n_506), .Y(n_582) );
AOI321xp33_ASAP7_75t_L g583 ( .A1(n_527), .A2(n_513), .A3(n_495), .B1(n_511), .B2(n_498), .C(n_484), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_541), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_522), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_523), .B(n_513), .Y(n_586) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_525), .A2(n_497), .B(n_495), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_532), .B(n_498), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_561), .B(n_484), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_520), .B(n_482), .C(n_514), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_523), .B(n_484), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_547), .A2(n_501), .B(n_484), .Y(n_592) );
INVx2_ASAP7_75t_SL g593 ( .A(n_523), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_523), .A2(n_501), .B(n_510), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_546), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_544), .B(n_510), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_565), .B(n_66), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_543), .B(n_296), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_560), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_552), .B(n_72), .Y(n_601) );
OAI22xp33_ASAP7_75t_SL g602 ( .A1(n_537), .A2(n_226), .B1(n_266), .B2(n_79), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_520), .A2(n_226), .B1(n_193), .B2(n_196), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_521), .A2(n_226), .B1(n_263), .B2(n_269), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_528), .B(n_226), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_568), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_539), .A2(n_269), .B(n_263), .C(n_249), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_563), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_559), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_559), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_518), .A2(n_236), .B1(n_237), .B2(n_196), .C(n_231), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_557), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_572), .B(n_549), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_571), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_606), .Y(n_615) );
AOI21xp33_ASAP7_75t_SL g616 ( .A1(n_599), .A2(n_531), .B(n_549), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_583), .B(n_524), .Y(n_617) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_599), .A2(n_593), .B(n_569), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_574), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_609), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_582), .B(n_531), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_578), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_584), .Y(n_625) );
BUFx2_ASAP7_75t_L g626 ( .A(n_586), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_595), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_582), .B(n_545), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_596), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_581), .B(n_545), .Y(n_630) );
NOR4xp25_ASAP7_75t_SL g631 ( .A(n_612), .B(n_543), .C(n_524), .D(n_535), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_579), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_573), .B(n_551), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_575), .A2(n_539), .B(n_564), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_586), .B(n_553), .Y(n_635) );
NOR3xp33_ASAP7_75t_SL g636 ( .A(n_570), .B(n_590), .C(n_575), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_585), .Y(n_637) );
INVx4_ASAP7_75t_L g638 ( .A(n_601), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_602), .B(n_567), .C(n_558), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_591), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_587), .A2(n_551), .B1(n_550), .B2(n_553), .C(n_539), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_600), .B(n_551), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_591), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_569), .A2(n_553), .B(n_542), .C(n_540), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_589), .B(n_535), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_608), .B(n_535), .Y(n_647) );
O2A1O1Ixp5_ASAP7_75t_SL g648 ( .A1(n_618), .A2(n_605), .B(n_604), .C(n_562), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_615), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_623), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_633), .A2(n_588), .B1(n_577), .B2(n_597), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_617), .B(n_607), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_624), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_634), .B(n_603), .C(n_592), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_619), .Y(n_655) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_635), .B(n_536), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_625), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_636), .B(n_594), .C(n_611), .Y(n_658) );
XNOR2x2_ASAP7_75t_L g659 ( .A(n_617), .B(n_598), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_627), .Y(n_660) );
BUFx3_ASAP7_75t_L g661 ( .A(n_626), .Y(n_661) );
NAND2xp33_ASAP7_75t_SL g662 ( .A(n_631), .B(n_610), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_645), .A2(n_607), .B1(n_538), .B2(n_548), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_614), .B(n_538), .Y(n_665) );
XOR2x2_ASAP7_75t_L g666 ( .A(n_659), .B(n_635), .Y(n_666) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_652), .A2(n_632), .B1(n_622), .B2(n_637), .C1(n_642), .C2(n_644), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_654), .A2(n_641), .B1(n_640), .B2(n_639), .C(n_628), .Y(n_668) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_655), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_656), .A2(n_616), .B1(n_621), .B2(n_638), .Y(n_670) );
NOR2xp33_ASAP7_75t_R g671 ( .A(n_662), .B(n_638), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_664), .A2(n_630), .B(n_646), .C(n_613), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_651), .B(n_643), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_661), .B(n_647), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_658), .A2(n_620), .B(n_237), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_650), .B(n_177), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_653), .Y(n_677) );
AO22x2_ASAP7_75t_L g678 ( .A1(n_657), .A2(n_660), .B1(n_663), .B2(n_665), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_648), .A2(n_656), .B1(n_661), .B2(n_617), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_649), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_652), .B(n_654), .C(n_658), .D(n_496), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_671), .B(n_666), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_669), .B(n_674), .Y(n_683) );
OR3x2_ASAP7_75t_L g684 ( .A(n_681), .B(n_679), .C(n_667), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_668), .A2(n_670), .B1(n_672), .B2(n_673), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_677), .B(n_680), .Y(n_686) );
NAND3x1_ASAP7_75t_L g687 ( .A(n_685), .B(n_669), .C(n_675), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_686), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_682), .B(n_678), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_688), .B(n_683), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_689), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_690), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_691), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_692), .A2(n_684), .B1(n_687), .B2(n_678), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_693), .B(n_676), .Y(n_695) );
endmodule