module real_aes_2935_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_22;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_8;
wire n_10;
AOI32xp33_ASAP7_75t_L g7 ( .A1(n_0), .A2(n_5), .A3(n_8), .B1(n_14), .B2(n_15), .Y(n_7) );
INVxp33_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NAND3xp33_ASAP7_75t_SL g17 ( .A(n_1), .B(n_18), .C(n_19), .Y(n_17) );
INVx3_ASAP7_75t_L g21 ( .A(n_2), .Y(n_21) );
INVx1_ASAP7_75t_L g18 ( .A(n_3), .Y(n_18) );
INVx1_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_4), .B(n_10), .Y(n_22) );
OAI21xp33_ASAP7_75t_SL g15 ( .A1(n_5), .A2(n_10), .B(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_9), .B(n_10), .Y(n_8) );
AOI21xp5_ASAP7_75t_SL g16 ( .A1(n_10), .A2(n_17), .B(n_22), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
INVx2_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
endmodule