module fake_jpeg_18120_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_27),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_26),
.B(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_2),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_19),
.B1(n_11),
.B2(n_13),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_20),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_25),
.B(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_19),
.B1(n_13),
.B2(n_11),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_41),
.B1(n_28),
.B2(n_12),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_11),
.B1(n_22),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_52),
.B1(n_57),
.B2(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_51),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_25),
.B(n_20),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_53),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_39),
.B(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_6),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_43),
.B1(n_42),
.B2(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_7),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_10),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_79),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_49),
.B1(n_57),
.B2(n_50),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_51),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_77),
.B(n_70),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_83),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_62),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_70),
.C(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_86),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_69),
.C(n_47),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_75),
.B(n_78),
.C(n_64),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_7),
.B(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_49),
.B1(n_71),
.B2(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_73),
.B1(n_46),
.B2(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_68),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_100),
.B(n_97),
.C(n_88),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_87),
.B(n_88),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_8),
.B(n_10),
.Y(n_102)
);


endmodule