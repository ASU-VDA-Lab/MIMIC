module real_jpeg_2211_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_25),
.C(n_38),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_7),
.B(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_7),
.B(n_23),
.C(n_30),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_54),
.C(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_7),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_7),
.B(n_58),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_7),
.B(n_65),
.Y(n_126)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_92),
.B1(n_143),
.B2(n_144),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_12),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_91),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_82),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_82),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_61),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_46),
.B2(n_60),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_35),
.B2(n_45),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_19),
.A2(n_20),
.B1(n_64),
.B2(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_19),
.A2(n_20),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_19),
.A2(n_64),
.B(n_72),
.C(n_134),
.Y(n_137)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_51),
.C(n_89),
.Y(n_88)
);

AO21x2_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_22)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

OA22x2_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_102),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_30),
.B(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_35),
.A2(n_45),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

AO21x2_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_44),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

AOI211xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_64),
.B(n_71),
.C(n_72),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_51),
.B1(n_89),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_51),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_50),
.A2(n_51),
.B1(n_100),
.B2(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_51),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_51),
.B(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_73),
.C(n_118),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_58),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_54),
.B(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_74),
.B2(n_75),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_73),
.B1(n_76),
.B2(n_81),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_64),
.A2(n_73),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_64),
.A2(n_73),
.B1(n_111),
.B2(n_112),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_64),
.A2(n_73),
.B1(n_99),
.B2(n_140),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B(n_70),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_69),
.Y(n_68)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_95),
.C(n_99),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_84),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_85),
.A2(n_86),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_106),
.B(n_142),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_103),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_136),
.B(n_141),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_130),
.B(n_135),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_120),
.B(n_129),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_114),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_138),
.Y(n_141)
);


endmodule