module fake_jpeg_3054_n_486 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_486);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_486;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx8_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_52),
.B(n_84),
.Y(n_122)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_53),
.Y(n_133)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_88),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_14),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_28),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_45),
.B1(n_30),
.B2(n_36),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_114),
.B1(n_115),
.B2(n_125),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_61),
.A2(n_45),
.B1(n_30),
.B2(n_36),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_38),
.B1(n_31),
.B2(n_39),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_27),
.B1(n_42),
.B2(n_22),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_116),
.B(n_140),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_22),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_59),
.B(n_37),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_57),
.A2(n_44),
.B1(n_28),
.B2(n_37),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_54),
.A2(n_23),
.B1(n_26),
.B2(n_39),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_126),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_55),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_151),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_27),
.B1(n_42),
.B2(n_35),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_39),
.B(n_26),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_44),
.B1(n_28),
.B2(n_35),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_63),
.B(n_44),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_65),
.A2(n_66),
.B1(n_93),
.B2(n_92),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_83),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_103),
.A2(n_94),
.B1(n_67),
.B2(n_69),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

BUFx4f_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_95),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_157),
.B(n_159),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_158),
.B(n_174),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_82),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_87),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_96),
.B(n_64),
.CI(n_73),
.CON(n_162),
.SN(n_162)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_162),
.B(n_188),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_77),
.B1(n_89),
.B2(n_86),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_91),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_80),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_167),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_97),
.A2(n_79),
.B1(n_78),
.B2(n_75),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_153),
.B1(n_165),
.B2(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_99),
.A2(n_25),
.B1(n_71),
.B2(n_72),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_171),
.A2(n_193),
.B1(n_200),
.B2(n_209),
.Y(n_246)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_0),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_197),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_34),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_106),
.C(n_104),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_134),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_113),
.B(n_2),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_190),
.Y(n_229)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_191),
.Y(n_225)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_202),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_111),
.A2(n_25),
.B1(n_29),
.B2(n_34),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_25),
.B(n_29),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_100),
.B(n_141),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_196),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_2),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_134),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_201),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_126),
.A2(n_34),
.B1(n_29),
.B2(n_24),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_199),
.A2(n_128),
.B1(n_102),
.B2(n_24),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_203),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_112),
.B(n_146),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_129),
.B(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_141),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_111),
.A2(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_236),
.B1(n_255),
.B2(n_257),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_230),
.B(n_167),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_100),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_234),
.C(n_167),
.Y(n_263)
);

OAI22x1_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_157),
.B1(n_164),
.B2(n_162),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_219),
.A2(n_162),
.B1(n_160),
.B2(n_205),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_104),
.B1(n_131),
.B2(n_128),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_222),
.A2(n_187),
.B1(n_183),
.B2(n_184),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_224),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_106),
.B(n_149),
.C(n_102),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_121),
.B1(n_105),
.B2(n_131),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_155),
.B(n_149),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_141),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g244 ( 
.A1(n_180),
.A2(n_102),
.B1(n_121),
.B2(n_105),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_256),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_204),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_253),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_163),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_159),
.B(n_3),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_197),
.A2(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

NOR2x1_ASAP7_75t_R g335 ( 
.A(n_259),
.B(n_278),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_213),
.A2(n_199),
.B(n_177),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_260),
.A2(n_282),
.B(n_293),
.C(n_249),
.Y(n_316)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_291),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_165),
.B(n_201),
.C(n_166),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_286),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_275),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_269),
.A2(n_283),
.B1(n_210),
.B2(n_229),
.Y(n_326)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_173),
.C(n_176),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_234),
.C(n_223),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_175),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_276),
.B(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_245),
.A2(n_177),
.B(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_238),
.B(n_208),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_219),
.A2(n_250),
.B1(n_226),
.B2(n_245),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_295),
.B1(n_261),
.B2(n_296),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_221),
.A2(n_190),
.B(n_156),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_226),
.A2(n_189),
.B1(n_192),
.B2(n_185),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_235),
.B(n_156),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_285),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_214),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_202),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_215),
.B(n_191),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_210),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_290),
.Y(n_319)
);

NAND2x1_ASAP7_75t_SL g289 ( 
.A(n_221),
.B(n_203),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g333 ( 
.A(n_289),
.B(n_227),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_235),
.B(n_186),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_254),
.A2(n_3),
.B(n_5),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_294),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_230),
.A2(n_6),
.B(n_7),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_212),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_7),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_251),
.Y(n_331)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_299),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_229),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_300),
.Y(n_309)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_301),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_273),
.A2(n_244),
.B1(n_212),
.B2(n_223),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_304),
.A2(n_315),
.B1(n_337),
.B2(n_338),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_317),
.C(n_325),
.Y(n_342)
);

OAI32xp33_ASAP7_75t_L g313 ( 
.A1(n_273),
.A2(n_256),
.A3(n_212),
.B1(n_236),
.B2(n_244),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_318),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_259),
.B1(n_261),
.B2(n_290),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_243),
.C(n_224),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_271),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_321),
.B(n_276),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_285),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_331),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_272),
.A2(n_246),
.B1(n_249),
.B2(n_243),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_216),
.C(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_271),
.B1(n_280),
.B2(n_260),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_328),
.A2(n_297),
.B1(n_299),
.B2(n_292),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_216),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_330),
.C(n_339),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_257),
.C(n_229),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_333),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_259),
.A2(n_255),
.B1(n_227),
.B2(n_251),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_293),
.A2(n_253),
.B1(n_225),
.B2(n_252),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_240),
.C(n_237),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_341),
.A2(n_343),
.B1(n_346),
.B2(n_348),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_302),
.A2(n_265),
.B1(n_264),
.B2(n_297),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_328),
.A2(n_265),
.B(n_289),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_345),
.A2(n_350),
.B(n_360),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_264),
.B(n_282),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_306),
.A2(n_277),
.B1(n_279),
.B2(n_284),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_321),
.A2(n_289),
.B(n_278),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_353),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_307),
.B(n_291),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_270),
.B1(n_266),
.B2(n_295),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_355),
.A2(n_320),
.B1(n_309),
.B2(n_312),
.Y(n_397)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_301),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_363),
.C(n_325),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_335),
.A2(n_294),
.B(n_267),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_287),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_366),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_298),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_258),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_262),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_312),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_369),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_315),
.A2(n_269),
.B1(n_283),
.B2(n_288),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_370),
.A2(n_326),
.B1(n_309),
.B2(n_324),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_288),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_371),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_333),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_311),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_379),
.C(n_380),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_381),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_363),
.C(n_368),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_377),
.C(n_386),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_317),
.C(n_305),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_359),
.B(n_330),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_339),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_331),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_344),
.A2(n_304),
.B1(n_316),
.B2(n_319),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_385),
.A2(n_387),
.B1(n_396),
.B2(n_397),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_332),
.C(n_334),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_344),
.A2(n_335),
.B1(n_334),
.B2(n_332),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_391),
.A2(n_393),
.B1(n_356),
.B2(n_364),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_349),
.A2(n_313),
.B1(n_320),
.B2(n_303),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_333),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_350),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_344),
.A2(n_352),
.B1(n_343),
.B2(n_372),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_349),
.A2(n_314),
.B1(n_240),
.B2(n_237),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_401),
.A2(n_403),
.B1(n_396),
.B2(n_387),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_393),
.A2(n_364),
.B1(n_346),
.B2(n_370),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_354),
.C(n_345),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_412),
.C(n_415),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_382),
.A2(n_347),
.B1(n_346),
.B2(n_371),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_407),
.A2(n_409),
.B1(n_417),
.B2(n_389),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_382),
.A2(n_347),
.B1(n_366),
.B2(n_365),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_410),
.B(n_411),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_379),
.B(n_351),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_369),
.C(n_361),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_358),
.C(n_357),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_394),
.A2(n_355),
.B1(n_314),
.B2(n_353),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_416),
.B(n_383),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_385),
.A2(n_220),
.B1(n_225),
.B2(n_10),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_8),
.B(n_9),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_418),
.A2(n_378),
.B(n_376),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_8),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_9),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_397),
.Y(n_421)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_421),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_429),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_426),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_403),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_399),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_401),
.A2(n_381),
.B1(n_386),
.B2(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_431),
.Y(n_442)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_409),
.Y(n_432)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_414),
.A2(n_395),
.B1(n_10),
.B2(n_11),
.Y(n_433)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_9),
.CI(n_12),
.CON(n_435),
.SN(n_435)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_436),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_418),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_417),
.Y(n_437)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_12),
.B(n_13),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_405),
.Y(n_448)
);

INVx11_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_452),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_428),
.B1(n_426),
.B2(n_437),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_402),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_451),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_402),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_412),
.C(n_400),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_414),
.Y(n_453)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_453),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_450),
.B(n_425),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_455),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_440),
.Y(n_455)
);

FAx1_ASAP7_75t_SL g456 ( 
.A(n_446),
.B(n_438),
.CI(n_410),
.CON(n_456),
.SN(n_456)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_463),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_442),
.A2(n_406),
.B(n_427),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_458),
.A2(n_452),
.B(n_400),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_427),
.B(n_432),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_459),
.A2(n_445),
.B(n_444),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_460),
.A2(n_449),
.B1(n_448),
.B2(n_447),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_443),
.A2(n_433),
.B1(n_439),
.B2(n_425),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_466),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_472),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_456),
.B(n_408),
.CI(n_438),
.CON(n_469),
.SN(n_469)
);

NOR3xp33_ASAP7_75t_SL g474 ( 
.A(n_469),
.B(n_408),
.C(n_456),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_444),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_471),
.B(n_463),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_464),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_476),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_462),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_471),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_462),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_478),
.A2(n_479),
.B(n_470),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_480),
.B(n_473),
.C(n_457),
.Y(n_481)
);

A2O1A1O1Ixp25_ASAP7_75t_L g483 ( 
.A1(n_481),
.A2(n_482),
.B(n_460),
.C(n_469),
.D(n_435),
.Y(n_483)
);

AOI321xp33_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_435),
.A3(n_420),
.B1(n_434),
.B2(n_419),
.C(n_13),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_434),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_485),
.A2(n_12),
.B(n_479),
.Y(n_486)
);


endmodule