module fake_netlist_6_2608_n_1015 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1015);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1015;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_795;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_970;
wire n_849;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_100),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_148),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_70),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_19),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_109),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_129),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_154),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_140),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_90),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_4),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_214),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_153),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_141),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_203),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_56),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_123),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_162),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_118),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_85),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_132),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_137),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_159),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_213),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_142),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_3),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_205),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_80),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_46),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_34),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_98),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_59),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_125),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_57),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_207),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_160),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_9),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_209),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_89),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_64),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_157),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_2),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_107),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_175),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_32),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_105),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_35),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_54),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_189),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_29),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_62),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_65),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_193),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_111),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_127),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_218),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_164),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_5),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_174),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_112),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_225),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_66),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_76),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_20),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_204),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_113),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_84),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_104),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_67),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_40),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_139),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_236),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_226),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_243),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_229),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_230),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_231),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_233),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_271),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_234),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_268),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_238),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_0),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_246),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_0),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_292),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_241),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_1),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_275),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_292),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_247),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_273),
.B(n_1),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_248),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_283),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_227),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_232),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_235),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_2),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_237),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_240),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_305),
.B(n_3),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_242),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_244),
.B(n_4),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_250),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_256),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_262),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_239),
.B(n_249),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_272),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_251),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_252),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_277),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_298),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_255),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_326),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

CKINVDCx8_ASAP7_75t_R g387 ( 
.A(n_359),
.Y(n_387)
);

CKINVDCx8_ASAP7_75t_R g388 ( 
.A(n_328),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_304),
.B(n_253),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_332),
.B(n_318),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_380),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_322),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_362),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_228),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_334),
.B(n_324),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_280),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_289),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_335),
.B(n_323),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_336),
.B(n_254),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_346),
.B(n_306),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_343),
.B(n_257),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_345),
.B(n_316),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_258),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_341),
.B(n_259),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_355),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_261),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_375),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_349),
.B(n_321),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_330),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_330),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_402),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_354),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_405),
.B(n_354),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_385),
.B(n_255),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_351),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_340),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_385),
.B(n_255),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_263),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_393),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_402),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_402),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_340),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_264),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_393),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_418),
.B(n_361),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_399),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_255),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_430),
.A2(n_361),
.B1(n_337),
.B2(n_296),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_431),
.A2(n_255),
.B1(n_320),
.B2(n_319),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_401),
.B(n_255),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_391),
.B(n_265),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_411),
.B(n_266),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_267),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_406),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_391),
.B(n_270),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_274),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_431),
.B(n_5),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_28),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_391),
.B(n_278),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_409),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_388),
.Y(n_483)
);

AO22x2_ASAP7_75t_L g484 ( 
.A1(n_426),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_484)
);

INVx6_ASAP7_75t_L g485 ( 
.A(n_409),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_399),
.B(n_279),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_400),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_421),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_400),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_404),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_388),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_407),
.B(n_281),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_436),
.B(n_282),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_284),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_428),
.B(n_285),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_383),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_392),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_424),
.A2(n_302),
.B1(n_314),
.B2(n_313),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_383),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_429),
.B(n_286),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_424),
.A2(n_301),
.B1(n_312),
.B2(n_310),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_437),
.B(n_290),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_392),
.B(n_291),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_433),
.B(n_31),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_383),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_383),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_424),
.A2(n_300),
.B1(n_309),
.B2(n_308),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_401),
.B(n_294),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_495),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_460),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_501),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_504),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_491),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_493),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_435),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_456),
.B(n_435),
.Y(n_531)
);

OAI221xp5_ASAP7_75t_L g532 ( 
.A1(n_471),
.A2(n_422),
.B1(n_441),
.B2(n_415),
.C(n_416),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_452),
.B(n_437),
.Y(n_533)
);

CKINVDCx11_ASAP7_75t_R g534 ( 
.A(n_489),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_466),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_503),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_483),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_496),
.B(n_437),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_469),
.A2(n_440),
.B1(n_441),
.B2(n_424),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_464),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_469),
.A2(n_440),
.B1(n_424),
.B2(n_401),
.Y(n_542)
);

AO22x2_ASAP7_75t_L g543 ( 
.A1(n_484),
.A2(n_432),
.B1(n_434),
.B2(n_433),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_503),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_478),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_461),
.B(n_403),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_514),
.Y(n_547)
);

OR2x2_ASAP7_75t_SL g548 ( 
.A(n_449),
.B(n_439),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g549 ( 
.A1(n_515),
.A2(n_396),
.B1(n_387),
.B2(n_438),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_461),
.B(n_475),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_451),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_497),
.B(n_427),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_497),
.B(n_412),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_498),
.B(n_414),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_494),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_447),
.Y(n_558)
);

AO22x2_ASAP7_75t_L g559 ( 
.A1(n_484),
.A2(n_325),
.B1(n_419),
.B2(n_8),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_484),
.A2(n_479),
.B1(n_472),
.B2(n_507),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_475),
.B(n_387),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_498),
.B(n_394),
.Y(n_562)
);

AO22x2_ASAP7_75t_L g563 ( 
.A1(n_479),
.A2(n_325),
.B1(n_7),
.B2(n_10),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_472),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_507),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_465),
.B(n_394),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_515),
.B(n_413),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_474),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_568)
);

BUFx8_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_449),
.Y(n_570)
);

AO22x2_ASAP7_75t_L g571 ( 
.A1(n_505),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_505),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_453),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_499),
.B(n_500),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_468),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_465),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_511),
.Y(n_580)
);

OAI221xp5_ASAP7_75t_L g581 ( 
.A1(n_471),
.A2(n_403),
.B1(n_416),
.B2(n_415),
.C(n_384),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_511),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_446),
.B(n_386),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_519),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_508),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_473),
.B(n_417),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_519),
.B(n_423),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_509),
.B(n_423),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_508),
.B(n_295),
.Y(n_591)
);

OAI221xp5_ASAP7_75t_L g592 ( 
.A1(n_518),
.A2(n_303),
.B1(n_297),
.B2(n_417),
.C(n_389),
.Y(n_592)
);

OAI221xp5_ASAP7_75t_L g593 ( 
.A1(n_518),
.A2(n_473),
.B1(n_477),
.B2(n_481),
.C(n_417),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_512),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_482),
.B(n_417),
.Y(n_595)
);

BUFx8_ASAP7_75t_L g596 ( 
.A(n_512),
.Y(n_596)
);

AO22x2_ASAP7_75t_L g597 ( 
.A1(n_512),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_512),
.B(n_417),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_487),
.Y(n_599)
);

BUFx8_ASAP7_75t_L g600 ( 
.A(n_512),
.Y(n_600)
);

BUFx8_ASAP7_75t_L g601 ( 
.A(n_480),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_487),
.Y(n_602)
);

NAND2x1p5_ASAP7_75t_L g603 ( 
.A(n_492),
.B(n_390),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_575),
.B(n_538),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_553),
.B(n_477),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_561),
.B(n_481),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_551),
.B(n_514),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_555),
.B(n_514),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_530),
.B(n_510),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_554),
.B(n_510),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_533),
.B(n_517),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_578),
.B(n_517),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_545),
.B(n_443),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_580),
.B(n_443),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_582),
.B(n_443),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_570),
.B(n_579),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_546),
.B(n_458),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_549),
.B(n_458),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_574),
.B(n_458),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_585),
.B(n_490),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_480),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_558),
.B(n_462),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_541),
.B(n_462),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_524),
.B(n_462),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_557),
.B(n_490),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_SL g626 ( 
.A(n_537),
.B(n_463),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_556),
.B(n_442),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_525),
.B(n_454),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_527),
.B(n_454),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_528),
.B(n_467),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_589),
.B(n_502),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_SL g632 ( 
.A(n_521),
.B(n_513),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_591),
.B(n_480),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_550),
.B(n_455),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_529),
.B(n_457),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_536),
.B(n_457),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_544),
.B(n_459),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_520),
.B(n_522),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_552),
.B(n_480),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_590),
.B(n_506),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_562),
.B(n_523),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_535),
.B(n_506),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_526),
.B(n_506),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_534),
.B(n_480),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_569),
.B(n_485),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_577),
.B(n_506),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_573),
.B(n_516),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_576),
.B(n_516),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_601),
.B(n_516),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_596),
.B(n_516),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_600),
.B(n_566),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_588),
.B(n_389),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_583),
.B(n_389),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_547),
.B(n_389),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_567),
.B(n_390),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_540),
.B(n_485),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_584),
.B(n_485),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_587),
.B(n_33),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_599),
.B(n_36),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_602),
.B(n_37),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_595),
.B(n_38),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_603),
.B(n_39),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_548),
.B(n_41),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_539),
.B(n_24),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_539),
.B(n_42),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_593),
.B(n_44),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_542),
.B(n_47),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_SL g668 ( 
.A(n_560),
.B(n_25),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_605),
.A2(n_598),
.B(n_592),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_609),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_666),
.A2(n_560),
.B1(n_594),
.B2(n_597),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_612),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_617),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_641),
.B(n_542),
.Y(n_674)
);

AO21x2_ASAP7_75t_L g675 ( 
.A1(n_666),
.A2(n_655),
.B(n_667),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_662),
.A2(n_532),
.B(n_581),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_639),
.A2(n_543),
.B(n_594),
.Y(n_677)
);

INVx3_ASAP7_75t_SL g678 ( 
.A(n_651),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_633),
.A2(n_597),
.B(n_543),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_664),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_608),
.A2(n_559),
.B(n_564),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_658),
.B(n_571),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_665),
.A2(n_586),
.B(n_572),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_634),
.A2(n_564),
.B(n_572),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_604),
.B(n_559),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_626),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_616),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_636),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_644),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_621),
.B(n_568),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_637),
.Y(n_691)
);

O2A1O1Ixp5_ASAP7_75t_L g692 ( 
.A1(n_618),
.A2(n_568),
.B(n_565),
.C(n_563),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_658),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_610),
.A2(n_565),
.B(n_563),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_630),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_658),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_645),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_652),
.A2(n_143),
.B(n_223),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_606),
.B(n_48),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_635),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_647),
.A2(n_136),
.B(n_222),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_668),
.A2(n_224),
.B(n_135),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_627),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_619),
.B(n_49),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_663),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_620),
.B(n_50),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_613),
.B(n_26),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_648),
.A2(n_134),
.B(n_215),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_646),
.A2(n_133),
.B(n_212),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_623),
.B(n_26),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_614),
.A2(n_615),
.B1(n_622),
.B2(n_643),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_659),
.A2(n_144),
.B(n_52),
.Y(n_712)
);

OA21x2_ASAP7_75t_L g713 ( 
.A1(n_640),
.A2(n_145),
.B(n_53),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_611),
.B(n_27),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_607),
.A2(n_55),
.B(n_58),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_656),
.A2(n_60),
.B(n_63),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_638),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_624),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_628),
.A2(n_72),
.B(n_73),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_632),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_670),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_705),
.B(n_649),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_680),
.B(n_650),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_657),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_685),
.B(n_689),
.Y(n_725)
);

AO31x2_ASAP7_75t_L g726 ( 
.A1(n_671),
.A2(n_625),
.A3(n_660),
.B(n_661),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_697),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_669),
.A2(n_653),
.B(n_629),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_696),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_676),
.A2(n_642),
.B(n_654),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_696),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_SL g732 ( 
.A1(n_702),
.A2(n_671),
.B(n_674),
.C(n_699),
.Y(n_732)
);

AO31x2_ASAP7_75t_L g733 ( 
.A1(n_679),
.A2(n_631),
.A3(n_75),
.B(n_77),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_701),
.A2(n_74),
.B(n_78),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_696),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_684),
.A2(n_79),
.B(n_81),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_695),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_674),
.A2(n_82),
.A3(n_83),
.B(n_86),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_692),
.A2(n_87),
.B(n_88),
.C(n_91),
.Y(n_739)
);

NAND2x1p5_ASAP7_75t_L g740 ( 
.A(n_717),
.B(n_92),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_708),
.A2(n_93),
.B(n_94),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_709),
.A2(n_95),
.B(n_96),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_693),
.Y(n_743)
);

OR3x4_ASAP7_75t_SL g744 ( 
.A(n_673),
.B(n_99),
.C(n_101),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_672),
.B(n_102),
.Y(n_745)
);

INVx4_ASAP7_75t_SL g746 ( 
.A(n_697),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_716),
.A2(n_103),
.B(n_106),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_707),
.Y(n_748)
);

OAI21x1_ASAP7_75t_SL g749 ( 
.A1(n_702),
.A2(n_108),
.B(n_110),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_686),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_678),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_694),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_688),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_690),
.B(n_117),
.Y(n_754)
);

INVxp33_ASAP7_75t_SL g755 ( 
.A(n_703),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_691),
.Y(n_756)
);

OAI222xp33_ASAP7_75t_L g757 ( 
.A1(n_682),
.A2(n_718),
.B1(n_720),
.B2(n_710),
.C1(n_717),
.C2(n_711),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_711),
.A2(n_119),
.A3(n_120),
.B(n_124),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_683),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_759)
);

OAI21x1_ASAP7_75t_SL g760 ( 
.A1(n_683),
.A2(n_131),
.B(n_146),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_700),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_704),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_714),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_677),
.A2(n_147),
.B(n_150),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_720),
.B(n_151),
.Y(n_765)
);

AOI21x1_ASAP7_75t_L g766 ( 
.A1(n_713),
.A2(n_217),
.B(n_155),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_682),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_704),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_753),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_768),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_756),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_755),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_761),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_768),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_729),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_737),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_743),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_766),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_728),
.A2(n_706),
.B(n_675),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_764),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_758),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_767),
.B(n_681),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_768),
.A2(n_712),
.B1(n_718),
.B2(n_715),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_734),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_721),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_758),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_741),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_742),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_767),
.Y(n_790)
);

AOI21xp33_ASAP7_75t_L g791 ( 
.A1(n_748),
.A2(n_681),
.B(n_675),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_763),
.B(n_706),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_743),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_725),
.B(n_754),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_733),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_758),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_733),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_731),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

AOI21x1_ASAP7_75t_L g800 ( 
.A1(n_728),
.A2(n_719),
.B(n_698),
.Y(n_800)
);

OA21x2_ASAP7_75t_L g801 ( 
.A1(n_736),
.A2(n_152),
.B(n_156),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_727),
.Y(n_802)
);

BUFx12f_ASAP7_75t_L g803 ( 
.A(n_750),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_745),
.Y(n_804)
);

AO21x2_ASAP7_75t_L g805 ( 
.A1(n_736),
.A2(n_158),
.B(n_163),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_729),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_731),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_745),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_738),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_735),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_729),
.B(n_723),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_738),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_738),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_726),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_732),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_749),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_816)
);

AO21x2_ASAP7_75t_L g817 ( 
.A1(n_757),
.A2(n_169),
.B(n_170),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_726),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_726),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_R g821 ( 
.A(n_802),
.B(n_751),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_770),
.B(n_774),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_794),
.B(n_748),
.Y(n_823)
);

AND2x2_ASAP7_75t_SL g824 ( 
.A(n_801),
.B(n_744),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_794),
.B(n_724),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_792),
.B(n_722),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_772),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_804),
.B(n_765),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_786),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_811),
.B(n_765),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_R g831 ( 
.A(n_772),
.B(n_770),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_798),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_R g833 ( 
.A(n_770),
.B(n_774),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_811),
.B(n_762),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_811),
.B(n_762),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_810),
.B(n_740),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_774),
.B(n_746),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_807),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_790),
.B(n_746),
.Y(n_839)
);

XOR2xp5_ASAP7_75t_L g840 ( 
.A(n_819),
.B(n_740),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_790),
.B(n_752),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_810),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_782),
.B(n_730),
.Y(n_843)
);

CKINVDCx16_ASAP7_75t_R g844 ( 
.A(n_803),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_782),
.B(n_730),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_804),
.B(n_759),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_803),
.B(n_757),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_776),
.B(n_739),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_775),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_775),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_793),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_SL g852 ( 
.A(n_817),
.B(n_739),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_806),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_R g854 ( 
.A(n_801),
.B(n_171),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_R g855 ( 
.A(n_801),
.B(n_172),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_808),
.B(n_760),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_815),
.B(n_173),
.Y(n_858)
);

BUFx2_ASAP7_75t_SL g859 ( 
.A(n_776),
.Y(n_859)
);

BUFx10_ASAP7_75t_L g860 ( 
.A(n_771),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_808),
.B(n_176),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_769),
.B(n_177),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_SL g864 ( 
.A(n_817),
.B(n_178),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_R g865 ( 
.A(n_801),
.B(n_179),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_843),
.B(n_796),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_851),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_843),
.B(n_781),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_824),
.A2(n_805),
.B1(n_817),
.B2(n_783),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_825),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_821),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_845),
.B(n_781),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_847),
.A2(n_779),
.B(n_816),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_832),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_845),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_777),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_862),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_838),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_859),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_848),
.B(n_787),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_860),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_842),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_860),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_857),
.Y(n_885)
);

CKINVDCx8_ASAP7_75t_R g886 ( 
.A(n_844),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_828),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_836),
.B(n_787),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_830),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_826),
.B(n_769),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_822),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_863),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_822),
.B(n_796),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_841),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_852),
.B(n_809),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_833),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_SL g897 ( 
.A1(n_858),
.A2(n_805),
.B1(n_815),
.B2(n_809),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_841),
.Y(n_898)
);

BUFx2_ASAP7_75t_SL g899 ( 
.A(n_886),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_875),
.B(n_812),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_896),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_866),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_867),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_875),
.B(n_812),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_867),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_897),
.A2(n_840),
.B1(n_846),
.B2(n_839),
.Y(n_906)
);

AOI31xp33_ASAP7_75t_L g907 ( 
.A1(n_873),
.A2(n_831),
.A3(n_855),
.B(n_865),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_874),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_878),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_883),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_885),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_885),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_887),
.B(n_791),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_868),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_892),
.B(n_864),
.C(n_861),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_869),
.B(n_835),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_902),
.B(n_866),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_902),
.B(n_866),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_902),
.B(n_914),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_914),
.B(n_868),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_903),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_901),
.B(n_889),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_901),
.B(n_877),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_905),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_899),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_903),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_906),
.B(n_884),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_910),
.B(n_870),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_908),
.B(n_882),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_911),
.B(n_880),
.Y(n_930)
);

AO221x2_ASAP7_75t_L g931 ( 
.A1(n_930),
.A2(n_909),
.B1(n_881),
.B2(n_886),
.C(n_907),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_929),
.B(n_930),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_925),
.B(n_871),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_923),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_928),
.B(n_912),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_920),
.B(n_827),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_924),
.B(n_919),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_921),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_934),
.B(n_917),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_933),
.B(n_927),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_932),
.B(n_927),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_931),
.B(n_917),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_937),
.B(n_927),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_938),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_936),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_935),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_934),
.B(n_918),
.Y(n_947)
);

NOR2x1_ASAP7_75t_SL g948 ( 
.A(n_940),
.B(n_916),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_939),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_946),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_945),
.B(n_890),
.Y(n_951)
);

OAI32xp33_ASAP7_75t_L g952 ( 
.A1(n_942),
.A2(n_916),
.A3(n_854),
.B1(n_915),
.B2(n_900),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_951),
.B(n_947),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_949),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_950),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_951),
.B(n_952),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_954),
.B(n_940),
.Y(n_957)
);

BUFx12f_ASAP7_75t_L g958 ( 
.A(n_955),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_956),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_953),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_955),
.Y(n_961)
);

OAI211xp5_ASAP7_75t_SL g962 ( 
.A1(n_959),
.A2(n_943),
.B(n_941),
.C(n_948),
.Y(n_962)
);

NOR3x1_ASAP7_75t_L g963 ( 
.A(n_961),
.B(n_896),
.C(n_944),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_957),
.A2(n_915),
.B(n_884),
.Y(n_964)
);

OAI221xp5_ASAP7_75t_L g965 ( 
.A1(n_960),
.A2(n_884),
.B1(n_913),
.B2(n_876),
.C(n_894),
.Y(n_965)
);

AND4x1_ASAP7_75t_L g966 ( 
.A(n_958),
.B(n_879),
.C(n_834),
.D(n_922),
.Y(n_966)
);

NOR4xp25_ASAP7_75t_SL g967 ( 
.A(n_960),
.B(n_853),
.C(n_879),
.D(n_926),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_959),
.B(n_919),
.Y(n_968)
);

NAND4xp25_ASAP7_75t_L g969 ( 
.A(n_959),
.B(n_898),
.C(n_837),
.D(n_839),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_968),
.Y(n_970)
);

NAND2xp33_ASAP7_75t_R g971 ( 
.A(n_967),
.B(n_180),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_962),
.A2(n_969),
.B1(n_965),
.B2(n_964),
.Y(n_972)
);

AOI222xp33_ASAP7_75t_L g973 ( 
.A1(n_963),
.A2(n_918),
.B1(n_880),
.B2(n_837),
.C1(n_872),
.C2(n_921),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_966),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_962),
.A2(n_891),
.B1(n_872),
.B2(n_893),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_962),
.A2(n_891),
.B(n_813),
.C(n_789),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_L g977 ( 
.A(n_962),
.B(n_893),
.C(n_904),
.Y(n_977)
);

NAND4xp75_ASAP7_75t_L g978 ( 
.A(n_970),
.B(n_888),
.C(n_797),
.D(n_799),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_971),
.A2(n_872),
.B1(n_805),
.B2(n_888),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_974),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_972),
.B(n_895),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_977),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_976),
.B(n_895),
.Y(n_983)
);

NOR2x1_ASAP7_75t_L g984 ( 
.A(n_973),
.B(n_813),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_975),
.B(n_856),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_980),
.B(n_181),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_797),
.C(n_799),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_982),
.B(n_182),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_981),
.B(n_856),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_SL g990 ( 
.A(n_985),
.B(n_850),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_984),
.B(n_183),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_983),
.B(n_184),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_986),
.B(n_978),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_992),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_988),
.Y(n_995)
);

AOI221xp5_ASAP7_75t_L g996 ( 
.A1(n_989),
.A2(n_820),
.B1(n_818),
.B2(n_795),
.C(n_778),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_SL g997 ( 
.A1(n_987),
.A2(n_849),
.B1(n_850),
.B2(n_820),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_991),
.B(n_849),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_998),
.Y(n_999)
);

AOI22x1_ASAP7_75t_L g1000 ( 
.A1(n_994),
.A2(n_995),
.B1(n_990),
.B2(n_993),
.Y(n_1000)
);

OR3x1_ASAP7_75t_L g1001 ( 
.A(n_997),
.B(n_996),
.C(n_818),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_L g1002 ( 
.A1(n_994),
.A2(n_795),
.B1(n_778),
.B2(n_800),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_999),
.A2(n_785),
.B(n_784),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_1000),
.A2(n_780),
.B1(n_814),
.B2(n_784),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_1001),
.A2(n_800),
.B(n_788),
.Y(n_1005)
);

AOI31xp33_ASAP7_75t_L g1006 ( 
.A1(n_1004),
.A2(n_1002),
.A3(n_187),
.B(n_188),
.Y(n_1006)
);

AOI31xp33_ASAP7_75t_L g1007 ( 
.A1(n_1003),
.A2(n_186),
.A3(n_191),
.B(n_192),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_1007),
.A2(n_1005),
.B(n_196),
.C(n_197),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1006),
.A2(n_785),
.B1(n_780),
.B2(n_789),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_1009),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1008),
.A2(n_789),
.B1(n_788),
.B2(n_814),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_1010),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_1011),
.Y(n_1013)
);

AOI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_1012),
.A2(n_195),
.B1(n_198),
.B2(n_200),
.C(n_202),
.Y(n_1014)
);

AOI211xp5_ASAP7_75t_L g1015 ( 
.A1(n_1014),
.A2(n_1013),
.B(n_206),
.C(n_208),
.Y(n_1015)
);


endmodule