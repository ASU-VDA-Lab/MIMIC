module real_jpeg_25979_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_35),
.B1(n_40),
.B2(n_44),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_35),
.B1(n_61),
.B2(n_67),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_3),
.A2(n_35),
.B1(n_55),
.B2(n_59),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_4),
.A2(n_40),
.B1(n_44),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_47),
.B1(n_55),
.B2(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_58),
.B(n_103),
.C(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_47),
.B1(n_62),
.B2(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_4),
.B(n_54),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_4),
.A2(n_59),
.B(n_74),
.C(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_24),
.C(n_43),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_4),
.B(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_32),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_4),
.B(n_45),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_55),
.B1(n_59),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_8),
.A2(n_40),
.B1(n_44),
.B2(n_63),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_63),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_26),
.B1(n_40),
.B2(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_11),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_11),
.B(n_185),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_133),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_131),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_108),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_108),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_80),
.B2(n_81),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_50),
.B2(n_51),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_36),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_29),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_22),
.A2(n_90),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_24),
.B(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_27),
.B(n_89),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_27),
.A2(n_33),
.B(n_89),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_27),
.B(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_30),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_30),
.B(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_48),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_37),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_46),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_38),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_38),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_44),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_40),
.B(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_44),
.A2(n_47),
.B(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_45),
.B(n_153),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_46),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_57),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_48),
.B(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_70),
.B1(n_71),
.B2(n_79),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_59),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_65),
.Y(n_95)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_77),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_72),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_76),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_78),
.B(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_83),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_83),
.B(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_85),
.B(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_87),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_90),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_106),
.Y(n_158)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_114),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_109),
.A2(n_110),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_113),
.Y(n_228)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_125),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_117),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_129),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_229),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_223),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_164),
.B(n_222),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_154),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_137),
.B(n_154),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.C(n_149),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_138),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_141),
.C(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_145),
.B(n_149),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_148),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_158),
.C(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_217),
.B(n_221),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_205),
.B(n_216),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_187),
.B(n_204),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_181),
.B2(n_186),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_180),
.C(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_193),
.B(n_203),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B(n_202),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_207),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);


endmodule