module fake_netlist_6_915_n_898 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_898);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_898;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_844;
wire n_343;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_719;
wire n_565;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_78),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_136),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_77),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_21),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_57),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_122),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_116),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_95),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_23),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_35),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_63),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_133),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_98),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_128),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_96),
.Y(n_237)
);

BUFx2_ASAP7_75t_SL g238 ( 
.A(n_6),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_46),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_115),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_55),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_11),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_184),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_152),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_151),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_105),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_15),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_114),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_125),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_76),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_101),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_80),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_119),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_89),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_166),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_97),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_132),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_47),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_153),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_70),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_68),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_43),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_185),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_59),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_186),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_179),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_196),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_1),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_164),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_117),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_197),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_198),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_212),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_201),
.B(n_0),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_236),
.Y(n_306)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_224),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_1),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_2),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_224),
.B(n_2),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_214),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_3),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_209),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_205),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_208),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_216),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_203),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_244),
.B(n_3),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_206),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_203),
.Y(n_323)
);

BUFx8_ASAP7_75t_SL g324 ( 
.A(n_206),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_210),
.B(n_4),
.Y(n_325)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_204),
.Y(n_326)
);

BUFx8_ASAP7_75t_L g327 ( 
.A(n_252),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_220),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_204),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_256),
.B(n_4),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_219),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_221),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_222),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_5),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_238),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_207),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_231),
.B(n_7),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_237),
.B(n_8),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g342 ( 
.A(n_225),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_207),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_325),
.B1(n_303),
.B2(n_305),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_242),
.B1(n_265),
.B2(n_268),
.Y(n_346)
);

AO22x2_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_297),
.B1(n_314),
.B2(n_310),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_336),
.A2(n_215),
.B1(n_229),
.B2(n_247),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_302),
.A2(n_249),
.B1(n_215),
.B2(n_286),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_R g350 ( 
.A1(n_301),
.A2(n_289),
.B1(n_288),
.B2(n_279),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_302),
.A2(n_229),
.B1(n_286),
.B2(n_249),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_292),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_302),
.A2(n_247),
.B1(n_250),
.B2(n_245),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_310),
.A2(n_240),
.B1(n_251),
.B2(n_259),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_302),
.A2(n_250),
.B1(n_261),
.B2(n_263),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_255),
.B1(n_281),
.B2(n_280),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_199),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_211),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_292),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_287),
.B1(n_278),
.B2(n_277),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_314),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_12),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_303),
.A2(n_276),
.B1(n_272),
.B2(n_271),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_308),
.A2(n_270),
.B1(n_269),
.B2(n_267),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g373 ( 
.A(n_300),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_303),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_303),
.A2(n_264),
.B1(n_262),
.B2(n_258),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_305),
.A2(n_257),
.B1(n_253),
.B2(n_248),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_291),
.Y(n_377)
);

NAND3x1_ASAP7_75t_L g378 ( 
.A(n_309),
.B(n_15),
.C(n_16),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_305),
.A2(n_246),
.B1(n_241),
.B2(n_239),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_L g381 ( 
.A1(n_305),
.A2(n_235),
.B1(n_234),
.B2(n_232),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_320),
.B(n_228),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g383 ( 
.A1(n_292),
.A2(n_226),
.B1(n_218),
.B2(n_213),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_339),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_384)
);

AO22x2_ASAP7_75t_L g385 ( 
.A1(n_341),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_309),
.A2(n_334),
.B1(n_342),
.B2(n_321),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_334),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_293),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_298),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_293),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_293),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_292),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_341),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_300),
.A2(n_330),
.B1(n_296),
.B2(n_316),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_330),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_296),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_320),
.B(n_30),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_348),
.B(n_295),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_379),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_390),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_388),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_324),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_307),
.Y(n_413)
);

INVx4_ASAP7_75t_SL g414 ( 
.A(n_398),
.Y(n_414)
);

AOI21x1_ASAP7_75t_L g415 ( 
.A1(n_382),
.A2(n_316),
.B(n_313),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_296),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_373),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_307),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_386),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_356),
.B(n_307),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_356),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_295),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_355),
.B(n_320),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_371),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_362),
.B(n_296),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_349),
.B(n_324),
.Y(n_431)
);

XOR2x2_ASAP7_75t_L g432 ( 
.A(n_369),
.B(n_335),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_369),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_366),
.B(n_307),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_294),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_367),
.A2(n_311),
.B(n_337),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_358),
.B(n_320),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_335),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_352),
.B(n_340),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_344),
.B(n_323),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_347),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_350),
.B(n_323),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

XOR2x2_ASAP7_75t_L g457 ( 
.A(n_378),
.B(n_327),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_383),
.B(n_304),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_387),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_396),
.B(n_304),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_351),
.B(n_311),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_401),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_313),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_423),
.B(n_304),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_441),
.B(n_337),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_340),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_423),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_417),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_467),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_318),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_414),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_312),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_416),
.B(n_312),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_312),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_317),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_433),
.A2(n_343),
.B(n_323),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_414),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_343),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_433),
.B(n_317),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_439),
.B(n_317),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_31),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_439),
.B(n_318),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_318),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_429),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_413),
.B(n_323),
.Y(n_505)
);

INVx3_ASAP7_75t_SL g506 ( 
.A(n_457),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_463),
.B(n_464),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_454),
.B(n_319),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_427),
.B(n_319),
.Y(n_511)
);

BUFx5_ASAP7_75t_L g512 ( 
.A(n_460),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_459),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_461),
.B(n_319),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_425),
.B(n_326),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_428),
.B(n_331),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_436),
.B(n_331),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_438),
.B(n_440),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_459),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_434),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_442),
.B(n_331),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_444),
.B(n_332),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_445),
.B(n_332),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_448),
.B(n_332),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_449),
.B(n_333),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_402),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_425),
.A2(n_450),
.B(n_456),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_450),
.B(n_424),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_451),
.B(n_333),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_424),
.B(n_326),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_479),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_479),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_L g539 ( 
.A(n_497),
.B(n_426),
.Y(n_539)
);

BUFx8_ASAP7_75t_SL g540 ( 
.A(n_522),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_479),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_493),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g543 ( 
.A(n_471),
.B(n_426),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_471),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_483),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_474),
.B(n_424),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_493),
.Y(n_547)
);

AND2x6_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_458),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_471),
.Y(n_549)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_497),
.B(n_443),
.Y(n_550)
);

NAND2x1_ASAP7_75t_SL g551 ( 
.A(n_513),
.B(n_455),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_474),
.B(n_424),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_493),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_503),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_483),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_463),
.Y(n_556)
);

BUFx12f_ASAP7_75t_L g557 ( 
.A(n_478),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_516),
.B(n_424),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_497),
.B(n_421),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_514),
.B(n_419),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_421),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_476),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_496),
.B(n_435),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_471),
.B(n_326),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_488),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_491),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_521),
.B(n_462),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_471),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_534),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_472),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_491),
.Y(n_575)
);

AND2x2_ASAP7_75t_SL g576 ( 
.A(n_514),
.B(n_431),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_468),
.B(n_411),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_534),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_475),
.B(n_326),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_469),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_495),
.Y(n_581)
);

NAND2x1_ASAP7_75t_SL g582 ( 
.A(n_520),
.B(n_327),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_472),
.B(n_329),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_475),
.B(n_329),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_468),
.B(n_434),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_489),
.B(n_333),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_480),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_514),
.B(n_329),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_500),
.Y(n_592)
);

NAND2x1p5_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_329),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_567),
.Y(n_594)
);

BUFx4_ASAP7_75t_SL g595 ( 
.A(n_587),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_542),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_575),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_507),
.Y(n_598)
);

CKINVDCx11_ASAP7_75t_R g599 ( 
.A(n_557),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_586),
.Y(n_600)
);

BUFx2_ASAP7_75t_SL g601 ( 
.A(n_563),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_591),
.Y(n_602)
);

BUFx2_ASAP7_75t_SL g603 ( 
.A(n_563),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_570),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_538),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_541),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_556),
.A2(n_512),
.B1(n_498),
.B2(n_482),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_547),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_549),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_540),
.Y(n_611)
);

CKINVDCx8_ASAP7_75t_R g612 ( 
.A(n_554),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_588),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_472),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_549),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_560),
.A2(n_512),
.B1(n_498),
.B2(n_482),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_577),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_568),
.Y(n_619)
);

CKINVDCx8_ASAP7_75t_R g620 ( 
.A(n_587),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_581),
.Y(n_621)
);

CKINVDCx6p67_ASAP7_75t_R g622 ( 
.A(n_587),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_573),
.A2(n_530),
.B1(n_512),
.B2(n_487),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_584),
.Y(n_624)
);

BUFx2_ASAP7_75t_SL g625 ( 
.A(n_544),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

BUFx4_ASAP7_75t_SL g627 ( 
.A(n_559),
.Y(n_627)
);

BUFx12f_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_576),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_544),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_570),
.B(n_472),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_574),
.B(n_477),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

INVx2_ASAP7_75t_R g634 ( 
.A(n_571),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_574),
.Y(n_635)
);

BUFx4f_ASAP7_75t_L g636 ( 
.A(n_548),
.Y(n_636)
);

INVx8_ASAP7_75t_L g637 ( 
.A(n_548),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_590),
.B(n_560),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_559),
.Y(n_639)
);

BUFx12f_ASAP7_75t_L g640 ( 
.A(n_550),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_551),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_637),
.Y(n_642)
);

CKINVDCx6p67_ASAP7_75t_R g643 ( 
.A(n_611),
.Y(n_643)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_637),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_612),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_638),
.A2(n_530),
.B1(n_546),
.B2(n_552),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_633),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_602),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_596),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_619),
.A2(n_589),
.B1(n_506),
.B2(n_480),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_598),
.B(n_578),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_617),
.A2(n_546),
.B1(n_552),
.B2(n_589),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_601),
.B(n_496),
.Y(n_654)
);

INVx6_ASAP7_75t_L g655 ( 
.A(n_613),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_637),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_600),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_595),
.Y(n_658)
);

BUFx8_ASAP7_75t_L g659 ( 
.A(n_611),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_619),
.A2(n_548),
.B1(n_550),
.B2(n_512),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_594),
.Y(n_662)
);

INVx6_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_623),
.A2(n_539),
.B1(n_561),
.B2(n_558),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_621),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_594),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_603),
.A2(n_512),
.B1(n_639),
.B2(n_628),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_624),
.B(n_545),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_635),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_609),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_623),
.A2(n_561),
.B(n_558),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_608),
.B(n_512),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_609),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_637),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_628),
.A2(n_512),
.B1(n_564),
.B2(n_548),
.Y(n_675)
);

BUFx12f_ASAP7_75t_L g676 ( 
.A(n_599),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_621),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_636),
.A2(n_539),
.B1(n_492),
.B2(n_481),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_624),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_605),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_614),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_599),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_636),
.B(n_574),
.Y(n_683)
);

INVx8_ASAP7_75t_L g684 ( 
.A(n_635),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_652),
.B(n_469),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_679),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_668),
.B(n_641),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_652),
.B(n_473),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_651),
.A2(n_506),
.B1(n_629),
.B2(n_639),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_647),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_660),
.A2(n_620),
.B1(n_629),
.B2(n_618),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_646),
.A2(n_506),
.B1(n_555),
.B2(n_512),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_681),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_654),
.B(n_487),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_660),
.A2(n_620),
.B1(n_618),
.B2(n_622),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_668),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_662),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_653),
.A2(n_622),
.B1(n_640),
.B2(n_473),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_665),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_653),
.A2(n_640),
.B1(n_517),
.B2(n_564),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_644),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_677),
.B(n_533),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_648),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_667),
.A2(n_517),
.B1(n_490),
.B2(n_536),
.Y(n_704)
);

BUFx4f_ASAP7_75t_SL g705 ( 
.A(n_676),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_645),
.A2(n_490),
.B1(n_512),
.B2(n_536),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_675),
.A2(n_533),
.B1(n_606),
.B2(n_607),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_669),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_SL g709 ( 
.A1(n_671),
.A2(n_501),
.B(n_511),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_672),
.A2(n_671),
.B1(n_649),
.B2(n_680),
.Y(n_710)
);

BUFx4f_ASAP7_75t_L g711 ( 
.A(n_643),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_664),
.A2(n_501),
.B1(n_634),
.B2(n_502),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_664),
.A2(n_634),
.B1(n_502),
.B2(n_499),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_650),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_672),
.A2(n_499),
.B1(n_592),
.B2(n_515),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_678),
.A2(n_484),
.B1(n_486),
.B2(n_515),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_644),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_657),
.B(n_504),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_678),
.A2(n_579),
.B1(n_585),
.B2(n_610),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_666),
.B(n_511),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_661),
.A2(n_484),
.B1(n_486),
.B2(n_585),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_670),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_673),
.A2(n_579),
.B1(n_531),
.B2(n_504),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_657),
.B(n_518),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_655),
.A2(n_531),
.B1(n_508),
.B2(n_504),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_642),
.B(n_626),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_659),
.A2(n_510),
.B1(n_500),
.B2(n_509),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_659),
.A2(n_510),
.B1(n_500),
.B2(n_509),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_656),
.A2(n_509),
.B1(n_529),
.B2(n_518),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_656),
.A2(n_529),
.B1(n_525),
.B2(n_527),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_655),
.B(n_519),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_683),
.A2(n_663),
.B1(n_642),
.B2(n_674),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_695),
.A2(n_682),
.B1(n_663),
.B2(n_644),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_689),
.A2(n_529),
.B1(n_519),
.B2(n_523),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_SL g736 ( 
.A1(n_689),
.A2(n_683),
.B(n_524),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_691),
.A2(n_524),
.B1(n_523),
.B2(n_525),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_688),
.B(n_508),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_698),
.A2(n_508),
.B1(n_528),
.B2(n_674),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_697),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_700),
.A2(n_627),
.B1(n_616),
.B2(n_610),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_694),
.B(n_669),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_SL g743 ( 
.A1(n_685),
.A2(n_610),
.B1(n_616),
.B2(n_625),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_706),
.A2(n_528),
.B1(n_505),
.B2(n_532),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_693),
.B(n_669),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_692),
.A2(n_528),
.B1(n_505),
.B2(n_532),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_692),
.A2(n_532),
.B1(n_485),
.B2(n_527),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_727),
.A2(n_543),
.B1(n_616),
.B2(n_604),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_710),
.A2(n_485),
.B1(n_526),
.B2(n_553),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_696),
.A2(n_485),
.B1(n_526),
.B2(n_684),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_727),
.A2(n_604),
.B1(n_615),
.B2(n_631),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_687),
.A2(n_485),
.B1(n_684),
.B2(n_470),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_704),
.A2(n_684),
.B1(n_604),
.B2(n_626),
.Y(n_753)
);

AOI221xp5_ASAP7_75t_L g754 ( 
.A1(n_709),
.A2(n_520),
.B1(n_477),
.B2(n_470),
.C(n_630),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_728),
.A2(n_631),
.B1(n_615),
.B2(n_630),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_687),
.A2(n_730),
.B1(n_728),
.B2(n_716),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_712),
.A2(n_470),
.B1(n_630),
.B2(n_626),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_721),
.A2(n_470),
.B1(n_477),
.B2(n_569),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_724),
.A2(n_477),
.B1(n_572),
.B2(n_569),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_690),
.B(n_582),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_703),
.B(n_635),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_719),
.A2(n_712),
.B1(n_713),
.B2(n_705),
.Y(n_762)
);

OAI221xp5_ASAP7_75t_L g763 ( 
.A1(n_732),
.A2(n_583),
.B1(n_565),
.B2(n_593),
.C(n_632),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_713),
.A2(n_635),
.B1(n_572),
.B2(n_477),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_705),
.A2(n_477),
.B1(n_593),
.B2(n_343),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_SL g766 ( 
.A(n_699),
.B(n_632),
.C(n_494),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_686),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_714),
.A2(n_343),
.B1(n_33),
.B2(n_34),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_702),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_733),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_770)
);

OAI222xp33_ASAP7_75t_L g771 ( 
.A1(n_707),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.C1(n_49),
.C2(n_50),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_738),
.B(n_722),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_740),
.B(n_715),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_760),
.B(n_718),
.C(n_701),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_742),
.B(n_715),
.Y(n_775)
);

OAI221xp5_ASAP7_75t_SL g776 ( 
.A1(n_736),
.A2(n_731),
.B1(n_725),
.B2(n_723),
.C(n_729),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_762),
.A2(n_731),
.B(n_729),
.Y(n_777)
);

OAI221xp5_ASAP7_75t_SL g778 ( 
.A1(n_756),
.A2(n_720),
.B1(n_708),
.B2(n_717),
.C(n_701),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_734),
.A2(n_711),
.B1(n_726),
.B2(n_717),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_735),
.B(n_726),
.C(n_711),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_767),
.B(n_51),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_745),
.B(n_54),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_761),
.B(n_56),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_741),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_743),
.B(n_64),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_753),
.B(n_65),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_754),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_71),
.Y(n_788)
);

OA21x2_ASAP7_75t_L g789 ( 
.A1(n_749),
.A2(n_764),
.B(n_757),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_SL g790 ( 
.A1(n_771),
.A2(n_72),
.B(n_73),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_757),
.B(n_735),
.Y(n_791)
);

AOI21xp33_ASAP7_75t_L g792 ( 
.A1(n_768),
.A2(n_74),
.B(n_75),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_764),
.B(n_79),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_758),
.B(n_81),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_746),
.B(n_82),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_770),
.B(n_83),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_737),
.B(n_84),
.C(n_87),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_763),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_747),
.B(n_88),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_737),
.B(n_90),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_775),
.B(n_759),
.Y(n_801)
);

OAI211xp5_ASAP7_75t_SL g802 ( 
.A1(n_774),
.A2(n_752),
.B(n_750),
.C(n_739),
.Y(n_802)
);

AOI211xp5_ASAP7_75t_L g803 ( 
.A1(n_790),
.A2(n_769),
.B(n_766),
.C(n_751),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_790),
.B(n_748),
.C(n_755),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_798),
.B(n_778),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_772),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_798),
.B(n_765),
.C(n_93),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_780),
.B(n_91),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_772),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_797),
.A2(n_94),
.B1(n_99),
.B2(n_100),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_775),
.B(n_102),
.Y(n_811)
);

AND2x2_ASAP7_75t_SL g812 ( 
.A(n_793),
.B(n_103),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_780),
.B(n_104),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_773),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_792),
.B(n_106),
.C(n_107),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_783),
.B(n_108),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_783),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_792),
.B(n_109),
.C(n_110),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_813),
.B(n_797),
.C(n_796),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_806),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_805),
.B(n_776),
.C(n_800),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_806),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_817),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_814),
.B(n_789),
.Y(n_824)
);

XNOR2xp5_ASAP7_75t_L g825 ( 
.A(n_812),
.B(n_779),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_812),
.Y(n_826)
);

NAND4xp75_ASAP7_75t_SL g827 ( 
.A(n_808),
.B(n_786),
.C(n_789),
.D(n_793),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_809),
.Y(n_828)
);

XOR2x2_ASAP7_75t_L g829 ( 
.A(n_825),
.B(n_805),
.Y(n_829)
);

XNOR2x1_ASAP7_75t_L g830 ( 
.A(n_821),
.B(n_811),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_820),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_828),
.Y(n_832)
);

XNOR2x1_ASAP7_75t_L g833 ( 
.A(n_821),
.B(n_801),
.Y(n_833)
);

OAI22x1_ASAP7_75t_L g834 ( 
.A1(n_832),
.A2(n_826),
.B1(n_823),
.B2(n_813),
.Y(n_834)
);

XNOR2xp5_ASAP7_75t_L g835 ( 
.A(n_829),
.B(n_827),
.Y(n_835)
);

XOR2x2_ASAP7_75t_L g836 ( 
.A(n_833),
.B(n_826),
.Y(n_836)
);

XOR2x2_ASAP7_75t_L g837 ( 
.A(n_830),
.B(n_819),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_831),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_836),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_838),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_837),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_834),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_840),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_842),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_841),
.A2(n_835),
.B1(n_804),
.B2(n_808),
.Y(n_845)
);

AOI221xp5_ASAP7_75t_L g846 ( 
.A1(n_844),
.A2(n_839),
.B1(n_843),
.B2(n_835),
.C(n_845),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_844),
.Y(n_847)
);

AOI22x1_ASAP7_75t_SL g848 ( 
.A1(n_844),
.A2(n_831),
.B1(n_822),
.B2(n_803),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_844),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_846),
.A2(n_824),
.B1(n_815),
.B2(n_818),
.Y(n_850)
);

AO22x2_ASAP7_75t_L g851 ( 
.A1(n_848),
.A2(n_807),
.B1(n_781),
.B2(n_786),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_847),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_849),
.A2(n_816),
.B1(n_810),
.B2(n_802),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_846),
.A2(n_777),
.B1(n_788),
.B2(n_782),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_846),
.A2(n_777),
.B1(n_788),
.B2(n_785),
.Y(n_855)
);

NOR2x1_ASAP7_75t_L g856 ( 
.A(n_847),
.B(n_794),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_852),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_856),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_853),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_851),
.A2(n_784),
.B1(n_795),
.B2(n_799),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_854),
.B(n_794),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_855),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_850),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_852),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_860),
.A2(n_787),
.B1(n_791),
.B2(n_795),
.Y(n_865)
);

AO22x2_ASAP7_75t_L g866 ( 
.A1(n_858),
.A2(n_799),
.B1(n_118),
.B2(n_120),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_857),
.Y(n_867)
);

NAND4xp25_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_113),
.C(n_121),
.D(n_123),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_863),
.A2(n_789),
.B1(n_126),
.B2(n_127),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_SL g870 ( 
.A(n_859),
.B(n_124),
.C(n_129),
.Y(n_870)
);

OAI211xp5_ASAP7_75t_L g871 ( 
.A1(n_864),
.A2(n_789),
.B(n_134),
.C(n_135),
.Y(n_871)
);

AO22x2_ASAP7_75t_L g872 ( 
.A1(n_861),
.A2(n_860),
.B1(n_137),
.B2(n_138),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_867),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_872),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_866),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_869),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_865),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_870),
.A2(n_131),
.B1(n_140),
.B2(n_141),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_871),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_879)
);

AO22x2_ASAP7_75t_L g880 ( 
.A1(n_874),
.A2(n_868),
.B1(n_147),
.B2(n_148),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_875),
.Y(n_881)
);

OAI22x1_ASAP7_75t_L g882 ( 
.A1(n_877),
.A2(n_146),
.B1(n_150),
.B2(n_154),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_873),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_878),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_876),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_879),
.A2(n_162),
.B1(n_167),
.B2(n_169),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_881),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_883),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_882),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_880),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_887),
.A2(n_880),
.B1(n_886),
.B2(n_884),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_889),
.A2(n_885),
.B1(n_172),
.B2(n_173),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_891),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_892),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_893),
.A2(n_890),
.B1(n_888),
.B2(n_175),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_895),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_896),
.A2(n_894),
.B1(n_174),
.B2(n_176),
.C(n_178),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_897),
.A2(n_171),
.B1(n_182),
.B2(n_183),
.Y(n_898)
);


endmodule