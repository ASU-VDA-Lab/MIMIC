module real_jpeg_1509_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_70),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_38),
.B1(n_48),
.B2(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_38),
.B1(n_65),
.B2(n_66),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_5),
.A2(n_50),
.B1(n_65),
.B2(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_50),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_23),
.C(n_45),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_6),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_25),
.B1(n_48),
.B2(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_6),
.A2(n_25),
.B1(n_65),
.B2(n_66),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_43),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_6),
.B(n_29),
.C(n_31),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_66),
.C(n_84),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_27),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_6),
.B(n_63),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_88),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_130),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_129),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_107),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_16),
.B(n_107),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.C(n_90),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_17),
.B(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_57),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_41),
.B2(n_56),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_56),
.C(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_22),
.A2(n_27),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_22),
.B(n_117),
.Y(n_182)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_23),
.A2(n_26),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_23),
.B(n_162),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_27),
.B(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_28),
.B(n_104),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_30),
.A2(n_31),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_31),
.B(n_191),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_35),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_39),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_47),
.B(n_53),
.Y(n_115)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B(n_71),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_73),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_62),
.A2(n_72),
.B(n_128),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_62),
.B(n_197),
.Y(n_211)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_63),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_72),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_66),
.B1(n_83),
.B2(n_84),
.Y(n_86)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_66),
.B(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_71),
.B(n_210),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_72),
.B(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_90),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_77),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_79),
.B(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_80),
.B(n_88),
.Y(n_166)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_81),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_87),
.B(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_88),
.B(n_168),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_102),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI21x1_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_120),
.B2(n_121),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_126),
.B(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_150),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_148),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_148),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_140),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_135),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_140),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_147),
.B(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_172),
.B(n_229),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_169),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_154),
.B(n_169),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.C(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_156),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_164),
.B1(n_165),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21x1_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_185),
.B(n_228),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_181),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_226),
.Y(n_225)
);

OAI21x1_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_223),
.B(n_227),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_205),
.B(n_222),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_198),
.B1(n_199),
.B2(n_204),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_202),
.C(n_204),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_212),
.B(n_221),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_209),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B(n_220),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_225),
.Y(n_227)
);


endmodule