module real_aes_15855_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g877 ( .A(n_0), .B(n_878), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_1), .A2(n_86), .B1(n_855), .B2(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g856 ( .A(n_1), .Y(n_856) );
AOI22x1_ASAP7_75t_SL g127 ( .A1(n_2), .A2(n_128), .B1(n_129), .B2(n_135), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_2), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_3), .A2(n_6), .B1(n_257), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_4), .A2(n_46), .B1(n_152), .B2(n_154), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_5), .A2(n_26), .B1(n_154), .B2(n_197), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_7), .A2(n_18), .B1(n_179), .B2(n_248), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_8), .A2(n_64), .B1(n_199), .B2(n_224), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_9), .A2(n_19), .B1(n_152), .B2(n_183), .Y(n_614) );
INVx1_ASAP7_75t_L g878 ( .A(n_10), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_11), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_12), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_13), .A2(n_20), .B1(n_181), .B2(n_223), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_14), .A2(n_90), .B1(n_852), .B2(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_14), .Y(n_852) );
OR2x2_ASAP7_75t_L g115 ( .A(n_15), .B(n_41), .Y(n_115) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_16), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_17), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_21), .A2(n_101), .B1(n_179), .B2(n_257), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_22), .A2(n_42), .B1(n_215), .B2(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_23), .B(n_180), .Y(n_212) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_24), .A2(n_61), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_25), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_27), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_28), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_29), .B(n_158), .Y(n_522) );
INVx4_ASAP7_75t_R g577 ( .A(n_30), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_31), .A2(n_51), .B1(n_160), .B2(n_162), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_32), .A2(n_105), .B1(n_873), .B2(n_879), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_33), .A2(n_57), .B1(n_162), .B2(n_179), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_34), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_35), .B(n_215), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_36), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_37), .B(n_154), .Y(n_529) );
INVx1_ASAP7_75t_L g538 ( .A(n_38), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_SL g595 ( .A1(n_39), .A2(n_152), .B(n_164), .C(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_40), .A2(n_58), .B1(n_152), .B2(n_162), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_43), .A2(n_88), .B1(n_152), .B2(n_196), .Y(n_195) );
AOI22x1_ASAP7_75t_SL g131 ( .A1(n_44), .A2(n_59), .B1(n_132), .B2(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_44), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_45), .A2(n_50), .B1(n_152), .B2(n_183), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_47), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_48), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_49), .A2(n_63), .B1(n_179), .B2(n_234), .Y(n_259) );
INVx1_ASAP7_75t_L g526 ( .A(n_52), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_53), .B(n_152), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_54), .Y(n_547) );
INVx2_ASAP7_75t_L g121 ( .A(n_55), .Y(n_121) );
INVx1_ASAP7_75t_L g113 ( .A(n_56), .Y(n_113) );
BUFx3_ASAP7_75t_L g124 ( .A(n_56), .Y(n_124) );
INVx1_ASAP7_75t_L g133 ( .A(n_59), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_60), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_62), .A2(n_89), .B1(n_152), .B2(n_162), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_65), .A2(n_77), .B1(n_160), .B2(n_234), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_66), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_67), .A2(n_79), .B1(n_152), .B2(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_68), .A2(n_99), .B1(n_179), .B2(n_181), .Y(n_178) );
AND2x4_ASAP7_75t_L g148 ( .A(n_69), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g169 ( .A(n_70), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_71), .A2(n_92), .B1(n_160), .B2(n_162), .Y(n_534) );
AO22x1_ASAP7_75t_L g564 ( .A1(n_72), .A2(n_78), .B1(n_245), .B2(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g149 ( .A(n_73), .Y(n_149) );
AND2x2_ASAP7_75t_L g598 ( .A(n_74), .B(n_166), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_75), .B(n_199), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_76), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_80), .B(n_154), .Y(n_548) );
INVx2_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_82), .B(n_166), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_83), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_84), .A2(n_100), .B1(n_162), .B2(n_199), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_85), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_86), .B(n_176), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_86), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_87), .Y(n_171) );
INVx1_ASAP7_75t_L g853 ( .A(n_90), .Y(n_853) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_91), .B(n_166), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_93), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_94), .B(n_166), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_95), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g497 ( .A(n_95), .Y(n_497) );
NAND2xp33_ASAP7_75t_L g216 ( .A(n_96), .B(n_180), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_97), .A2(n_185), .B(n_199), .C(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_98), .B(n_580), .Y(n_579) );
NAND2xp33_ASAP7_75t_L g552 ( .A(n_102), .B(n_161), .Y(n_552) );
OAI22x1_ASAP7_75t_L g129 ( .A1(n_103), .A2(n_130), .B1(n_131), .B2(n_134), .Y(n_129) );
INVxp67_ASAP7_75t_SL g134 ( .A(n_103), .Y(n_134) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_116), .Y(n_105) );
INVx1_ASAP7_75t_L g860 ( .A(n_106), .Y(n_860) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
BUFx12f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g848 ( .A(n_110), .Y(n_848) );
AND2x6_ASAP7_75t_SL g110 ( .A(n_111), .B(n_114), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_114), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NOR2x1_ASAP7_75t_L g872 ( .A(n_115), .B(n_124), .Y(n_872) );
OAI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_125), .B(n_844), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g864 ( .A(n_121), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_121), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_136), .B2(n_843), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g843 ( .A(n_136), .Y(n_843) );
OA22x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_493), .B1(n_498), .B2(n_500), .Y(n_136) );
INVx2_ASAP7_75t_L g858 ( .A(n_137), .Y(n_858) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_137), .B(n_847), .C(n_850), .Y(n_859) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_389), .Y(n_137) );
NOR2x1_ASAP7_75t_L g138 ( .A(n_139), .B(n_341), .Y(n_138) );
NAND3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_288), .C(n_326), .Y(n_139) );
AOI221xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_219), .B1(n_239), .B2(n_267), .C(n_273), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_141), .A2(n_466), .B1(n_469), .B2(n_470), .Y(n_465) );
INVx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_190), .Y(n_142) );
INVx1_ASAP7_75t_L g380 ( .A(n_143), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_172), .Y(n_143) );
INVx1_ASAP7_75t_L g332 ( .A(n_144), .Y(n_332) );
AND2x4_ASAP7_75t_L g375 ( .A(n_144), .B(n_296), .Y(n_375) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g303 ( .A(n_145), .B(n_206), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_145), .B(n_272), .Y(n_363) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g271 ( .A(n_146), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g287 ( .A(n_146), .B(n_192), .Y(n_287) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_146), .Y(n_294) );
INVx1_ASAP7_75t_L g350 ( .A(n_146), .Y(n_350) );
AO31x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .A3(n_165), .B(n_170), .Y(n_146) );
INVx2_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
AO31x2_ASAP7_75t_L g220 ( .A1(n_147), .A2(n_174), .A3(n_221), .B(n_227), .Y(n_220) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_147), .A2(n_193), .A3(n_243), .B(n_250), .Y(n_242) );
AO31x2_ASAP7_75t_L g612 ( .A1(n_147), .A2(n_238), .A3(n_613), .B(n_616), .Y(n_612) );
BUFx10_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
BUFx10_ASAP7_75t_L g513 ( .A(n_148), .Y(n_513) );
INVx1_ASAP7_75t_L g568 ( .A(n_148), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B1(n_159), .B2(n_163), .Y(n_150) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx4_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx1_ASAP7_75t_L g234 ( .A(n_152), .Y(n_234) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_153), .Y(n_154) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
INVx2_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
INVx1_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
INVx1_ASAP7_75t_L g225 ( .A(n_153), .Y(n_225) );
INVx1_ASAP7_75t_L g246 ( .A(n_153), .Y(n_246) );
INVx1_ASAP7_75t_L g249 ( .A(n_153), .Y(n_249) );
INVx1_ASAP7_75t_L g258 ( .A(n_153), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_154), .B(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_155), .A2(n_163), .B1(n_233), .B2(n_235), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_155), .A2(n_163), .B1(n_244), .B2(n_247), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_155), .A2(n_163), .B1(n_256), .B2(n_259), .Y(n_255) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g512 ( .A(n_156), .Y(n_512) );
BUFx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g550 ( .A(n_157), .Y(n_550) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx8_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
INVx1_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
INVx1_ASAP7_75t_L g525 ( .A(n_158), .Y(n_525) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_161), .A2(n_249), .B1(n_577), .B2(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_162), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g536 ( .A(n_162), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_163), .A2(n_178), .B1(n_182), .B2(n_184), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_163), .A2(n_195), .B1(n_198), .B2(n_200), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_163), .A2(n_214), .B(n_216), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_163), .A2(n_184), .B1(n_222), .B2(n_226), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_163), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_163), .A2(n_200), .B1(n_534), .B2(n_535), .Y(n_533) );
OAI22x1_ASAP7_75t_L g613 ( .A1(n_163), .A2(n_200), .B1(n_614), .B2(n_615), .Y(n_613) );
INVx6_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g210 ( .A1(n_164), .A2(n_183), .B(n_211), .C(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_164), .A2(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_164), .B(n_564), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_164), .A2(n_560), .B(n_564), .C(n_567), .Y(n_626) );
AO31x2_ASAP7_75t_L g508 ( .A1(n_165), .A2(n_509), .A3(n_513), .B(n_514), .Y(n_508) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_166), .B(n_555), .Y(n_554) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_167), .B(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_167), .B(n_189), .Y(n_188) );
BUFx3_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
INVx2_ASAP7_75t_SL g208 ( .A(n_167), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_167), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g530 ( .A(n_167), .B(n_513), .Y(n_530) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g176 ( .A(n_168), .Y(n_176) );
INVx3_ASAP7_75t_L g270 ( .A(n_172), .Y(n_270) );
AND2x2_ASAP7_75t_L g285 ( .A(n_172), .B(n_206), .Y(n_285) );
INVx2_ASAP7_75t_L g291 ( .A(n_172), .Y(n_291) );
AND2x4_ASAP7_75t_L g353 ( .A(n_172), .B(n_192), .Y(n_353) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_172), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_172), .B(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g302 ( .A(n_173), .B(n_192), .Y(n_302) );
AND2x2_ASAP7_75t_L g330 ( .A(n_173), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g409 ( .A(n_173), .Y(n_409) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .A3(n_186), .B(n_188), .Y(n_173) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_174), .A2(n_201), .A3(n_533), .B(n_537), .Y(n_532) );
AOI21x1_ASAP7_75t_L g587 ( .A1(n_174), .A2(n_588), .B(n_598), .Y(n_587) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_175), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_175), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g580 ( .A(n_175), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_175), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g204 ( .A(n_176), .Y(n_204) );
INVx2_ASAP7_75t_L g238 ( .A(n_176), .Y(n_238) );
OAI21xp33_ASAP7_75t_L g567 ( .A1(n_176), .A2(n_562), .B(n_568), .Y(n_567) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVxp67_ASAP7_75t_SL g565 ( .A(n_180), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_183), .A2(n_547), .B(n_548), .C(n_549), .Y(n_546) );
INVx1_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g200 ( .A(n_185), .Y(n_200) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_230), .A3(n_255), .B(n_260), .Y(n_254) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_187), .A2(n_572), .B(n_575), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_206), .Y(n_190) );
INVx1_ASAP7_75t_L g365 ( .A(n_191), .Y(n_365) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_191), .B(n_285), .Y(n_393) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g295 ( .A(n_192), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g331 ( .A(n_192), .Y(n_331) );
INVx1_ASAP7_75t_L g407 ( .A(n_192), .Y(n_407) );
AO31x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .A3(n_201), .B(n_203), .Y(n_192) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_197), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_200), .B(n_576), .Y(n_575) );
AO31x2_ASAP7_75t_L g229 ( .A1(n_201), .A2(n_230), .A3(n_232), .B(n_236), .Y(n_229) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_SL g217 ( .A(n_202), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_SL g227 ( .A(n_204), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g231 ( .A(n_204), .Y(n_231) );
AND2x4_ASAP7_75t_L g346 ( .A(n_206), .B(n_331), .Y(n_346) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g368 ( .A(n_207), .Y(n_368) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_218), .Y(n_207) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_208), .A2(n_209), .B(n_218), .Y(n_272) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_213), .B(n_217), .Y(n_209) );
AND2x4_ASAP7_75t_L g240 ( .A(n_219), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
INVx4_ASAP7_75t_SL g264 ( .A(n_220), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_220), .B(n_266), .Y(n_276) );
BUFx2_ASAP7_75t_L g340 ( .A(n_220), .Y(n_340) );
AND2x2_ASAP7_75t_L g384 ( .A(n_220), .B(n_242), .Y(n_384) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_225), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
OR2x2_ASAP7_75t_L g300 ( .A(n_229), .B(n_242), .Y(n_300) );
INVx2_ASAP7_75t_L g311 ( .A(n_229), .Y(n_311) );
AND2x4_ASAP7_75t_L g314 ( .A(n_229), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_229), .Y(n_355) );
INVx1_ASAP7_75t_L g396 ( .A(n_229), .Y(n_396) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_230), .A2(n_571), .B(n_579), .Y(n_570) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_238), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_252), .Y(n_239) );
INVx2_ASAP7_75t_L g489 ( .A(n_240), .Y(n_489) );
AND2x4_ASAP7_75t_L g450 ( .A(n_241), .B(n_253), .Y(n_450) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
INVx2_ASAP7_75t_L g315 ( .A(n_242), .Y(n_315) );
INVx1_ASAP7_75t_L g371 ( .A(n_242), .Y(n_371) );
AND2x2_ASAP7_75t_L g397 ( .A(n_242), .B(n_322), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_242), .B(n_310), .Y(n_401) );
OAI21xp33_ASAP7_75t_SL g521 ( .A1(n_245), .A2(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_263), .Y(n_252) );
INVx3_ASAP7_75t_L g378 ( .A(n_253), .Y(n_378) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_262), .Y(n_253) );
INVx2_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
INVx2_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_258), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_262), .B(n_264), .Y(n_323) );
AND2x2_ASAP7_75t_L g351 ( .A(n_262), .B(n_322), .Y(n_351) );
INVx1_ASAP7_75t_L g277 ( .A(n_263), .Y(n_277) );
NAND2x1_ASAP7_75t_L g413 ( .A(n_263), .B(n_387), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_263), .B(n_351), .Y(n_462) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g280 ( .A(n_264), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_264), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g370 ( .A(n_264), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_264), .Y(n_447) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_267), .A2(n_460), .B1(n_461), .B2(n_463), .Y(n_459) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_269), .B(n_303), .Y(n_338) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g361 ( .A(n_270), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g460 ( .A(n_270), .B(n_271), .Y(n_460) );
AND2x2_ASAP7_75t_L g333 ( .A(n_271), .B(n_302), .Y(n_333) );
AND2x4_ASAP7_75t_L g352 ( .A(n_271), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g403 ( .A(n_271), .B(n_330), .Y(n_403) );
INVx1_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
AOI31xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .A3(n_278), .B(n_283), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_275), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_275), .Y(n_469) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_275), .A2(n_277), .B(n_307), .Y(n_487) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g464 ( .A(n_279), .B(n_300), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
INVx1_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_281), .Y(n_426) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
OR2x2_ASAP7_75t_L g336 ( .A(n_282), .B(n_311), .Y(n_336) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2x1p5_ASAP7_75t_L g325 ( .A(n_287), .B(n_291), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_297), .B1(n_301), .B2(n_304), .C(n_316), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2x1_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g405 ( .A(n_294), .B(n_308), .Y(n_405) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g335 ( .A(n_298), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g422 ( .A(n_298), .B(n_314), .Y(n_422) );
AND2x4_ASAP7_75t_L g339 ( .A(n_299), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g358 ( .A(n_300), .B(n_321), .Y(n_358) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x4_ASAP7_75t_SL g374 ( .A(n_302), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g415 ( .A(n_302), .Y(n_415) );
INVx2_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
AND2x2_ASAP7_75t_L g438 ( .A(n_302), .B(n_368), .Y(n_438) );
INVx1_ASAP7_75t_L g416 ( .A(n_303), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_312), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_306), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_307), .B(n_314), .Y(n_348) );
AND2x2_ASAP7_75t_L g369 ( .A(n_307), .B(n_370), .Y(n_369) );
NAND2x1_ASAP7_75t_L g477 ( .A(n_307), .B(n_339), .Y(n_477) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B(n_324), .Y(n_316) );
NAND2x1_ASAP7_75t_L g478 ( .A(n_318), .B(n_422), .Y(n_478) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_319), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx4_ASAP7_75t_L g387 ( .A(n_321), .Y(n_387) );
AND2x2_ASAP7_75t_L g457 ( .A(n_321), .B(n_362), .Y(n_457) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g354 ( .A(n_322), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g367 ( .A(n_325), .B(n_368), .Y(n_367) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_325), .B(n_438), .Y(n_437) );
AOI322xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .A3(n_332), .B1(n_333), .B2(n_334), .C1(n_337), .C2(n_339), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g420 ( .A(n_330), .B(n_368), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_330), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g444 ( .A(n_330), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g449 ( .A(n_330), .B(n_434), .Y(n_449) );
INVx1_ASAP7_75t_L g458 ( .A(n_330), .Y(n_458) );
OR2x2_ASAP7_75t_L g344 ( .A(n_332), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g471 ( .A(n_332), .Y(n_471) );
AND2x2_ASAP7_75t_L g474 ( .A(n_333), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_336), .B(n_350), .C(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g452 ( .A(n_336), .Y(n_452) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND3xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_356), .C(n_366), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_349), .B2(n_351), .C1(n_352), .C2(n_354), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI22x1_ASAP7_75t_L g488 ( .A1(n_345), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g349 ( .A(n_346), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_346), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g442 ( .A(n_346), .B(n_408), .Y(n_442) );
AND2x4_ASAP7_75t_L g472 ( .A(n_346), .B(n_409), .Y(n_472) );
AND2x2_ASAP7_75t_L g453 ( .A(n_347), .B(n_420), .Y(n_453) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g445 ( .A(n_350), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_351), .B(n_384), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_351), .B(n_370), .Y(n_468) );
INVx1_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
INVx2_ASAP7_75t_L g432 ( .A(n_354), .Y(n_432) );
INVx1_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .Y(n_360) );
AOI221xp5_ASAP7_75t_SL g448 ( .A1(n_361), .A2(n_449), .B1(n_450), .B2(n_451), .C(n_453), .Y(n_448) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g434 ( .A(n_363), .Y(n_434) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_363), .Y(n_486) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_365), .B(n_471), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_372), .B2(n_383), .C(n_385), .Y(n_366) );
OR2x2_ASAP7_75t_L g423 ( .A(n_368), .B(n_424), .Y(n_423) );
AOI32xp33_ASAP7_75t_L g404 ( .A1(n_370), .A2(n_384), .A3(n_405), .B1(n_406), .B2(n_410), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_370), .B(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B1(n_379), .B2(n_381), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_375), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g446 ( .A(n_378), .B(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g439 ( .A(n_382), .B(n_384), .Y(n_439) );
AND2x2_ASAP7_75t_L g492 ( .A(n_382), .B(n_397), .Y(n_492) );
AND2x2_ASAP7_75t_L g451 ( .A(n_383), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_384), .B(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_454), .Y(n_389) );
NAND4xp75_ASAP7_75t_L g390 ( .A(n_391), .B(n_417), .C(n_435), .D(n_448), .Y(n_390) );
AOI211x1_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_398), .C(n_412), .Y(n_391) );
INVxp67_ASAP7_75t_L g490 ( .A(n_392), .Y(n_490) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
BUFx2_ASAP7_75t_L g411 ( .A(n_407), .Y(n_411) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g483 ( .A(n_411), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .C(n_416), .Y(n_412) );
INVx2_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_427), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_423), .B2(n_425), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_432), .B2(n_433), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_440), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_447), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
NAND4xp75_ASAP7_75t_SL g454 ( .A(n_455), .B(n_465), .C(n_473), .D(n_481), .Y(n_454) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
NOR2xp67_ASAP7_75t_SL g473 ( .A(n_474), .B(n_476), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_479), .Y(n_476) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
AOI21x1_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_487), .B(n_488), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx8_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx12f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
BUFx8_ASAP7_75t_SL g499 ( .A(n_496), .Y(n_499) );
AND2x2_ASAP7_75t_L g871 ( .A(n_496), .B(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_733), .Y(n_500) );
NOR4xp25_ASAP7_75t_L g501 ( .A(n_502), .B(n_633), .C(n_675), .D(n_707), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_539), .B(n_581), .C(n_618), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_516), .Y(n_505) );
INVx2_ASAP7_75t_L g646 ( .A(n_506), .Y(n_646) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g725 ( .A(n_507), .B(n_518), .Y(n_725) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_508), .B(n_532), .Y(n_584) );
AND2x2_ASAP7_75t_L g607 ( .A(n_508), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_SL g632 ( .A(n_508), .Y(n_632) );
OR2x2_ASAP7_75t_L g695 ( .A(n_508), .B(n_532), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_512), .A2(n_528), .B(n_529), .Y(n_527) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_512), .A2(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g555 ( .A(n_513), .Y(n_555) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g629 ( .A(n_517), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g641 ( .A(n_517), .Y(n_641) );
INVxp67_ASAP7_75t_SL g819 ( .A(n_517), .Y(n_819) );
OR2x2_ASAP7_75t_L g832 ( .A(n_517), .B(n_833), .Y(n_832) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_531), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_518), .B(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g605 ( .A(n_518), .Y(n_605) );
AND2x2_ASAP7_75t_L g652 ( .A(n_518), .B(n_653), .Y(n_652) );
NAND2x1p5_ASAP7_75t_SL g671 ( .A(n_518), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_518), .B(n_606), .Y(n_721) );
INVx1_ASAP7_75t_L g810 ( .A(n_518), .Y(n_810) );
AND2x2_ASAP7_75t_L g839 ( .A(n_518), .B(n_532), .Y(n_839) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_527), .B(n_530), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
BUFx4f_ASAP7_75t_L g594 ( .A(n_525), .Y(n_594) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g606 ( .A(n_532), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_532), .B(n_632), .Y(n_654) );
INVx1_ASAP7_75t_L g674 ( .A(n_532), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_532), .B(n_608), .Y(n_726) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_556), .Y(n_540) );
OR2x2_ASAP7_75t_L g623 ( .A(n_541), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g730 ( .A(n_541), .B(n_679), .Y(n_730) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g639 ( .A(n_542), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_542), .B(n_659), .Y(n_658) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_542), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g602 ( .A(n_543), .Y(n_602) );
BUFx3_ASAP7_75t_L g650 ( .A(n_543), .Y(n_650) );
AND2x2_ASAP7_75t_L g686 ( .A(n_543), .B(n_667), .Y(n_686) );
AND2x2_ASAP7_75t_L g766 ( .A(n_543), .B(n_612), .Y(n_766) );
AND2x2_ASAP7_75t_L g779 ( .A(n_543), .B(n_570), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_551), .B(n_554), .Y(n_545) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g719 ( .A(n_556), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_556), .B(n_649), .Y(n_727) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_569), .Y(n_556) );
AND2x2_ASAP7_75t_L g638 ( .A(n_557), .B(n_570), .Y(n_638) );
INVx1_ASAP7_75t_L g746 ( .A(n_557), .Y(n_746) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g600 ( .A(n_558), .B(n_570), .Y(n_600) );
AND2x2_ASAP7_75t_L g663 ( .A(n_558), .B(n_569), .Y(n_663) );
AOI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_563), .B(n_566), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_568), .A2(n_589), .B(n_595), .Y(n_588) );
AND2x2_ASAP7_75t_L g621 ( .A(n_569), .B(n_612), .Y(n_621) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g611 ( .A(n_570), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g679 ( .A(n_570), .B(n_612), .Y(n_679) );
INVx1_ASAP7_75t_L g690 ( .A(n_570), .Y(n_690) );
AND2x2_ASAP7_75t_L g753 ( .A(n_570), .B(n_602), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_599), .B1(n_603), .B2(n_609), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_582), .A2(n_652), .B1(n_655), .B2(n_657), .Y(n_651) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OR2x2_ASAP7_75t_L g731 ( .A(n_584), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g837 ( .A(n_584), .Y(n_837) );
INVx1_ASAP7_75t_L g696 ( .A(n_585), .Y(n_696) );
OR2x2_ASAP7_75t_L g759 ( .A(n_585), .B(n_654), .Y(n_759) );
OR2x2_ASAP7_75t_L g630 ( .A(n_586), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_586), .B(n_605), .Y(n_706) );
AND2x2_ASAP7_75t_L g723 ( .A(n_586), .B(n_650), .Y(n_723) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_586), .Y(n_740) );
INVxp67_ASAP7_75t_L g788 ( .A(n_586), .Y(n_788) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g608 ( .A(n_587), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_594), .Y(n_589) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_600), .Y(n_698) );
INVx3_ASAP7_75t_L g703 ( .A(n_600), .Y(n_703) );
AND2x2_ASAP7_75t_L g716 ( .A(n_600), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g816 ( .A(n_600), .B(n_778), .Y(n_816) );
INVx1_ASAP7_75t_L g610 ( .A(n_601), .Y(n_610) );
OR2x2_ASAP7_75t_L g793 ( .A(n_601), .B(n_768), .Y(n_793) );
BUFx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g717 ( .A(n_602), .B(n_627), .Y(n_717) );
AND2x2_ASAP7_75t_L g738 ( .A(n_602), .B(n_663), .Y(n_738) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_604), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g739 ( .A(n_604), .Y(n_739) );
AND2x2_ASAP7_75t_L g781 ( .A(n_604), .B(n_782), .Y(n_781) );
AND2x4_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx2_ASAP7_75t_L g682 ( .A(n_605), .Y(n_682) );
AND2x2_ASAP7_75t_L g713 ( .A(n_605), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_605), .B(n_672), .Y(n_732) );
AND2x2_ASAP7_75t_L g681 ( .A(n_607), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g797 ( .A(n_607), .Y(n_797) );
AND2x2_ASAP7_75t_L g820 ( .A(n_607), .B(n_810), .Y(n_820) );
INVx1_ASAP7_75t_L g833 ( .A(n_607), .Y(n_833) );
INVx2_ASAP7_75t_L g672 ( .A(n_608), .Y(n_672) );
OR2x2_ASAP7_75t_L g768 ( .A(n_608), .B(n_632), .Y(n_768) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_611), .B(n_649), .Y(n_656) );
INVx2_ASAP7_75t_L g627 ( .A(n_612), .Y(n_627) );
INVx2_ASAP7_75t_L g667 ( .A(n_612), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_612), .B(n_625), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_628), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_621), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g762 ( .A(n_624), .B(n_763), .Y(n_762) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g668 ( .A(n_625), .Y(n_668) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g659 ( .A(n_627), .Y(n_659) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g642 ( .A(n_630), .Y(n_642) );
INVxp67_ASAP7_75t_L g813 ( .A(n_630), .Y(n_813) );
OR2x2_ASAP7_75t_L g715 ( .A(n_631), .B(n_672), .Y(n_715) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_634), .B(n_643), .C(n_651), .D(n_660), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_640), .C(n_642), .Y(n_634) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g829 ( .A1(n_636), .A2(n_830), .B(n_832), .C(n_834), .Y(n_829) );
OR2x6_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_638), .B(n_686), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_638), .B(n_742), .C(n_744), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_638), .B(n_717), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_638), .A2(n_743), .B1(n_835), .B2(n_838), .C(n_840), .Y(n_834) );
INVx1_ASAP7_75t_L g825 ( .A(n_639), .Y(n_825) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_644), .A2(n_652), .B1(n_687), .B2(n_761), .C(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_646), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g711 ( .A(n_647), .Y(n_711) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_649), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g826 ( .A(n_649), .B(n_677), .Y(n_826) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g662 ( .A(n_650), .Y(n_662) );
AND3x1_ASAP7_75t_L g835 ( .A(n_650), .B(n_836), .C(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g705 ( .A(n_654), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g775 ( .A(n_657), .Y(n_775) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g751 ( .A(n_659), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g778 ( .A(n_659), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_669), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2x1_ASAP7_75t_L g676 ( .A(n_662), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g743 ( .A(n_663), .Y(n_743) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g699 ( .A(n_667), .Y(n_699) );
OR2x2_ASAP7_75t_L g678 ( .A(n_668), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g791 ( .A(n_668), .Y(n_791) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_670), .B(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
OR2x2_ASAP7_75t_L g747 ( .A(n_671), .B(n_695), .Y(n_747) );
INVx2_ASAP7_75t_L g836 ( .A(n_671), .Y(n_836) );
INVx1_ASAP7_75t_L g710 ( .A(n_672), .Y(n_710) );
NOR4xp25_ASAP7_75t_L g840 ( .A(n_672), .B(n_703), .C(n_841), .D(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_673), .Y(n_842) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx3_ASAP7_75t_L g828 ( .A(n_674), .Y(n_828) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_680), .B(n_683), .C(n_691), .Y(n_675) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g815 ( .A(n_678), .Y(n_815) );
INVx2_ASAP7_75t_L g800 ( .A(n_679), .Y(n_800) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_681), .A2(n_684), .B(n_687), .Y(n_683) );
OR2x2_ASAP7_75t_L g767 ( .A(n_682), .B(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g785 ( .A(n_682), .B(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g701 ( .A(n_686), .Y(n_701) );
AND2x4_ASAP7_75t_SL g790 ( .A(n_686), .B(n_791), .Y(n_790) );
INVx3_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_689), .Y(n_756) );
INVx1_ASAP7_75t_L g763 ( .A(n_690), .Y(n_763) );
AOI32xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_697), .A3(n_699), .B1(n_700), .B2(n_704), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_694), .B(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_694), .Y(n_755) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g772 ( .A(n_695), .B(n_710), .Y(n_772) );
INVx2_ASAP7_75t_L g786 ( .A(n_695), .Y(n_786) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g765 ( .A(n_703), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B(n_712), .C(n_728), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .B(n_718), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g769 ( .A(n_717), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_717), .B(n_804), .Y(n_803) );
OAI32xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .A3(n_722), .B1(n_724), .B2(n_727), .Y(n_718) );
INVx1_ASAP7_75t_L g804 ( .A(n_719), .Y(n_804) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g796 ( .A(n_721), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_805), .Y(n_733) );
NAND4xp25_ASAP7_75t_L g734 ( .A(n_735), .B(n_760), .C(n_773), .D(n_801), .Y(n_734) );
NOR2xp67_ASAP7_75t_L g735 ( .A(n_736), .B(n_748), .Y(n_735) );
OAI32xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .A3(n_740), .B1(n_741), .B2(n_747), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g787 ( .A(n_739), .B(n_788), .Y(n_787) );
OAI32xp33_ASAP7_75t_L g792 ( .A1(n_739), .A2(n_793), .A3(n_794), .B1(n_796), .B2(n_798), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_740), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_742), .B(n_807), .Y(n_806) );
INVx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g799 ( .A(n_745), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g831 ( .A(n_745), .Y(n_831) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g795 ( .A(n_746), .Y(n_795) );
OAI22x1_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_754), .B1(n_756), .B2(n_757), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_758), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2x1_ASAP7_75t_L g824 ( .A(n_762), .B(n_825), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B1(n_769), .B2(n_770), .Y(n_764) );
NAND2x1_ASAP7_75t_L g830 ( .A(n_766), .B(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g841 ( .A(n_766), .Y(n_841) );
INVx2_ASAP7_75t_L g782 ( .A(n_768), .Y(n_782) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NOR3xp33_ASAP7_75t_SL g773 ( .A(n_774), .B(n_783), .C(n_792), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_780), .Y(n_774) );
NAND2xp33_ASAP7_75t_L g802 ( .A(n_776), .B(n_803), .Y(n_802) );
INVx2_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND2x4_ASAP7_75t_L g838 ( .A(n_782), .B(n_839), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B(n_789), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AND2x4_ASAP7_75t_L g809 ( .A(n_786), .B(n_810), .Y(n_809) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_788), .Y(n_808) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND3xp33_ASAP7_75t_SL g805 ( .A(n_806), .B(n_811), .C(n_823), .Y(n_805) );
AND2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g814 ( .A(n_810), .Y(n_814) );
AOI222xp33_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_815), .B1(n_816), .B2(n_817), .C1(n_820), .C2(n_821), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
O2A1O1Ixp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_826), .B(n_827), .C(n_829), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_861), .B(n_865), .Y(n_844) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_857), .B(n_859), .C(n_860), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_849), .Y(n_846) );
INVx5_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
XOR2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_854), .Y(n_850) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx6f_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
CKINVDCx11_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx10_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AND2x6_ASAP7_75t_L g876 ( .A(n_871), .B(n_877), .Y(n_876) );
BUFx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
INVx5_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
BUFx8_ASAP7_75t_L g880 ( .A(n_876), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_880), .Y(n_879) );
endmodule