module fake_jpeg_17995_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_43),
.B(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_56),
.Y(n_69)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_10),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_60),
.Y(n_71)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_9),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_64),
.Y(n_88)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_9),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_67),
.Y(n_94)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_15),
.B1(n_39),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_68),
.A2(n_74),
.B1(n_80),
.B2(n_89),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_30),
.B1(n_37),
.B2(n_33),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_76),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_99),
.B1(n_110),
.B2(n_113),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_23),
.B1(n_22),
.B2(n_20),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_101),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_85),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_37),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_63),
.B1(n_45),
.B2(n_47),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_23),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_95),
.B(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_54),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_27),
.B1(n_26),
.B2(n_8),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_105),
.B1(n_80),
.B2(n_72),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_0),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_18),
.B1(n_8),
.B2(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_38),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_112),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_27),
.B1(n_26),
.B2(n_8),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_59),
.A2(n_36),
.B1(n_34),
.B2(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_38),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_38),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_118),
.A2(n_151),
.B(n_76),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_123),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_41),
.A3(n_66),
.B1(n_26),
.B2(n_54),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_77),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_131),
.B1(n_133),
.B2(n_137),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_149),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_87),
.B1(n_97),
.B2(n_109),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_84),
.A2(n_5),
.B1(n_7),
.B2(n_28),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_28),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_71),
.B(n_7),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_51),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_51),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_152),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_48),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_48),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_106),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_95),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_175),
.C(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_149),
.B1(n_147),
.B2(n_127),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_162),
.B1(n_165),
.B2(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_102),
.B1(n_73),
.B2(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_102),
.B1(n_73),
.B2(n_84),
.Y(n_165)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_169),
.B(n_100),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_103),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_48),
.C(n_51),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_97),
.B1(n_109),
.B2(n_87),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_142),
.B1(n_126),
.B2(n_134),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_141),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_120),
.A2(n_77),
.B1(n_108),
.B2(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_111),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_151),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_116),
.Y(n_197)
);

XOR2x1_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_118),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_190),
.A2(n_208),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_127),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_130),
.C(n_122),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_216),
.C(n_119),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_156),
.C(n_188),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_135),
.B(n_148),
.C(n_124),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_203),
.B1(n_171),
.B2(n_167),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_115),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_201),
.B(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_145),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_135),
.B1(n_124),
.B2(n_151),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_206),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_136),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_128),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_163),
.B(n_139),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_125),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_114),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_132),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_224),
.C(n_229),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_183),
.B1(n_184),
.B2(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_209),
.B1(n_192),
.B2(n_203),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_185),
.C(n_158),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_232),
.B(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_175),
.C(n_162),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_SL g234 ( 
.A1(n_190),
.A2(n_176),
.A3(n_216),
.B1(n_204),
.B2(n_197),
.C1(n_206),
.C2(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_195),
.C(n_212),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.C(n_178),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_194),
.C(n_213),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_215),
.B1(n_171),
.B2(n_205),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_251),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_199),
.A3(n_208),
.B1(n_192),
.B2(n_217),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_254),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_208),
.B1(n_200),
.B2(n_211),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_228),
.B1(n_229),
.B2(n_236),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_202),
.B1(n_207),
.B2(n_166),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_172),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_250),
.C(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_172),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_178),
.B(n_166),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_189),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_233),
.B(n_189),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_181),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_257),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_226),
.B(n_157),
.Y(n_258)
);

NOR3xp33_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_230),
.C(n_222),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_234),
.A3(n_231),
.B1(n_218),
.B2(n_227),
.C1(n_221),
.C2(n_223),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_260),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_227),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_251),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_255),
.B(n_225),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_246),
.B1(n_243),
.B2(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_244),
.B1(n_242),
.B2(n_220),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_231),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_270),
.C(n_253),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_218),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_250),
.C(n_248),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_245),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_281),
.B1(n_282),
.B2(n_262),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_262),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_225),
.B1(n_238),
.B2(n_76),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_269),
.B1(n_263),
.B2(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_261),
.B1(n_267),
.B2(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_287),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_288),
.B(n_287),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_294),
.C(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_289),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_297),
.B(n_298),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_300),
.Y(n_302)
);


endmodule