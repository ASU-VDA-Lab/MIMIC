module fake_jpeg_17660_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_36),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_30),
.B1(n_20),
.B2(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_48),
.B1(n_46),
.B2(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_32),
.B1(n_30),
.B2(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_22),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_19),
.B1(n_28),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_79),
.Y(n_99)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

NAND2x1p5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_35),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_74),
.B(n_85),
.Y(n_96)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_66),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_28),
.B1(n_19),
.B2(n_26),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_64),
.B1(n_81),
.B2(n_60),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_19),
.B1(n_16),
.B2(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_73),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_35),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_25),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_18),
.C(n_24),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_2),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_35),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_108),
.Y(n_133)
);

AOI21x1_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_29),
.B(n_21),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_106),
.B(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_110),
.B1(n_58),
.B2(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_18),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_125),
.B1(n_134),
.B2(n_8),
.Y(n_146)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_18),
.C(n_78),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_22),
.C(n_9),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_69),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_101),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_4),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_106),
.A3(n_105),
.B1(n_88),
.B2(n_93),
.C1(n_110),
.C2(n_100),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_68),
.B(n_65),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_121),
.B(n_131),
.Y(n_141)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_22),
.Y(n_127)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_90),
.B(n_72),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_95),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_150),
.B(n_132),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_142),
.C(n_146),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_101),
.B1(n_109),
.B2(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_143),
.B1(n_113),
.B2(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_151),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_106),
.B(n_109),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_93),
.B1(n_9),
.B2(n_8),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_62),
.B(n_67),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_10),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_22),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_126),
.C(n_125),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_142),
.B1(n_154),
.B2(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_112),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_170),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_135),
.B(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_116),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_174),
.C(n_156),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_111),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_141),
.B(n_140),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_167),
.B(n_159),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_173),
.B1(n_171),
.B2(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_186),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_174),
.B(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_173),
.C(n_128),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_118),
.C(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_183),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_194),
.B(n_180),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_180),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_161),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_182),
.C(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_205),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_12),
.B(n_13),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_198),
.C(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_185),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_186),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_200),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_204),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_213),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_214),
.B(n_215),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_202),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_201),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_217),
.C(n_216),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_14),
.C(n_15),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_220),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_221),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_222),
.Y(n_225)
);


endmodule