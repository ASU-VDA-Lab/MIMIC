module real_jpeg_27889_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_0),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_0),
.A2(n_30),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_0),
.B(n_32),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_0),
.A2(n_61),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_0),
.B(n_61),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_0),
.B(n_74),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_0),
.A2(n_136),
.B1(n_138),
.B2(n_204),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_0),
.A2(n_33),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_2),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_2),
.A2(n_56),
.B1(n_58),
.B2(n_96),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_96),
.Y(n_224)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_5),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_101),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_5),
.A2(n_56),
.B1(n_58),
.B2(n_101),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_101),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_7),
.A2(n_37),
.B1(n_56),
.B2(n_58),
.Y(n_157)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_9),
.A2(n_56),
.B1(n_58),
.B2(n_104),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_104),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_104),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_10),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_28),
.B1(n_56),
.B2(n_58),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_10),
.A2(n_28),
.B1(n_61),
.B2(n_62),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_94),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_11),
.A2(n_56),
.B1(n_58),
.B2(n_94),
.Y(n_197)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_13),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_111),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_111),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_111),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_17),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_17),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_22),
.B(n_43),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_24),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_35),
.B(n_108),
.C(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_32),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_32),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_29),
.A2(n_32),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_29),
.A2(n_32),
.B1(n_145),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_29),
.A2(n_32),
.B1(n_164),
.B2(n_259),
.Y(n_258)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_68),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_68),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_33),
.A2(n_62),
.A3(n_68),
.B1(n_221),
.B2(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_34),
.B(n_108),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_82),
.B(n_333),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_75),
.C(n_77),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_44),
.A2(n_45),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_64),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_46),
.B(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_48),
.A2(n_79),
.B1(n_81),
.B2(n_286),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_52),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_52),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_52),
.A2(n_64),
.B1(n_312),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_63),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_59),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_53),
.A2(n_59),
.B1(n_134),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_53),
.A2(n_59),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_53),
.A2(n_59),
.B1(n_178),
.B2(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_53),
.B(n_108),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_53),
.A2(n_59),
.B1(n_100),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_53),
.A2(n_59),
.B1(n_63),
.B2(n_268),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_54),
.A2(n_58),
.A3(n_61),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_55),
.B(n_56),
.Y(n_182)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_56),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_61),
.B(n_72),
.Y(n_229)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_64),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_73),
.B2(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_65),
.A2(n_66),
.B1(n_74),
.B2(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_66),
.A2(n_74),
.B1(n_93),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_74),
.B1(n_148),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_66),
.A2(n_74),
.B1(n_166),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_71),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_71),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_67),
.A2(n_71),
.B1(n_95),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_67),
.A2(n_71),
.B1(n_125),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_67),
.A2(n_71),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_75),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_79),
.A2(n_81),
.B1(n_110),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_79),
.A2(n_81),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_326),
.B(n_332),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_303),
.A3(n_322),
.B1(n_324),
.B2(n_325),
.C(n_336),
.Y(n_83)
);

AOI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_255),
.A3(n_292),
.B1(n_297),
.B2(n_302),
.C(n_337),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_150),
.C(n_168),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_129),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_87),
.B(n_129),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_112),
.C(n_121),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_88),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_106),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_98),
.C(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_102),
.A2(n_105),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_102),
.A2(n_105),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_108),
.B(n_138),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_112),
.A2(n_121),
.B1(n_122),
.B2(n_253),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_112),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_116),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g205 ( 
.A(n_117),
.Y(n_205)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_123),
.B(n_240),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_126),
.B(n_128),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_127),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_140),
.C(n_141),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_135),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_136),
.A2(n_138),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_136),
.A2(n_197),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_136),
.A2(n_138),
.B1(n_192),
.B2(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_136),
.A2(n_138),
.B(n_157),
.Y(n_270)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_146),
.C(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_151),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_152),
.B(n_153),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_167),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_155),
.B(n_160),
.C(n_167),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_156),
.B(n_158),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_159),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_249),
.B(n_254),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_235),
.B(n_248),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_214),
.B(n_234),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_193),
.B(n_213),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_183),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_173),
.B(n_183),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_191),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_201),
.B(n_212),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_200),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_207),
.B(n_211),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_226),
.C(n_233),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_244),
.C(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_272),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.C(n_271),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_263),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_257),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.CI(n_262),
.CON(n_257),
.SN(n_257)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_260),
.C(n_262),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_269),
.B2(n_270),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_264),
.B(n_270),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_270),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_284),
.B(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_290),
.B2(n_291),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_281),
.C(n_291),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.B(n_280),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_279),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

FAx1_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_305),
.CI(n_314),
.CON(n_304),
.SN(n_304)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_315),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_315),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_313),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_307),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_309),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_320),
.C(n_321),
.Y(n_327)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule