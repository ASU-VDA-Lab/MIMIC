module fake_jpeg_17105_n_97 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_97);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_24),
.Y(n_49)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_35)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_32),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_5),
.B1(n_11),
.B2(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_15),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_9),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_19),
.B1(n_15),
.B2(n_17),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_45),
.B1(n_50),
.B2(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_17),
.B1(n_21),
.B2(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_42),
.B1(n_35),
.B2(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_18),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_26),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_18),
.C(n_22),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_18),
.B(n_11),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_42),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_29),
.B(n_31),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_66),
.B2(n_51),
.Y(n_70)
);

AOI22x1_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_45),
.B1(n_50),
.B2(n_47),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_52),
.B(n_49),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_36),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_39),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_72),
.C(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_74),
.B1(n_66),
.B2(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_77),
.B(n_64),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_57),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_75),
.C(n_62),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_61),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_81),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_55),
.B(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

OAI31xp67_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_62),
.A3(n_76),
.B(n_80),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_78),
.C(n_79),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_87),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_87),
.C(n_86),
.Y(n_94)
);

AOI211xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.C(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_92),
.B(n_96),
.Y(n_97)
);


endmodule