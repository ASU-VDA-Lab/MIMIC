module fake_netlist_6_3794_n_1658 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1658);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1658;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_142;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_141;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_17),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_25),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_39),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_55),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_54),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_2),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_131),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_30),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_74),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_19),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_28),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_35),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_15),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_39),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_71),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_12),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_35),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_21),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_24),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_34),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_25),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_18),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_22),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_58),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_123),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_57),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_47),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_66),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_52),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_38),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_64),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_10),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_53),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_42),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_10),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_24),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_49),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_120),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_135),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_11),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_59),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_137),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_117),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_21),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_6),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_43),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_27),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_103),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_68),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_45),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_14),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_79),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_18),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_22),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_7),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_29),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_51),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_23),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_100),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_14),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_121),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_133),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_136),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_90),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_95),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_28),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_60),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_16),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_122),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_26),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_87),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_84),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_114),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_34),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_104),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_7),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_61),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_77),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_23),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_112),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_33),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_50),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_45),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_29),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_19),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_38),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_36),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_9),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_132),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_3),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_93),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_183),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_187),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_174),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_183),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_183),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_179),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_181),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_166),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_189),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_193),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_147),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_200),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_151),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_243),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_250),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_147),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_212),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_214),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_158),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_187),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_241),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_152),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_152),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_216),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_145),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_145),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_145),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_217),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_224),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_146),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_203),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_160),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_203),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_225),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_170),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_151),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_234),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_160),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_185),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_191),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_195),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_256),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_320),
.A2(n_208),
.B(n_202),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_288),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_312),
.A2(n_229),
.B1(n_259),
.B2(n_155),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_256),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_286),
.Y(n_365)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_234),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_184),
.Y(n_368)
);

AND3x2_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_283),
.C(n_188),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_289),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_289),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_290),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_287),
.B(n_159),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_188),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_292),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_291),
.B(n_141),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_144),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_293),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_295),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_296),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_296),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_300),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_300),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_294),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_302),
.B(n_141),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_302),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_287),
.B(n_219),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_333),
.B(n_306),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_333),
.B(n_148),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_307),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_142),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_324),
.B(n_227),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_310),
.B(n_163),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_310),
.B(n_142),
.Y(n_403)
);

AOI22x1_ASAP7_75t_SL g404 ( 
.A1(n_314),
.A2(n_167),
.B1(n_172),
.B2(n_171),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_311),
.B(n_143),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_297),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_313),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_383),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_383),
.Y(n_411)
);

AO21x2_ASAP7_75t_L g412 ( 
.A1(n_378),
.A2(n_175),
.B(n_164),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_357),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_358),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_377),
.B(n_298),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g416 ( 
.A1(n_400),
.A2(n_343),
.B(n_308),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_394),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_360),
.A2(n_172),
.B1(n_171),
.B2(n_264),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_390),
.B(n_303),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_337),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

AOI22x1_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_343),
.B1(n_344),
.B2(n_274),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_394),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_351),
.B(n_177),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

BUFx6f_ASAP7_75t_SL g440 ( 
.A(n_374),
.Y(n_440)
);

BUFx6f_ASAP7_75t_SL g441 ( 
.A(n_374),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_350),
.B(n_317),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_363),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_350),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_395),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_349),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_395),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_371),
.B(n_318),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_349),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_352),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_389),
.A2(n_173),
.B1(n_272),
.B2(n_236),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_389),
.B(n_330),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_362),
.B(n_334),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_358),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_354),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_395),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_393),
.B(n_362),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_356),
.B(n_301),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

AND3x2_ASAP7_75t_L g476 ( 
.A(n_356),
.B(n_149),
.C(n_304),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_378),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_353),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_353),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_355),
.Y(n_484)
);

NOR2x1p5_ASAP7_75t_L g485 ( 
.A(n_391),
.B(n_155),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_404),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_361),
.B(n_316),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_363),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_361),
.B(n_335),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_367),
.B(n_315),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_407),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_393),
.B(n_340),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_367),
.B(n_315),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_355),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_374),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_363),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_391),
.B(n_321),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_359),
.Y(n_503)
);

AOI21x1_ASAP7_75t_L g504 ( 
.A1(n_375),
.A2(n_323),
.B(n_322),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_380),
.A2(n_275),
.B1(n_231),
.B2(n_244),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_380),
.A2(n_273),
.B1(n_268),
.B2(n_281),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_363),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_366),
.B(n_322),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_375),
.B(n_180),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_359),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_374),
.Y(n_513)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_399),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_365),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_399),
.B(n_321),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_365),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g519 ( 
.A1(n_403),
.A2(n_192),
.B(n_190),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_403),
.B(n_327),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_366),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_366),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_402),
.B(n_143),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_405),
.B(n_323),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_405),
.A2(n_232),
.B1(n_213),
.B2(n_218),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_409),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_372),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_372),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_380),
.B(n_321),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_380),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_397),
.A2(n_167),
.B1(n_258),
.B2(n_162),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_373),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_408),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_373),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_376),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_376),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_381),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_375),
.B(n_162),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_381),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_397),
.B(n_344),
.C(n_336),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_369),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_382),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_382),
.B(n_328),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_408),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_397),
.B(n_150),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_397),
.B(n_150),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_386),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_368),
.B(n_153),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_439),
.B(n_342),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_514),
.B(n_369),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_425),
.B(n_194),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_410),
.B(n_270),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_L g556 ( 
.A(n_492),
.B(n_211),
.C(n_156),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_439),
.B(n_442),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_433),
.A2(n_254),
.B1(n_267),
.B2(n_252),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_478),
.B(n_402),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_439),
.B(n_386),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_433),
.A2(n_247),
.B1(n_228),
.B2(n_158),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_442),
.B(n_387),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_425),
.B(n_198),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_410),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_442),
.B(n_387),
.Y(n_566)
);

AND2x4_ASAP7_75t_SL g567 ( 
.A(n_426),
.B(n_279),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_454),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_454),
.B(n_392),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_454),
.B(n_392),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_455),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_471),
.B(n_398),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_419),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_471),
.B(n_398),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_462),
.B(n_199),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_520),
.B(n_284),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_531),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_411),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_520),
.B(n_342),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_417),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_529),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_466),
.B(n_153),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_531),
.Y(n_584)
);

OAI22xp33_ASAP7_75t_L g585 ( 
.A1(n_464),
.A2(n_168),
.B1(n_165),
.B2(n_258),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_471),
.B(n_401),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_464),
.A2(n_278),
.B1(n_261),
.B2(n_264),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_457),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_430),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_444),
.B(n_154),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_460),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_433),
.A2(n_435),
.B1(n_438),
.B2(n_431),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_417),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_499),
.A2(n_154),
.B1(n_157),
.B2(n_161),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_431),
.A2(n_158),
.B1(n_205),
.B2(n_257),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_524),
.B(n_363),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_457),
.B(n_363),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_419),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_419),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_461),
.B(n_364),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_470),
.B(n_364),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_452),
.Y(n_603)
);

BUFx5_ASAP7_75t_L g604 ( 
.A(n_435),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_475),
.B(n_209),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_458),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_423),
.B(n_364),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_423),
.B(n_364),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_413),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_499),
.A2(n_513),
.B1(n_475),
.B2(n_441),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

BUFx8_ASAP7_75t_L g612 ( 
.A(n_428),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_428),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_513),
.A2(n_230),
.B1(n_262),
.B2(n_265),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_452),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_483),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_453),
.B(n_158),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_456),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_456),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_416),
.B(n_157),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_453),
.B(n_158),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_453),
.B(n_158),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_438),
.B(n_364),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_493),
.B(n_364),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_426),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_469),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_497),
.B(n_364),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_416),
.B(n_161),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_485),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_453),
.B(n_158),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_543),
.B(n_485),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_468),
.B(n_158),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_465),
.B(n_169),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_483),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_429),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_530),
.B(n_388),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_484),
.B(n_498),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_538),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_426),
.B(n_169),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_496),
.B(n_472),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_498),
.B(n_503),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_511),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_473),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_525),
.B(n_246),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_542),
.B(n_279),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_462),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_440),
.A2(n_260),
.B1(n_246),
.B2(n_253),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_512),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_512),
.B(n_388),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_543),
.B(n_346),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_SL g654 ( 
.A(n_468),
.B(n_505),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_426),
.B(n_279),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_468),
.B(n_388),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_468),
.B(n_505),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_515),
.B(n_388),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_511),
.B(n_253),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_487),
.B(n_260),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_540),
.B(n_346),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_476),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_551),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_456),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_518),
.B(n_388),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_459),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_527),
.B(n_215),
.Y(n_668)
);

BUFx5_ASAP7_75t_L g669 ( 
.A(n_462),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_468),
.B(n_238),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_242),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_427),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_531),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_536),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_468),
.B(n_248),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_537),
.B(n_541),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_459),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_537),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_501),
.B(n_263),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_488),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_440),
.A2(n_282),
.B1(n_263),
.B2(n_255),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_541),
.B(n_368),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_549),
.B(n_328),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_532),
.B(n_517),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_532),
.B(n_347),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_549),
.B(n_329),
.Y(n_688)
);

AO221x1_ASAP7_75t_L g689 ( 
.A1(n_418),
.A2(n_404),
.B1(n_348),
.B2(n_347),
.C(n_339),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_459),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_547),
.B(n_348),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_522),
.B(n_412),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_415),
.B(n_282),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_474),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_420),
.B(n_176),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_538),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_505),
.B(n_329),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_505),
.B(n_178),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_505),
.B(n_182),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_531),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_522),
.B(n_186),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_412),
.B(n_197),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_412),
.B(n_201),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_519),
.B(n_339),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_548),
.B(n_337),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_505),
.B(n_204),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_440),
.B(n_441),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_544),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_562),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_571),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_578),
.Y(n_712)
);

AND2x6_ASAP7_75t_SL g713 ( 
.A(n_647),
.B(n_486),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_592),
.B(n_519),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_582),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_582),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_552),
.B(n_488),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_609),
.B(n_510),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_552),
.B(n_488),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_588),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_SL g722 ( 
.A1(n_591),
.A2(n_165),
.B1(n_168),
.B2(n_261),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_592),
.B(n_519),
.Y(n_723)
);

AND2x2_ASAP7_75t_SL g724 ( 
.A(n_567),
.B(n_440),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_565),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_629),
.B(n_506),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_649),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_626),
.A2(n_504),
.B(n_511),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_649),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_604),
.B(n_544),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_649),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_682),
.Y(n_732)
);

BUFx4f_ASAP7_75t_L g733 ( 
.A(n_634),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_604),
.B(n_511),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_604),
.B(n_511),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_682),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_578),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_601),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_614),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_593),
.Y(n_740)
);

INVx5_ASAP7_75t_L g741 ( 
.A(n_682),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_557),
.A2(n_441),
.B1(n_511),
.B2(n_523),
.Y(n_742)
);

OAI21xp5_ASAP7_75t_L g743 ( 
.A1(n_561),
.A2(n_504),
.B(n_511),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_606),
.B(n_427),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_593),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_604),
.B(n_534),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_613),
.Y(n_747)
);

NAND3xp33_ASAP7_75t_SL g748 ( 
.A(n_556),
.B(n_576),
.C(n_660),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_682),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_576),
.B(n_441),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_613),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_646),
.B(n_583),
.Y(n_752)
);

INVx5_ASAP7_75t_L g753 ( 
.A(n_554),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_628),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_604),
.B(n_550),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_568),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_614),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_629),
.B(n_414),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_612),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_634),
.B(n_508),
.Y(n_760)
);

OR2x2_ASAP7_75t_SL g761 ( 
.A(n_687),
.B(n_269),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_SL g762 ( 
.A(n_585),
.B(n_276),
.C(n_277),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_628),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_632),
.B(n_508),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_604),
.B(n_550),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_558),
.B(n_550),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_641),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_709),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_605),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_605),
.B(n_430),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_558),
.B(n_534),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_709),
.Y(n_772)
);

OR2x2_ASAP7_75t_SL g773 ( 
.A(n_643),
.B(n_277),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_581),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_590),
.B(n_414),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_672),
.A2(n_528),
.B(n_508),
.C(n_535),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_590),
.B(n_414),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_561),
.B(n_546),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_663),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_686),
.B(n_414),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_636),
.B(n_443),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_610),
.A2(n_528),
.B1(n_545),
.B2(n_280),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_580),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_568),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_555),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_623),
.A2(n_528),
.B(n_535),
.C(n_534),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_553),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_595),
.A2(n_507),
.B1(n_210),
.B2(n_245),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_653),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_SL g791 ( 
.A(n_585),
.B(n_206),
.C(n_240),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_708),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_653),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_669),
.B(n_445),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_579),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_694),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_579),
.B(n_674),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_611),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_573),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_546),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_615),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_636),
.B(n_443),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_619),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_655),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_669),
.B(n_445),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_648),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_637),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_651),
.Y(n_808)
);

BUFx2_ASAP7_75t_SL g809 ( 
.A(n_674),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_642),
.B(n_443),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_661),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_598),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_644),
.B(n_546),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_678),
.B(n_535),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_704),
.B(n_443),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_700),
.B(n_490),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_664),
.A2(n_467),
.B1(n_490),
.B2(n_500),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_673),
.B(n_467),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_691),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_705),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_567),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_R g822 ( 
.A(n_707),
.B(n_490),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_599),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_675),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_669),
.B(n_445),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_662),
.Y(n_826)
);

AND2x6_ASAP7_75t_SL g827 ( 
.A(n_647),
.B(n_207),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_705),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_700),
.B(n_490),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_577),
.B(n_467),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_677),
.B(n_467),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_680),
.B(n_500),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_693),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_693),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_SL g835 ( 
.A(n_587),
.B(n_220),
.C(n_221),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_607),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_560),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_608),
.B(n_500),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_669),
.B(n_500),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_563),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_623),
.B(n_631),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_603),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_669),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_617),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_631),
.A2(n_526),
.B(n_421),
.C(n_422),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_669),
.B(n_421),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_566),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_681),
.A2(n_526),
.B(n_422),
.C(n_424),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_695),
.A2(n_436),
.B1(n_446),
.B2(n_509),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_695),
.B(n_424),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_645),
.B(n_445),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_569),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_684),
.B(n_432),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_570),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_627),
.B(n_432),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_645),
.B(n_521),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_630),
.B(n_437),
.Y(n_857)
);

CKINVDCx8_ASAP7_75t_R g858 ( 
.A(n_681),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_702),
.A2(n_509),
.B1(n_436),
.B2(n_446),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_645),
.B(n_521),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_577),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_596),
.B(n_437),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_618),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_559),
.B(n_447),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_645),
.B(n_521),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_639),
.B(n_447),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_701),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_616),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_703),
.A2(n_436),
.B1(n_446),
.B2(n_509),
.Y(n_869)
);

OR2x4_ASAP7_75t_L g870 ( 
.A(n_689),
.B(n_222),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_595),
.B(n_448),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_584),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_572),
.B(n_448),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_L g874 ( 
.A(n_554),
.B(n_429),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_652),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_658),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_707),
.A2(n_436),
.B1(n_446),
.B2(n_509),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_666),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_575),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_597),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_574),
.B(n_451),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_584),
.B(n_683),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_638),
.B(n_521),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_668),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_752),
.B(n_671),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_710),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_748),
.A2(n_650),
.B1(n_659),
.B2(n_594),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_SL g888 ( 
.A(n_833),
.B(n_587),
.C(n_239),
.Y(n_888)
);

OAI22x1_ASAP7_75t_L g889 ( 
.A1(n_834),
.A2(n_237),
.B1(n_226),
.B2(n_233),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_725),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_841),
.A2(n_633),
.B(n_625),
.C(n_624),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_R g892 ( 
.A(n_754),
.B(n_554),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_711),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_750),
.A2(n_586),
.B(n_692),
.C(n_600),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_714),
.A2(n_589),
.B1(n_575),
.B2(n_602),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_714),
.A2(n_589),
.B1(n_620),
.B2(n_625),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_828),
.B(n_621),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_730),
.A2(n_620),
.B(n_624),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_759),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_784),
.B(n_685),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_745),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_721),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_883),
.A2(n_657),
.B(n_633),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_769),
.B(n_688),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_747),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_843),
.A2(n_657),
.B(n_656),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_790),
.B(n_622),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_858),
.B(n_698),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_769),
.B(n_698),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_741),
.A2(n_656),
.B(n_434),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_786),
.B(n_737),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_741),
.A2(n_429),
.B(n_434),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_840),
.B(n_554),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_715),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_826),
.B(n_712),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_744),
.A2(n_706),
.B(n_699),
.C(n_635),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_726),
.B(n_819),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_738),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_741),
.A2(n_749),
.B(n_794),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_727),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_723),
.A2(n_665),
.B1(n_690),
.B2(n_679),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_740),
.B(n_667),
.Y(n_922)
);

OAI21xp33_ASAP7_75t_L g923 ( 
.A1(n_762),
.A2(n_223),
.B(n_235),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_868),
.A2(n_676),
.B(n_670),
.C(n_697),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_760),
.B(n_564),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_741),
.A2(n_429),
.B(n_434),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_793),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_727),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_779),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_806),
.B(n_564),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_717),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_749),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_847),
.B(n_564),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_763),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_852),
.A2(n_854),
.B(n_780),
.C(n_802),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_749),
.A2(n_429),
.B(n_434),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_739),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_757),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_SL g939 ( 
.A(n_722),
.B(n_676),
.C(n_670),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_723),
.A2(n_697),
.B1(n_429),
.B2(n_434),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_763),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_751),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_763),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_788),
.A2(n_451),
.B(n_463),
.C(n_502),
.Y(n_944)
);

XOR2xp5_ASAP7_75t_L g945 ( 
.A(n_724),
.B(n_56),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_767),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_749),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_805),
.A2(n_825),
.B(n_735),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_836),
.B(n_884),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_734),
.A2(n_434),
.B(n_449),
.Y(n_950)
);

INVx6_ASAP7_75t_L g951 ( 
.A(n_713),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_795),
.A2(n_449),
.B1(n_450),
.B2(n_502),
.Y(n_952)
);

NOR2x1_ASAP7_75t_R g953 ( 
.A(n_804),
.B(n_449),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_867),
.B(n_480),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_880),
.B(n_480),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_774),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_798),
.B(n_481),
.Y(n_957)
);

AO32x2_ASAP7_75t_L g958 ( 
.A1(n_789),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_958)
);

INVx6_ASAP7_75t_L g959 ( 
.A(n_827),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_727),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_787),
.A2(n_776),
.B(n_728),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_733),
.B(n_449),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_760),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_801),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_882),
.A2(n_781),
.B(n_775),
.C(n_777),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_795),
.A2(n_449),
.B1(n_450),
.B2(n_495),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_820),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_803),
.B(n_481),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_734),
.A2(n_449),
.B(n_450),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_807),
.B(n_489),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_735),
.A2(n_450),
.B(n_654),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_789),
.A2(n_489),
.B(n_495),
.C(n_494),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_809),
.B(n_450),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_837),
.A2(n_477),
.B1(n_494),
.B2(n_463),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_728),
.A2(n_516),
.B(n_491),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_743),
.A2(n_450),
.B(n_491),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_808),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_758),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_797),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_811),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_766),
.A2(n_477),
.B1(n_516),
.B2(n_479),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_824),
.B(n_516),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_743),
.A2(n_491),
.B(n_479),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_797),
.Y(n_984)
);

AO32x2_ASAP7_75t_L g985 ( 
.A1(n_756),
.A2(n_1),
.A3(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_864),
.A2(n_479),
.B(n_474),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_SL g987 ( 
.A1(n_761),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_730),
.A2(n_474),
.B(n_83),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_718),
.A2(n_82),
.B1(n_127),
.B2(n_125),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_SL g990 ( 
.A1(n_783),
.A2(n_13),
.B(n_20),
.C(n_31),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_791),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_718),
.B(n_85),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_782),
.A2(n_20),
.B(n_32),
.C(n_37),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_839),
.A2(n_86),
.B(n_124),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_SL g995 ( 
.A1(n_773),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_837),
.B(n_44),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_837),
.B(n_44),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_839),
.A2(n_846),
.B(n_815),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_846),
.A2(n_91),
.B(n_113),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_768),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_835),
.A2(n_46),
.B(n_48),
.C(n_50),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_720),
.A2(n_63),
.B1(n_67),
.B2(n_69),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_879),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_815),
.A2(n_72),
.B(n_76),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_764),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_746),
.A2(n_88),
.B(n_96),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_864),
.A2(n_845),
.B(n_881),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_866),
.A2(n_97),
.B(n_101),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_772),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_792),
.A2(n_107),
.B(n_108),
.C(n_109),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_716),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_796),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_866),
.A2(n_110),
.B(n_111),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_832),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_850),
.A2(n_742),
.B(n_810),
.C(n_771),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_719),
.B(n_879),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_832),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_821),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_799),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_932),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_961),
.A2(n_848),
.B(n_770),
.Y(n_1021)
);

AO22x1_ASAP7_75t_L g1022 ( 
.A1(n_991),
.A2(n_764),
.B1(n_879),
.B2(n_753),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_885),
.B(n_878),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1014),
.B(n_876),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1017),
.B(n_875),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_SL g1026 ( 
.A1(n_996),
.A2(n_766),
.B(n_771),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_942),
.B(n_756),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_946),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_976),
.A2(n_838),
.B(n_855),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_950),
.A2(n_969),
.B(n_983),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_942),
.B(n_736),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_886),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1007),
.A2(n_874),
.B(n_857),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_948),
.A2(n_838),
.B(n_862),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_893),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_935),
.B(n_814),
.Y(n_1036)
);

AOI31xp67_ASAP7_75t_L g1037 ( 
.A1(n_909),
.A2(n_887),
.A3(n_933),
.B(n_913),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_998),
.A2(n_872),
.B(n_861),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_895),
.A2(n_871),
.A3(n_765),
.B(n_755),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_896),
.A2(n_814),
.B(n_813),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_927),
.B(n_736),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_949),
.B(n_813),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_927),
.B(n_785),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_901),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1007),
.A2(n_881),
.B(n_873),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_917),
.B(n_812),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_930),
.A2(n_853),
.B(n_817),
.C(n_778),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_908),
.A2(n_870),
.B1(n_861),
.B2(n_785),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_898),
.A2(n_800),
.B(n_853),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_915),
.B(n_870),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_890),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_978),
.B(n_863),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_905),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_967),
.B(n_844),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_902),
.B(n_800),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_1001),
.A2(n_873),
.B(n_818),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_R g1057 ( 
.A(n_892),
.B(n_822),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_963),
.B(n_716),
.Y(n_1058)
);

AO21x2_ASAP7_75t_L g1059 ( 
.A1(n_961),
.A2(n_859),
.B(n_869),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_891),
.A2(n_753),
.B(n_856),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_918),
.B(n_729),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_932),
.B(n_729),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_981),
.A2(n_831),
.B(n_746),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_964),
.Y(n_1064)
);

NOR4xp25_ASAP7_75t_L g1065 ( 
.A(n_993),
.B(n_755),
.C(n_765),
.D(n_871),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_977),
.B(n_731),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_941),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_900),
.B(n_823),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_956),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_911),
.B(n_842),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_980),
.B(n_731),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_981),
.A2(n_816),
.B(n_829),
.Y(n_1072)
);

AOI221xp5_ASAP7_75t_SL g1073 ( 
.A1(n_987),
.A2(n_732),
.B1(n_851),
.B2(n_860),
.C(n_865),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1000),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_SL g1075 ( 
.A(n_888),
.B(n_849),
.C(n_877),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_894),
.A2(n_903),
.B(n_916),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_971),
.A2(n_753),
.B(n_732),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1009),
.B(n_830),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_1018),
.B(n_753),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_986),
.A2(n_830),
.B(n_975),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_945),
.A2(n_830),
.B1(n_997),
.B2(n_904),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_972),
.A2(n_830),
.B(n_975),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_923),
.B(n_830),
.C(n_939),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_940),
.A2(n_921),
.A3(n_924),
.B(n_988),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_955),
.B(n_914),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_931),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_937),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_986),
.A2(n_919),
.B(n_936),
.Y(n_1088)
);

AO31x2_ASAP7_75t_L g1089 ( 
.A1(n_952),
.A2(n_966),
.A3(n_1013),
.B(n_1008),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_934),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_947),
.A2(n_906),
.B(n_973),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_938),
.B(n_954),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_912),
.A2(n_926),
.B(n_910),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1006),
.A2(n_944),
.B(n_982),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_SL g1095 ( 
.A(n_934),
.B(n_943),
.Y(n_1095)
);

AOI221x1_ASAP7_75t_L g1096 ( 
.A1(n_987),
.A2(n_995),
.B1(n_889),
.B2(n_1004),
.C(n_999),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_929),
.B(n_899),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_994),
.A2(n_970),
.A3(n_968),
.B(n_957),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_974),
.A2(n_962),
.B(n_1019),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_SL g1100 ( 
.A(n_934),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_1010),
.B(n_1012),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1005),
.B(n_963),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_992),
.A2(n_989),
.B(n_1002),
.C(n_907),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_973),
.A2(n_925),
.B(n_1011),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_922),
.Y(n_1105)
);

AO32x2_ASAP7_75t_L g1106 ( 
.A1(n_995),
.A2(n_958),
.A3(n_985),
.B1(n_990),
.B2(n_953),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_963),
.B(n_984),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_920),
.A2(n_928),
.B(n_973),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_979),
.B(n_984),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_979),
.B(n_984),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_979),
.B(n_992),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_897),
.A2(n_959),
.B1(n_951),
.B2(n_1003),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_897),
.A2(n_960),
.B(n_1003),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_943),
.B(n_960),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_985),
.A2(n_958),
.B(n_960),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_943),
.A2(n_985),
.B(n_958),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_959),
.B(n_951),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_886),
.Y(n_1118)
);

AO21x2_ASAP7_75t_L g1119 ( 
.A1(n_961),
.A2(n_1007),
.B(n_1015),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_885),
.B(n_841),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_885),
.B(n_606),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1015),
.A2(n_895),
.A3(n_896),
.B(n_935),
.Y(n_1122)
);

OAI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_949),
.A2(n_576),
.B(n_752),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_901),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_963),
.B(n_979),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1015),
.A2(n_965),
.B(n_841),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_935),
.A2(n_841),
.B(n_748),
.C(n_909),
.Y(n_1127)
);

BUFx8_ASAP7_75t_SL g1128 ( 
.A(n_890),
.Y(n_1128)
);

AO21x1_ASAP7_75t_L g1129 ( 
.A1(n_896),
.A2(n_841),
.B(n_895),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_885),
.A2(n_558),
.B1(n_834),
.B2(n_833),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_976),
.A2(n_969),
.B(n_950),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_976),
.A2(n_969),
.B(n_950),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_885),
.B(n_841),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_L g1134 ( 
.A(n_941),
.Y(n_1134)
);

BUFx2_ASAP7_75t_SL g1135 ( 
.A(n_890),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_886),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_901),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_929),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_946),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1015),
.A2(n_589),
.B(n_1007),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_885),
.B(n_606),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_917),
.B(n_784),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_885),
.A2(n_748),
.B(n_841),
.C(n_606),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_886),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_885),
.A2(n_748),
.B(n_841),
.C(n_606),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_942),
.B(n_833),
.Y(n_1146)
);

OAI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_887),
.A2(n_834),
.B1(n_833),
.B2(n_858),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_901),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_886),
.Y(n_1149)
);

AOI211x1_ASAP7_75t_L g1150 ( 
.A1(n_949),
.A2(n_585),
.B(n_587),
.C(n_841),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_901),
.Y(n_1151)
);

AOI221x1_ASAP7_75t_L g1152 ( 
.A1(n_1015),
.A2(n_841),
.B1(n_748),
.B2(n_935),
.C(n_896),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_886),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1143),
.A2(n_1145),
.B(n_1123),
.C(n_1120),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1076),
.A2(n_1152),
.B(n_1126),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1046),
.B(n_1052),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1124),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1100),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1129),
.A2(n_1076),
.A3(n_1140),
.B(n_1116),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1032),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_1126),
.A2(n_1140),
.B(n_1033),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1130),
.A2(n_1147),
.B1(n_1133),
.B2(n_1120),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1148),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1035),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1128),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_SL g1166 ( 
.A1(n_1103),
.A2(n_1047),
.B(n_1133),
.C(n_1075),
.Y(n_1166)
);

OAI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1121),
.A2(n_1141),
.B(n_1130),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1150),
.A2(n_1127),
.B1(n_1065),
.B2(n_1050),
.C(n_1056),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1093),
.A2(n_1088),
.B(n_1038),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1072),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1102),
.B(n_1068),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_SL g1172 ( 
.A(n_1134),
.B(n_1097),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1077),
.A2(n_1094),
.B(n_1034),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1023),
.B(n_1042),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1116),
.A2(n_1033),
.A3(n_1045),
.B(n_1096),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1138),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1064),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1118),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1077),
.A2(n_1029),
.B(n_1091),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1023),
.A2(n_1053),
.B1(n_1137),
.B2(n_1024),
.Y(n_1180)
);

CKINVDCx11_ASAP7_75t_R g1181 ( 
.A(n_1067),
.Y(n_1181)
);

CKINVDCx9p33_ASAP7_75t_R g1182 ( 
.A(n_1051),
.Y(n_1182)
);

CKINVDCx6p67_ASAP7_75t_R g1183 ( 
.A(n_1135),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1136),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1144),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1024),
.A2(n_1025),
.B1(n_1055),
.B2(n_1083),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1149),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1153),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1058),
.Y(n_1189)
);

BUFx8_ASAP7_75t_SL g1190 ( 
.A(n_1134),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1074),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1028),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1111),
.B(n_1125),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1117),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1069),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1139),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1049),
.A2(n_1063),
.B(n_1026),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1040),
.A2(n_1060),
.B(n_1080),
.Y(n_1198)
);

BUFx8_ASAP7_75t_SL g1199 ( 
.A(n_1044),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_1112),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1036),
.A2(n_1081),
.A3(n_1025),
.B(n_1055),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1082),
.A2(n_1101),
.B(n_1036),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1082),
.A2(n_1059),
.B(n_1021),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1059),
.A2(n_1042),
.B(n_1119),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1104),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1142),
.A2(n_1151),
.B1(n_1146),
.B2(n_1111),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1078),
.A2(n_1115),
.B(n_1085),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1085),
.A2(n_1061),
.B(n_1071),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1125),
.B(n_1058),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_1054),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1057),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1073),
.A2(n_1071),
.B(n_1066),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1037),
.A2(n_1043),
.B(n_1105),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1086),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1070),
.B(n_1087),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1061),
.A2(n_1066),
.B(n_1099),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1114),
.Y(n_1217)
);

BUFx2_ASAP7_75t_SL g1218 ( 
.A(n_1079),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1020),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1092),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1109),
.B(n_1110),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1020),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1041),
.A2(n_1027),
.B1(n_1031),
.B2(n_1109),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1110),
.B(n_1107),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1113),
.A2(n_1099),
.B(n_1062),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1114),
.A2(n_1022),
.B(n_1106),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1090),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1119),
.A2(n_1021),
.B(n_1062),
.C(n_1122),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1095),
.B(n_1122),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1039),
.A2(n_1089),
.B(n_1084),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1084),
.A2(n_1039),
.B(n_1089),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1098),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1089),
.A2(n_1030),
.B(n_1131),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1098),
.B(n_1124),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1032),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1130),
.A2(n_833),
.B1(n_834),
.B2(n_748),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1111),
.B(n_1125),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1046),
.B(n_1052),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1032),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1134),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1032),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1124),
.B(n_1148),
.Y(n_1242)
);

AO21x2_ASAP7_75t_L g1243 ( 
.A1(n_1076),
.A2(n_1126),
.B(n_1140),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1076),
.A2(n_1152),
.B(n_1126),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1143),
.A2(n_841),
.B(n_769),
.C(n_1145),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1130),
.A2(n_833),
.B1(n_834),
.B2(n_858),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1111),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1124),
.Y(n_1248)
);

OAI22x1_ASAP7_75t_L g1249 ( 
.A1(n_1048),
.A2(n_833),
.B1(n_834),
.B2(n_1121),
.Y(n_1249)
);

AOI221xp5_ASAP7_75t_L g1250 ( 
.A1(n_1130),
.A2(n_585),
.B1(n_587),
.B2(n_576),
.C(n_833),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1121),
.B(n_1141),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1124),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1121),
.B(n_1141),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1121),
.B(n_833),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1138),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1130),
.A2(n_833),
.B1(n_834),
.B2(n_748),
.Y(n_1256)
);

BUFx4_ASAP7_75t_R g1257 ( 
.A(n_1128),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1020),
.B(n_741),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1072),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1051),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1142),
.B(n_609),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1134),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1111),
.B(n_1125),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1138),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1124),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1032),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1121),
.B(n_1141),
.Y(n_1267)
);

CKINVDCx14_ASAP7_75t_R g1268 ( 
.A(n_1138),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1030),
.A2(n_1132),
.B(n_1131),
.Y(n_1269)
);

BUFx4f_ASAP7_75t_SL g1270 ( 
.A(n_1067),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1032),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1076),
.A2(n_1152),
.B(n_1126),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1134),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1030),
.A2(n_1132),
.B(n_1131),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1164),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1217),
.B(n_1193),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1217),
.B(n_1193),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_SL g1278 ( 
.A1(n_1251),
.A2(n_1267),
.B(n_1253),
.Y(n_1278)
);

CKINVDCx14_ASAP7_75t_R g1279 ( 
.A(n_1268),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1171),
.B(n_1156),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1221),
.B(n_1224),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1245),
.A2(n_1154),
.B(n_1249),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1164),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1211),
.B(n_1240),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1209),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1254),
.A2(n_1256),
.B1(n_1236),
.B2(n_1250),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1245),
.A2(n_1154),
.B(n_1186),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1210),
.B(n_1167),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1254),
.A2(n_1246),
.B(n_1168),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1162),
.A2(n_1200),
.B1(n_1211),
.B2(n_1180),
.Y(n_1290)
);

AND2x2_ASAP7_75t_SL g1291 ( 
.A(n_1155),
.B(n_1244),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1238),
.B(n_1215),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1242),
.B(n_1234),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1162),
.B(n_1220),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1262),
.A2(n_1273),
.B(n_1223),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1237),
.B(n_1263),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1237),
.B(n_1263),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1191),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1176),
.Y(n_1299)
);

AND2x4_ASAP7_75t_SL g1300 ( 
.A(n_1183),
.B(n_1157),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1163),
.B(n_1248),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1261),
.A2(n_1228),
.B(n_1206),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1241),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1241),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1209),
.B(n_1192),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1230),
.A2(n_1231),
.B(n_1197),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1270),
.A2(n_1194),
.B1(n_1195),
.B2(n_1252),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1199),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1229),
.A2(n_1244),
.B(n_1155),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1231),
.A2(n_1197),
.B(n_1198),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1160),
.Y(n_1311)
);

NOR2x1_ASAP7_75t_SL g1312 ( 
.A(n_1243),
.B(n_1161),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1265),
.B(n_1192),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1260),
.B(n_1201),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1204),
.A2(n_1202),
.B(n_1213),
.C(n_1166),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1270),
.A2(n_1194),
.B1(n_1195),
.B2(n_1218),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1177),
.A2(n_1185),
.B1(n_1184),
.B2(n_1266),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1178),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1187),
.A2(n_1235),
.B1(n_1271),
.B2(n_1188),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1196),
.B(n_1189),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1196),
.B(n_1214),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1227),
.B(n_1165),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1201),
.B(n_1239),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1189),
.B(n_1247),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1268),
.A2(n_1264),
.B1(n_1176),
.B2(n_1165),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1172),
.A2(n_1226),
.B(n_1225),
.C(n_1272),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1247),
.B(n_1219),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1198),
.A2(n_1202),
.B(n_1173),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1208),
.B(n_1201),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1232),
.A2(n_1207),
.B(n_1216),
.C(n_1205),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1201),
.B(n_1222),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1158),
.A2(n_1203),
.B(n_1212),
.C(n_1219),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1158),
.A2(n_1264),
.B1(n_1222),
.B2(n_1219),
.Y(n_1333)
);

AOI221x1_ASAP7_75t_SL g1334 ( 
.A1(n_1182),
.A2(n_1175),
.B1(n_1255),
.B2(n_1190),
.C(n_1181),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1222),
.B(n_1259),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1170),
.B(n_1259),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1175),
.A2(n_1179),
.B(n_1233),
.C(n_1159),
.Y(n_1337)
);

O2A1O1Ixp5_ASAP7_75t_L g1338 ( 
.A1(n_1170),
.A2(n_1175),
.B(n_1203),
.C(n_1212),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1258),
.B(n_1181),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1233),
.B(n_1169),
.Y(n_1340)
);

CKINVDCx16_ASAP7_75t_R g1341 ( 
.A(n_1274),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1269),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1171),
.B(n_1156),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1254),
.A2(n_833),
.B1(n_834),
.B2(n_858),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1254),
.A2(n_833),
.B1(n_834),
.B2(n_858),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1254),
.A2(n_833),
.B1(n_834),
.B2(n_858),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1174),
.B(n_1251),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1254),
.A2(n_833),
.B1(n_834),
.B2(n_858),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1257),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1221),
.B(n_1224),
.Y(n_1350)
);

INVx4_ASAP7_75t_SL g1351 ( 
.A(n_1201),
.Y(n_1351)
);

OAI31xp33_ASAP7_75t_L g1352 ( 
.A1(n_1167),
.A2(n_987),
.A3(n_1147),
.B(n_1130),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1255),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1336),
.B(n_1335),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1291),
.B(n_1331),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1314),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1336),
.B(n_1335),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1293),
.B(n_1323),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1291),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1286),
.A2(n_1290),
.B1(n_1288),
.B2(n_1294),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1276),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1311),
.B(n_1347),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1352),
.A2(n_1333),
.B1(n_1353),
.B2(n_1277),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1337),
.A2(n_1330),
.B(n_1315),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1329),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1289),
.B(n_1287),
.C(n_1282),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1328),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1351),
.B(n_1309),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1311),
.B(n_1275),
.Y(n_1369)
);

OAI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1334),
.A2(n_1348),
.B1(n_1346),
.B2(n_1344),
.C(n_1345),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1312),
.A2(n_1315),
.B(n_1337),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1283),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1351),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1340),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1318),
.B(n_1298),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1303),
.B(n_1304),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1276),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1281),
.B(n_1350),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1321),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1306),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1326),
.B(n_1301),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1351),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1332),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1313),
.B(n_1302),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1306),
.Y(n_1386)
);

AO22x1_ASAP7_75t_L g1387 ( 
.A1(n_1316),
.A2(n_1349),
.B1(n_1277),
.B2(n_1339),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1310),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1341),
.B(n_1342),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1338),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1328),
.B(n_1305),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1378),
.B(n_1307),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1378),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1366),
.A2(n_1353),
.B1(n_1285),
.B2(n_1279),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1372),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1365),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1365),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1355),
.B(n_1292),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1358),
.B(n_1343),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1358),
.B(n_1280),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1366),
.B(n_1279),
.C(n_1325),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1382),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1367),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1382),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1362),
.B(n_1320),
.Y(n_1405)
);

NOR2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1385),
.B(n_1285),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1356),
.B(n_1324),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1355),
.B(n_1297),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1373),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1372),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1356),
.B(n_1300),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1391),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1391),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1361),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1362),
.B(n_1327),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1371),
.B(n_1295),
.Y(n_1416)
);

INVxp67_ASAP7_75t_R g1417 ( 
.A(n_1368),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1391),
.B(n_1296),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1360),
.A2(n_1296),
.B1(n_1322),
.B2(n_1327),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1388),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1374),
.B(n_1300),
.Y(n_1421)
);

INVx5_ASAP7_75t_L g1422 ( 
.A(n_1368),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1402),
.B(n_1380),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1395),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1412),
.B(n_1384),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1402),
.B(n_1404),
.C(n_1360),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1404),
.A2(n_1385),
.B(n_1370),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1396),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1416),
.A2(n_1370),
.B1(n_1363),
.B2(n_1299),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1401),
.A2(n_1384),
.B1(n_1379),
.B2(n_1284),
.C(n_1371),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1395),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1418),
.B(n_1359),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1421),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1393),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1401),
.B(n_1379),
.C(n_1390),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1405),
.B(n_1380),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1396),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1421),
.Y(n_1438)
);

AOI221xp5_ASAP7_75t_L g1439 ( 
.A1(n_1392),
.A2(n_1387),
.B1(n_1369),
.B2(n_1390),
.C(n_1375),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1399),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1393),
.A2(n_1359),
.B1(n_1361),
.B2(n_1377),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1399),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1416),
.A2(n_1359),
.B1(n_1377),
.B2(n_1361),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1410),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1400),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1416),
.A2(n_1387),
.B1(n_1364),
.B2(n_1359),
.Y(n_1446)
);

AOI31xp33_ASAP7_75t_L g1447 ( 
.A1(n_1394),
.A2(n_1308),
.A3(n_1368),
.B(n_1389),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1416),
.A2(n_1359),
.B1(n_1377),
.B2(n_1373),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1416),
.B(n_1389),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1419),
.A2(n_1357),
.B1(n_1354),
.B2(n_1383),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1414),
.Y(n_1451)
);

INVxp67_ASAP7_75t_SL g1452 ( 
.A(n_1397),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1397),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1403),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1393),
.A2(n_1354),
.B1(n_1357),
.B2(n_1364),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1422),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1420),
.A2(n_1386),
.B(n_1381),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1424),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1456),
.B(n_1413),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_SL g1460 ( 
.A(n_1439),
.B(n_1411),
.C(n_1409),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1424),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1428),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1437),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1457),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1431),
.Y(n_1465)
);

NOR2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1411),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1456),
.B(n_1422),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_SL g1468 ( 
.A(n_1427),
.B(n_1409),
.C(n_1415),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1431),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1432),
.B(n_1398),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1457),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1426),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1457),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1432),
.B(n_1398),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1426),
.B(n_1415),
.C(n_1369),
.Y(n_1475)
);

INVx4_ASAP7_75t_SL g1476 ( 
.A(n_1429),
.Y(n_1476)
);

OR2x6_ASAP7_75t_L g1477 ( 
.A(n_1449),
.B(n_1406),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1425),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1454),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1425),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1444),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1444),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1423),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1433),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1472),
.B(n_1440),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1472),
.B(n_1442),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1478),
.B(n_1452),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1476),
.B(n_1448),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1478),
.B(n_1480),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1484),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1482),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1466),
.B(n_1445),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1482),
.Y(n_1493)
);

NAND4xp25_ASAP7_75t_L g1494 ( 
.A(n_1460),
.B(n_1435),
.C(n_1430),
.D(n_1446),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1458),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1476),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1484),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1433),
.Y(n_1498)
);

AOI221x1_ASAP7_75t_L g1499 ( 
.A1(n_1460),
.A2(n_1429),
.B1(n_1450),
.B2(n_1436),
.C(n_1405),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1438),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1468),
.A2(n_1447),
.B(n_1455),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1458),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1477),
.B(n_1438),
.Y(n_1503)
);

NAND4xp25_ASAP7_75t_L g1504 ( 
.A(n_1468),
.B(n_1434),
.C(n_1441),
.D(n_1278),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1483),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1480),
.B(n_1453),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1483),
.B(n_1400),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1464),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1462),
.B(n_1463),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1477),
.B(n_1417),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1477),
.B(n_1417),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1477),
.B(n_1466),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1464),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1464),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1475),
.B(n_1408),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1458),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1475),
.B(n_1408),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1464),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1470),
.B(n_1474),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1461),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1461),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1476),
.B(n_1443),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1477),
.B(n_1434),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1476),
.Y(n_1524)
);

NAND4xp25_ASAP7_75t_L g1525 ( 
.A(n_1476),
.B(n_1375),
.C(n_1376),
.D(n_1407),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1477),
.B(n_1449),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1470),
.B(n_1474),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1495),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1527),
.B(n_1467),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

NOR2x1_ASAP7_75t_R g1531 ( 
.A(n_1496),
.B(n_1476),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1509),
.B(n_1462),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1527),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1490),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1505),
.B(n_1470),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1495),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1524),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1502),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

AOI32xp33_ASAP7_75t_L g1540 ( 
.A1(n_1496),
.A2(n_1524),
.A3(n_1488),
.B1(n_1522),
.B2(n_1512),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1494),
.A2(n_1476),
.B1(n_1406),
.B2(n_1449),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1516),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1524),
.B(n_1467),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1516),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1520),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1525),
.B(n_1463),
.Y(n_1547)
);

OAI21xp33_ASAP7_75t_L g1548 ( 
.A1(n_1494),
.A2(n_1449),
.B(n_1459),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1515),
.B(n_1459),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1520),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1467),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1521),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1510),
.B(n_1467),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1491),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1451),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1510),
.B(n_1467),
.Y(n_1558)
);

NOR2x1_ASAP7_75t_SL g1559 ( 
.A(n_1489),
.B(n_1422),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1489),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1500),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1491),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1547),
.A2(n_1517),
.B1(n_1486),
.B2(n_1485),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1534),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1560),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1538),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1538),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1561),
.B(n_1499),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1545),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1561),
.B(n_1499),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1523),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1519),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1545),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1557),
.A2(n_1504),
.B1(n_1525),
.B2(n_1523),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1557),
.A2(n_1504),
.B1(n_1364),
.B2(n_1526),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1548),
.A2(n_1511),
.B1(n_1526),
.B2(n_1503),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1560),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1528),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1536),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1507),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1537),
.B(n_1487),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1537),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1541),
.A2(n_1511),
.B1(n_1422),
.B2(n_1449),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1568),
.Y(n_1589)
);

O2A1O1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1573),
.A2(n_1556),
.B(n_1562),
.C(n_1532),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1577),
.A2(n_1551),
.B1(n_1543),
.B2(n_1555),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1564),
.B(n_1533),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1533),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1580),
.B(n_1535),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1578),
.A2(n_1531),
.B(n_1487),
.C(n_1549),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1586),
.B(n_1544),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1568),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1586),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1585),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1567),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1570),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1574),
.B(n_1543),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1574),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1585),
.B(n_1551),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1581),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1600),
.B(n_1594),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1592),
.B(n_1584),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1604),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1604),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1603),
.B(n_1579),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1603),
.B(n_1605),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1598),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1606),
.A2(n_1578),
.B1(n_1563),
.B2(n_1587),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1589),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1615),
.A2(n_1588),
.B1(n_1596),
.B2(n_1593),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1607),
.A2(n_1588),
.B(n_1595),
.C(n_1590),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1609),
.A2(n_1595),
.B(n_1610),
.C(n_1597),
.Y(n_1620)
);

OAI211xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1616),
.A2(n_1613),
.B(n_1608),
.C(n_1591),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1612),
.A2(n_1602),
.B1(n_1601),
.B2(n_1599),
.C(n_1583),
.Y(n_1622)
);

AO21x1_ASAP7_75t_L g1623 ( 
.A1(n_1617),
.A2(n_1576),
.B(n_1572),
.Y(n_1623)
);

AND3x1_ASAP7_75t_L g1624 ( 
.A(n_1611),
.B(n_1582),
.C(n_1571),
.Y(n_1624)
);

NOR2x1_ASAP7_75t_L g1625 ( 
.A(n_1614),
.B(n_1562),
.Y(n_1625)
);

HAxp5_ASAP7_75t_SL g1626 ( 
.A(n_1609),
.B(n_1542),
.CON(n_1626),
.SN(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1610),
.A2(n_1559),
.B(n_1552),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_L g1628 ( 
.A(n_1607),
.B(n_1558),
.C(n_1555),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1618),
.B(n_1506),
.Y(n_1629)
);

OAI32xp33_ASAP7_75t_L g1630 ( 
.A1(n_1626),
.A2(n_1558),
.A3(n_1554),
.B1(n_1550),
.B2(n_1546),
.Y(n_1630)
);

AOI21xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1619),
.A2(n_1506),
.B(n_1493),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1624),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1625),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1633),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1629),
.B(n_1628),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1632),
.A2(n_1621),
.B1(n_1623),
.B2(n_1622),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1631),
.B(n_1529),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1630),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1629),
.Y(n_1639)
);

INVx3_ASAP7_75t_SL g1640 ( 
.A(n_1639),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1634),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1637),
.B(n_1620),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1635),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1638),
.B(n_1493),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1640),
.A2(n_1636),
.B1(n_1627),
.B2(n_1529),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1642),
.B(n_1636),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1643),
.B(n_1641),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1646),
.B(n_1644),
.Y(n_1648)
);

AOI322xp5_ASAP7_75t_L g1649 ( 
.A1(n_1648),
.A2(n_1645),
.A3(n_1647),
.B1(n_1514),
.B2(n_1518),
.C1(n_1508),
.C2(n_1513),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1649),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1518),
.B(n_1514),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1651),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1652),
.A2(n_1559),
.B1(n_1513),
.B2(n_1508),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1653),
.A2(n_1498),
.B1(n_1467),
.B2(n_1479),
.Y(n_1654)
);

OAI21xp33_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1479),
.B(n_1459),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_SL g1656 ( 
.A1(n_1655),
.A2(n_1479),
.B1(n_1471),
.B2(n_1473),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1473),
.B1(n_1471),
.B2(n_1481),
.C(n_1465),
.Y(n_1657)
);

AOI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1473),
.B(n_1471),
.C(n_1469),
.Y(n_1658)
);


endmodule