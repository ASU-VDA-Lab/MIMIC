module real_jpeg_1957_n_17 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_106, n_11, n_14, n_110, n_7, n_3, n_5, n_4, n_102, n_105, n_109, n_101, n_1, n_16, n_15, n_13, n_103, n_17);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_106;
input n_11;
input n_14;
input n_110;
input n_7;
input n_3;
input n_5;
input n_4;
input n_102;
input n_105;
input n_109;
input n_101;
input n_1;
input n_16;
input n_15;
input n_13;
input n_103;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.C(n_53),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_3),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_3),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_4),
.Y(n_84)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_7),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_34),
.B1(n_68),
.B2(n_71),
.Y(n_33)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_9),
.A2(n_43),
.B(n_47),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_20),
.B1(n_21),
.B2(n_26),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_30),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_39),
.B1(n_41),
.B2(n_52),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.C(n_60),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_15),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_27),
.B1(n_98),
.B2(n_99),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_87),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_40),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_25),
.Y(n_55)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_27),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI221xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_74),
.C(n_88),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_64),
.C(n_65),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_56),
.C(n_57),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_51),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_82),
.Y(n_81)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_83),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_89),
.A3(n_90),
.B1(n_93),
.B2(n_94),
.C1(n_97),
.C2(n_111),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.C(n_80),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_101),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_102),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_103),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_104),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_105),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_106),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_107),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_108),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_109),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_110),
.Y(n_87)
);


endmodule