module fake_netlist_6_2597_n_925 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_925);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_925;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_465;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_742;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_608;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_527;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_663;
wire n_361;
wire n_508;
wire n_856;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_122),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_70),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_17),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_93),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_11),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_97),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

BUFx8_ASAP7_75t_SL g191 ( 
.A(n_90),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_126),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_133),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_13),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_14),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_23),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_59),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_2),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_54),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_9),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_89),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_87),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_114),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_50),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_33),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_74),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_134),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_77),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_91),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_82),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_125),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_115),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_16),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_103),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_143),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_49),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_29),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_104),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_7),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_51),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_17),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_28),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_76),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_118),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_150),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_3),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_138),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_81),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_78),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_53),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_99),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_135),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_38),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_5),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_111),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_139),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_130),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_0),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_174),
.B(n_0),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_176),
.B(n_1),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_176),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_224),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_190),
.B(n_1),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_169),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_196),
.B(n_2),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_190),
.B(n_3),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_196),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_230),
.B(n_215),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_215),
.B(n_4),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_36),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_4),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_179),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_181),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_5),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_185),
.B(n_37),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_200),
.B(n_40),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_172),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_177),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_214),
.B(n_41),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_6),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_228),
.B(n_7),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_42),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_191),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_170),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_194),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_43),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_201),
.B(n_8),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_171),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_173),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_203),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_187),
.B(n_44),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_205),
.B1(n_193),
.B2(n_219),
.Y(n_312)
);

AO22x2_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_259),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_195),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_205),
.B1(n_193),
.B2(n_238),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_175),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_178),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_262),
.A2(n_210),
.B1(n_225),
.B2(n_232),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_264),
.A2(n_261),
.B1(n_311),
.B2(n_272),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g324 ( 
.A1(n_294),
.A2(n_195),
.B1(n_184),
.B2(n_237),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_250),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_180),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_268),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_270),
.A2(n_257),
.B1(n_256),
.B2(n_255),
.Y(n_329)
);

AO22x2_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_182),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g333 ( 
.A1(n_267),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_294),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_284),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_183),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_253),
.B1(n_252),
.B2(n_251),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_259),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g342 ( 
.A1(n_267),
.A2(n_274),
.B1(n_292),
.B2(n_306),
.Y(n_342)
);

OA22x2_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_247),
.B1(n_245),
.B2(n_242),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_285),
.A2(n_241),
.B1(n_240),
.B2(n_236),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_310),
.A2(n_235),
.B1(n_233),
.B2(n_229),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_261),
.A2(n_311),
.B1(n_272),
.B2(n_307),
.Y(n_347)
);

OR2x6_ASAP7_75t_L g348 ( 
.A(n_279),
.B(n_20),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_288),
.A2(n_227),
.B1(n_223),
.B2(n_222),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

OR2x6_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_21),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_188),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_300),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_305),
.A2(n_221),
.B1(n_220),
.B2(n_217),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_189),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_21),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_276),
.A2(n_216),
.B1(n_212),
.B2(n_211),
.Y(n_358)
);

AO22x2_ASAP7_75t_L g359 ( 
.A1(n_274),
.A2(n_290),
.B1(n_306),
.B2(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_260),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_308),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_308),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_192),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_22),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_300),
.B(n_197),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_280),
.A2(n_209),
.B1(n_208),
.B2(n_207),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_298),
.B(n_199),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_336),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_308),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_314),
.Y(n_371)
);

INVx4_ASAP7_75t_SL g372 ( 
.A(n_362),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_292),
.B(n_290),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_319),
.A2(n_301),
.B(n_290),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_308),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_365),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_308),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_343),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_312),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_363),
.A2(n_306),
.B(n_301),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_317),
.B(n_300),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_339),
.B(n_301),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_357),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_277),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_322),
.B(n_277),
.Y(n_403)
);

INVx4_ASAP7_75t_SL g404 ( 
.A(n_351),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_316),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_299),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_304),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_343),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_342),
.Y(n_410)
);

BUFx8_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_358),
.B(n_202),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_313),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_303),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_346),
.B(n_304),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_313),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_324),
.B(n_206),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_348),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_318),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_318),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_366),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_353),
.B(n_45),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_320),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_346),
.B(n_358),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_321),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_304),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_327),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_367),
.A2(n_297),
.B(n_271),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_333),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_333),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_303),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_373),
.B(n_304),
.Y(n_448)
);

AO21x1_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_349),
.B(n_345),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_263),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_380),
.B(n_392),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_304),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_415),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_381),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_369),
.B(n_263),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_370),
.B(n_297),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_405),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_297),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_297),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_376),
.B(n_417),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_297),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_273),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_413),
.B(n_297),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_402),
.B(n_265),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_405),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_438),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_375),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_429),
.B(n_284),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_297),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_377),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_396),
.B(n_286),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_348),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_406),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_439),
.B(n_286),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_401),
.B(n_347),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_382),
.B(n_286),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

AND2x2_ASAP7_75t_SL g490 ( 
.A(n_432),
.B(n_323),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_273),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_391),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_389),
.B(n_275),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_421),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_409),
.B(n_275),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_421),
.B(n_286),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_421),
.B(n_286),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_414),
.B(n_281),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_383),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_407),
.B(n_258),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_432),
.A2(n_296),
.B(n_265),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_384),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_348),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_414),
.B(n_281),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_284),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_407),
.B(n_287),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_442),
.B(n_269),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_385),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_443),
.B(n_269),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_393),
.B(n_291),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_386),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_404),
.B(n_291),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_420),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_404),
.B(n_296),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_372),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_404),
.B(n_293),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_423),
.B(n_426),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_427),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_418),
.B(n_287),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_436),
.A2(n_293),
.B1(n_287),
.B2(n_289),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_428),
.B(n_293),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_387),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_433),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_434),
.B(n_46),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_388),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_492),
.B(n_411),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_452),
.B(n_418),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_455),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_456),
.B(n_425),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_447),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_455),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_494),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_456),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_504),
.A2(n_436),
.B(n_412),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_491),
.B(n_412),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_518),
.B(n_260),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_522),
.B(n_460),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_485),
.B(n_391),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_474),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_476),
.B(n_411),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_518),
.Y(n_552)
);

CKINVDCx8_ASAP7_75t_R g553 ( 
.A(n_459),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_518),
.B(n_260),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_476),
.B(n_372),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_454),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_422),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_491),
.B(n_372),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_518),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_522),
.B(n_467),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_422),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_526),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_522),
.B(n_287),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_502),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_494),
.B(n_260),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_475),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_467),
.B(n_430),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_454),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_475),
.B(n_47),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_450),
.B(n_287),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_528),
.B(n_289),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_460),
.B(n_258),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_490),
.B(n_22),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_514),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_289),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_494),
.B(n_260),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_450),
.B(n_23),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_475),
.B(n_48),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_489),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_514),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_473),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_489),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_489),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_514),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_513),
.B(n_293),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_493),
.Y(n_595)
);

NAND2x1_ASAP7_75t_L g596 ( 
.A(n_493),
.B(n_289),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_513),
.B(n_293),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_536),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

BUFx5_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_534),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_560),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_533),
.B(n_460),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_580),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_543),
.A2(n_490),
.B1(n_449),
.B2(n_504),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_560),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_570),
.B(n_547),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_553),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_544),
.B(n_460),
.Y(n_615)
);

NAND2x1p5_ASAP7_75t_L g616 ( 
.A(n_552),
.B(n_528),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_537),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_562),
.B(n_490),
.Y(n_618)
);

NOR2x1_ASAP7_75t_SL g619 ( 
.A(n_552),
.B(n_519),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_595),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_570),
.B(n_547),
.Y(n_621)
);

BUFx24_ASAP7_75t_L g622 ( 
.A(n_556),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_587),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_558),
.Y(n_625)
);

INVx8_ASAP7_75t_L g626 ( 
.A(n_572),
.Y(n_626)
);

INVx6_ASAP7_75t_SL g627 ( 
.A(n_575),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_585),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_585),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_565),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_592),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_553),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_542),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_585),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_585),
.Y(n_635)
);

CKINVDCx8_ASAP7_75t_R g636 ( 
.A(n_562),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_583),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_537),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_544),
.Y(n_640)
);

CKINVDCx11_ASAP7_75t_R g641 ( 
.A(n_588),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_592),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_572),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

BUFx2_ASAP7_75t_SL g645 ( 
.A(n_584),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_584),
.B(n_475),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_584),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_579),
.B(n_524),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_567),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_561),
.B(n_528),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_588),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

BUFx12f_ASAP7_75t_L g655 ( 
.A(n_588),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_636),
.A2(n_579),
.B1(n_530),
.B2(n_576),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_625),
.A2(n_564),
.B1(n_506),
.B2(n_569),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_620),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_648),
.A2(n_446),
.B1(n_484),
.B2(n_464),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_653),
.Y(n_661)
);

OAI21xp33_ASAP7_75t_L g662 ( 
.A1(n_618),
.A2(n_610),
.B(n_648),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_637),
.B(n_464),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_632),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_602),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_618),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_608),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_640),
.A2(n_569),
.B1(n_589),
.B2(n_567),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_623),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_654),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_606),
.B(n_446),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_603),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_610),
.A2(n_621),
.B1(n_612),
.B2(n_449),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_624),
.Y(n_674)
);

CKINVDCx14_ASAP7_75t_R g675 ( 
.A(n_633),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_617),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_630),
.Y(n_677)
);

BUFx12f_ASAP7_75t_L g678 ( 
.A(n_641),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_646),
.A2(n_484),
.B1(n_469),
.B2(n_589),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_600),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_643),
.A2(n_546),
.B1(n_581),
.B2(n_575),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_645),
.A2(n_546),
.B1(n_581),
.B2(n_575),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_599),
.Y(n_683)
);

CKINVDCx6p67_ASAP7_75t_R g684 ( 
.A(n_613),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_631),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_607),
.Y(n_686)
);

CKINVDCx6p67_ASAP7_75t_R g687 ( 
.A(n_641),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_609),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_655),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_622),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_642),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_606),
.B(n_573),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_SL g693 ( 
.A1(n_615),
.A2(n_484),
.B1(n_516),
.B2(n_502),
.Y(n_693)
);

BUFx2_ASAP7_75t_SL g694 ( 
.A(n_600),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_638),
.A2(n_581),
.B1(n_575),
.B2(n_559),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_600),
.Y(n_696)
);

CKINVDCx11_ASAP7_75t_R g697 ( 
.A(n_598),
.Y(n_697)
);

INVx8_ASAP7_75t_L g698 ( 
.A(n_598),
.Y(n_698)
);

CKINVDCx11_ASAP7_75t_R g699 ( 
.A(n_598),
.Y(n_699)
);

BUFx12f_ASAP7_75t_L g700 ( 
.A(n_628),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_646),
.A2(n_484),
.B1(n_473),
.B2(n_497),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_651),
.A2(n_497),
.B1(n_495),
.B2(n_516),
.Y(n_702)
);

CKINVDCx11_ASAP7_75t_R g703 ( 
.A(n_650),
.Y(n_703)
);

OAI22x1_ASAP7_75t_L g704 ( 
.A1(n_651),
.A2(n_521),
.B1(n_563),
.B2(n_548),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_626),
.A2(n_507),
.B1(n_500),
.B2(n_509),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_SL g706 ( 
.A1(n_615),
.A2(n_507),
.B(n_500),
.Y(n_706)
);

CKINVDCx8_ASAP7_75t_R g707 ( 
.A(n_629),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_661),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_662),
.A2(n_647),
.B1(n_457),
.B2(n_626),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_SL g710 ( 
.A1(n_660),
.A2(n_662),
.B(n_656),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_673),
.A2(n_457),
.B1(n_626),
.B2(n_590),
.Y(n_711)
);

OAI222xp33_ASAP7_75t_L g712 ( 
.A1(n_705),
.A2(n_581),
.B1(n_523),
.B2(n_616),
.C1(n_566),
.C2(n_586),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_666),
.A2(n_594),
.B1(n_591),
.B2(n_571),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_665),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_SL g715 ( 
.A1(n_693),
.A2(n_619),
.B1(n_622),
.B2(n_616),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_702),
.A2(n_495),
.B(n_516),
.Y(n_716)
);

INVxp33_ASAP7_75t_SL g717 ( 
.A(n_686),
.Y(n_717)
);

CKINVDCx6p67_ASAP7_75t_R g718 ( 
.A(n_664),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_666),
.A2(n_557),
.B1(n_571),
.B2(n_574),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_683),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_663),
.B(n_510),
.Y(n_721)
);

BUFx5_ASAP7_75t_L g722 ( 
.A(n_667),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_706),
.A2(n_540),
.B1(n_600),
.B2(n_496),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_669),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_SL g725 ( 
.A1(n_706),
.A2(n_523),
.B(n_448),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_671),
.A2(n_574),
.B1(n_578),
.B2(n_525),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_693),
.A2(n_614),
.B1(n_629),
.B2(n_635),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_657),
.A2(n_701),
.B1(n_679),
.B2(n_681),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_676),
.B(n_510),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_690),
.A2(n_614),
.B1(n_635),
.B2(n_629),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_678),
.A2(n_614),
.B1(n_652),
.B2(n_629),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_692),
.A2(n_578),
.B1(n_525),
.B2(n_529),
.Y(n_732)
);

BUFx4f_ASAP7_75t_SL g733 ( 
.A(n_687),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_704),
.A2(n_529),
.B1(n_482),
.B2(n_511),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_707),
.A2(n_668),
.B1(n_684),
.B2(n_672),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_658),
.Y(n_736)
);

AOI222xp33_ASAP7_75t_L g737 ( 
.A1(n_703),
.A2(n_508),
.B1(n_520),
.B2(n_527),
.C1(n_512),
.C2(n_539),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_670),
.Y(n_738)
);

BUFx8_ASAP7_75t_SL g739 ( 
.A(n_688),
.Y(n_739)
);

OAI21xp33_ASAP7_75t_L g740 ( 
.A1(n_675),
.A2(n_486),
.B(n_529),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_674),
.A2(n_482),
.B1(n_511),
.B2(n_508),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_685),
.A2(n_535),
.B1(n_627),
.B2(n_470),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_677),
.A2(n_627),
.B1(n_614),
.B2(n_652),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_682),
.A2(n_652),
.B1(n_635),
.B2(n_617),
.Y(n_744)
);

OAI222xp33_ASAP7_75t_L g745 ( 
.A1(n_691),
.A2(n_503),
.B1(n_471),
.B2(n_649),
.C1(n_639),
.C2(n_593),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_SL g746 ( 
.A1(n_677),
.A2(n_652),
.B1(n_635),
.B2(n_601),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_659),
.Y(n_747)
);

INVx4_ASAP7_75t_R g748 ( 
.A(n_697),
.Y(n_748)
);

AOI21xp33_ASAP7_75t_L g749 ( 
.A1(n_695),
.A2(n_597),
.B(n_483),
.Y(n_749)
);

INVxp33_ASAP7_75t_L g750 ( 
.A(n_689),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_694),
.A2(n_601),
.B1(n_604),
.B2(n_605),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_689),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_689),
.B(n_604),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_699),
.A2(n_478),
.B1(n_519),
.B2(n_501),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_698),
.A2(n_478),
.B1(n_505),
.B2(n_501),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_700),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_698),
.B(n_512),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_698),
.A2(n_472),
.B1(n_479),
.B2(n_470),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_659),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_659),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_680),
.B(n_520),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_680),
.A2(n_458),
.B(n_498),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_696),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_696),
.Y(n_764)
);

BUFx12f_ASAP7_75t_L g765 ( 
.A(n_703),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_658),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_662),
.A2(n_472),
.B1(n_479),
.B2(n_470),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_683),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_710),
.A2(n_639),
.B1(n_521),
.B2(n_471),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_728),
.A2(n_465),
.B1(n_472),
.B2(n_479),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_715),
.A2(n_471),
.B1(n_644),
.B2(n_634),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_720),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_736),
.B(n_649),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_SL g774 ( 
.A1(n_723),
.A2(n_605),
.B(n_604),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_711),
.A2(n_737),
.B1(n_716),
.B2(n_740),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_721),
.B(n_628),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_709),
.A2(n_601),
.B1(n_465),
.B2(n_501),
.Y(n_777)
);

OAI222xp33_ASAP7_75t_L g778 ( 
.A1(n_709),
.A2(n_596),
.B1(n_465),
.B2(n_505),
.C1(n_541),
.C2(n_549),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_727),
.A2(n_644),
.B1(n_634),
.B2(n_628),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_SL g780 ( 
.A1(n_735),
.A2(n_601),
.B1(n_605),
.B2(n_628),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_SL g781 ( 
.A1(n_744),
.A2(n_601),
.B1(n_605),
.B2(n_634),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_733),
.A2(n_765),
.B1(n_730),
.B2(n_717),
.Y(n_782)
);

OAI222xp33_ASAP7_75t_L g783 ( 
.A1(n_711),
.A2(n_505),
.B1(n_541),
.B2(n_531),
.C1(n_554),
.C2(n_538),
.Y(n_783)
);

OAI222xp33_ASAP7_75t_L g784 ( 
.A1(n_742),
.A2(n_754),
.B1(n_741),
.B2(n_729),
.C1(n_746),
.C2(n_734),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_733),
.A2(n_761),
.B1(n_757),
.B2(n_734),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_752),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_708),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_725),
.B(n_517),
.C(n_515),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_742),
.A2(n_601),
.B1(n_644),
.B2(n_634),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_719),
.A2(n_644),
.B1(n_611),
.B2(n_463),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_756),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_741),
.A2(n_554),
.B1(n_549),
.B2(n_538),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_732),
.A2(n_532),
.B1(n_531),
.B2(n_460),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_732),
.A2(n_532),
.B1(n_460),
.B2(n_488),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_714),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_738),
.B(n_499),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_726),
.A2(n_724),
.B1(n_766),
.B2(n_767),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_726),
.B(n_460),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_722),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_748),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_718),
.A2(n_515),
.B1(n_517),
.B2(n_480),
.Y(n_801)
);

OAI222xp33_ASAP7_75t_L g802 ( 
.A1(n_719),
.A2(n_582),
.B1(n_568),
.B2(n_611),
.C1(n_468),
.C2(n_466),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_767),
.A2(n_460),
.B1(n_480),
.B2(n_466),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_743),
.A2(n_480),
.B1(n_460),
.B2(n_466),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_722),
.A2(n_480),
.B1(n_453),
.B2(n_466),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_722),
.B(n_568),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_722),
.A2(n_468),
.B1(n_461),
.B2(n_582),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_713),
.A2(n_577),
.B1(n_555),
.B2(n_545),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_722),
.A2(n_468),
.B1(n_461),
.B2(n_477),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_722),
.A2(n_468),
.B1(n_461),
.B2(n_477),
.Y(n_810)
);

OAI222xp33_ASAP7_75t_L g811 ( 
.A1(n_713),
.A2(n_461),
.B1(n_25),
.B2(n_26),
.C1(n_27),
.C2(n_28),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_749),
.A2(n_477),
.B1(n_577),
.B2(n_545),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_750),
.A2(n_477),
.B1(n_555),
.B2(n_266),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_758),
.A2(n_266),
.B1(n_25),
.B2(n_27),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_753),
.B(n_24),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_755),
.A2(n_266),
.B1(n_258),
.B2(n_30),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_758),
.A2(n_266),
.B1(n_258),
.B2(n_30),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_772),
.B(n_773),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_788),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_791),
.B(n_739),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_775),
.A2(n_731),
.B1(n_751),
.B2(n_759),
.Y(n_821)
);

NAND3xp33_ASAP7_75t_L g822 ( 
.A(n_775),
.B(n_747),
.C(n_760),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_787),
.B(n_24),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_795),
.B(n_29),
.Y(n_824)
);

OAI221xp5_ASAP7_75t_L g825 ( 
.A1(n_785),
.A2(n_712),
.B1(n_32),
.B2(n_33),
.C(n_34),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_799),
.B(n_31),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_776),
.B(n_31),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_797),
.B(n_32),
.Y(n_828)
);

AOI21xp33_ASAP7_75t_L g829 ( 
.A1(n_769),
.A2(n_745),
.B(n_55),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_797),
.B(n_52),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_814),
.A2(n_266),
.B1(n_258),
.B2(n_60),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_796),
.B(n_56),
.Y(n_832)
);

OAI221xp5_ASAP7_75t_SL g833 ( 
.A1(n_814),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_780),
.B(n_64),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_806),
.B(n_65),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_791),
.B(n_66),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_816),
.A2(n_67),
.B(n_68),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_811),
.B(n_69),
.C(n_71),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_815),
.B(n_73),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_782),
.A2(n_258),
.B1(n_75),
.B2(n_79),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_781),
.B(n_80),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_777),
.B(n_83),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_770),
.B(n_85),
.Y(n_843)
);

NAND4xp25_ASAP7_75t_L g844 ( 
.A(n_786),
.B(n_94),
.C(n_95),
.D(n_96),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_SL g845 ( 
.A1(n_784),
.A2(n_98),
.B(n_100),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_798),
.B(n_101),
.Y(n_846)
);

OAI221xp5_ASAP7_75t_L g847 ( 
.A1(n_801),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.C(n_107),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_804),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_812),
.B(n_113),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_771),
.B(n_116),
.C(n_119),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_789),
.B(n_794),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_822),
.B(n_800),
.Y(n_852)
);

AO21x2_ASAP7_75t_L g853 ( 
.A1(n_829),
.A2(n_774),
.B(n_779),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_826),
.Y(n_854)
);

OA211x2_ASAP7_75t_L g855 ( 
.A1(n_837),
.A2(n_805),
.B(n_794),
.C(n_793),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_845),
.B(n_822),
.C(n_838),
.Y(n_856)
);

AO21x2_ASAP7_75t_L g857 ( 
.A1(n_850),
.A2(n_802),
.B(n_778),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_818),
.B(n_826),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_827),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_833),
.B(n_819),
.C(n_837),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_827),
.B(n_813),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_L g862 ( 
.A(n_828),
.B(n_817),
.C(n_810),
.Y(n_862)
);

XNOR2xp5_ASAP7_75t_L g863 ( 
.A(n_844),
.B(n_790),
.Y(n_863)
);

OAI211xp5_ASAP7_75t_SL g864 ( 
.A1(n_823),
.A2(n_807),
.B(n_809),
.C(n_793),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_828),
.B(n_825),
.C(n_830),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_841),
.B(n_803),
.Y(n_866)
);

NOR2x1_ASAP7_75t_L g867 ( 
.A(n_824),
.B(n_783),
.Y(n_867)
);

AO21x2_ASAP7_75t_L g868 ( 
.A1(n_846),
.A2(n_808),
.B(n_792),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_839),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_835),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_851),
.B(n_821),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_835),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_831),
.B(n_803),
.C(n_792),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_854),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_858),
.B(n_841),
.Y(n_875)
);

NAND4xp75_ASAP7_75t_SL g876 ( 
.A(n_866),
.B(n_834),
.C(n_836),
.D(n_820),
.Y(n_876)
);

NOR2x1_ASAP7_75t_L g877 ( 
.A(n_852),
.B(n_832),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_858),
.B(n_834),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_854),
.Y(n_879)
);

NAND4xp75_ASAP7_75t_L g880 ( 
.A(n_855),
.B(n_849),
.C(n_842),
.D(n_843),
.Y(n_880)
);

NAND4xp75_ASAP7_75t_SL g881 ( 
.A(n_866),
.B(n_849),
.C(n_842),
.D(n_847),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_872),
.Y(n_882)
);

XOR2xp5_ASAP7_75t_L g883 ( 
.A(n_871),
.B(n_840),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_859),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_859),
.B(n_848),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_870),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_870),
.Y(n_887)
);

AO22x1_ASAP7_75t_L g888 ( 
.A1(n_877),
.A2(n_867),
.B1(n_869),
.B2(n_861),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_886),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_883),
.B(n_856),
.Y(n_890)
);

XOR2x2_ASAP7_75t_L g891 ( 
.A(n_883),
.B(n_860),
.Y(n_891)
);

XOR2x2_ASAP7_75t_L g892 ( 
.A(n_876),
.B(n_856),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_882),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_884),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_890),
.A2(n_880),
.B1(n_865),
.B2(n_863),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_893),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_890),
.A2(n_880),
.B1(n_865),
.B2(n_863),
.Y(n_897)
);

OA22x2_ASAP7_75t_L g898 ( 
.A1(n_894),
.A2(n_879),
.B1(n_874),
.B2(n_887),
.Y(n_898)
);

XNOR2x1_ASAP7_75t_L g899 ( 
.A(n_891),
.B(n_881),
.Y(n_899)
);

XNOR2x2_ASAP7_75t_L g900 ( 
.A(n_892),
.B(n_867),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_894),
.A2(n_878),
.B1(n_862),
.B2(n_855),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_898),
.Y(n_902)
);

XOR2xp5_ASAP7_75t_L g903 ( 
.A(n_899),
.B(n_862),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_900),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_903),
.A2(n_897),
.B1(n_895),
.B2(n_901),
.Y(n_905)
);

OAI322xp33_ASAP7_75t_L g906 ( 
.A1(n_904),
.A2(n_896),
.A3(n_878),
.B1(n_889),
.B2(n_888),
.C1(n_879),
.C2(n_874),
.Y(n_906)
);

AOI221xp5_ASAP7_75t_L g907 ( 
.A1(n_906),
.A2(n_904),
.B1(n_902),
.B2(n_885),
.C(n_875),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_905),
.A2(n_853),
.B1(n_857),
.B2(n_873),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_907),
.A2(n_857),
.B1(n_868),
.B2(n_864),
.Y(n_909)
);

OAI22xp33_ASAP7_75t_L g910 ( 
.A1(n_908),
.A2(n_868),
.B1(n_120),
.B2(n_123),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_909),
.B(n_128),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_910),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_912),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_911),
.B(n_131),
.C(n_132),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_913),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_914),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_916),
.A2(n_140),
.B1(n_142),
.B2(n_144),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_915),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_918),
.Y(n_919)
);

AO22x1_ASAP7_75t_L g920 ( 
.A1(n_919),
.A2(n_917),
.B1(n_146),
.B2(n_147),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_920),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_921),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_922),
.Y(n_923)
);

AOI221xp5_ASAP7_75t_L g924 ( 
.A1(n_923),
.A2(n_153),
.B1(n_157),
.B2(n_158),
.C(n_159),
.Y(n_924)
);

AOI211xp5_ASAP7_75t_L g925 ( 
.A1(n_924),
.A2(n_161),
.B(n_164),
.C(n_165),
.Y(n_925)
);


endmodule