module fake_jpeg_8151_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_43),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_21),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_19),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_52),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_66),
.B(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_34),
.B1(n_21),
.B2(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_45),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_65),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_34),
.B1(n_23),
.B2(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_23),
.B1(n_25),
.B2(n_20),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_32),
.B1(n_25),
.B2(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_62),
.Y(n_100)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_74),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_77),
.B1(n_63),
.B2(n_45),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_41),
.B1(n_35),
.B2(n_28),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_79),
.B1(n_83),
.B2(n_63),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_35),
.B1(n_28),
.B2(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_89),
.B1(n_67),
.B2(n_39),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_33),
.B1(n_20),
.B2(n_24),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_45),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_56),
.C(n_38),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_33),
.B1(n_24),
.B2(n_17),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_102),
.B1(n_104),
.B2(n_109),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx24_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_108),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_84),
.B(n_76),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_100),
.B(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_48),
.B1(n_53),
.B2(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_63),
.B1(n_56),
.B2(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_75),
.B1(n_91),
.B2(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_61),
.B1(n_57),
.B2(n_46),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_114),
.Y(n_119)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_2),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_72),
.B(n_31),
.C(n_4),
.D(n_5),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_127),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_90),
.B1(n_87),
.B2(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_104),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_103),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_136),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_87),
.B1(n_70),
.B2(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_36),
.B1(n_38),
.B2(n_17),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_113),
.B1(n_117),
.B2(n_112),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_36),
.B(n_38),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_118),
.B(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_17),
.B1(n_29),
.B2(n_31),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_74),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_139),
.Y(n_186)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_115),
.B(n_97),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_154),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_114),
.C(n_111),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_147),
.C(n_158),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_130),
.C(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_149),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_164),
.B1(n_131),
.B2(n_118),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_120),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_105),
.B(n_95),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_163),
.B(n_125),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_141),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_97),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_96),
.C(n_101),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_162),
.C(n_157),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_74),
.C(n_86),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_29),
.B(n_3),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_124),
.A2(n_113),
.B1(n_3),
.B2(n_4),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_172),
.Y(n_198)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_182),
.C(n_146),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_177),
.B1(n_185),
.B2(n_159),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_186),
.B(n_143),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_137),
.B1(n_140),
.B2(n_121),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_183),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_153),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_127),
.B1(n_123),
.B2(n_113),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_188),
.C(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_147),
.C(n_162),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_202),
.B(n_203),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_159),
.B1(n_143),
.B2(n_156),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_200),
.B1(n_183),
.B2(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_170),
.B(n_139),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_158),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_161),
.B(n_139),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_212),
.B1(n_190),
.B2(n_203),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_207),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_167),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_216),
.C(n_29),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_173),
.B(n_176),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_202),
.B(n_198),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_180),
.B1(n_174),
.B2(n_173),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_167),
.B(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_191),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_171),
.C(n_86),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_195),
.C(n_189),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_217),
.B(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_221),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_220),
.A2(n_208),
.B(n_227),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_224),
.C(n_225),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_196),
.B(n_86),
.C(n_29),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_2),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_11),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_210),
.C(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_208),
.C(n_206),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_12),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_233),
.C(n_223),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_15),
.Y(n_238)
);

AOI21x1_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_5),
.B(n_7),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_12),
.C(n_16),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_238),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_7),
.B(n_8),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_229),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_232),
.B1(n_8),
.B2(n_10),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_244),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_239),
.B(n_110),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_237),
.CI(n_234),
.CON(n_247),
.SN(n_247)
);

OAI311xp33_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_246),
.A3(n_13),
.B1(n_14),
.C1(n_7),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_250),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_110),
.Y(n_253)
);


endmodule