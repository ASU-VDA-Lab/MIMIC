module real_jpeg_33599_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

INVx2_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_0),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_1),
.B(n_103),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_SL g107 ( 
.A(n_1),
.B(n_108),
.C(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_108),
.C(n_110),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_1),
.B(n_110),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_6),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_6),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_6),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_7),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_8),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_10),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_11),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_11),
.B(n_155),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_11),
.B(n_254),
.Y(n_253)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_12),
.A2(n_13),
.B1(n_127),
.B2(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_13),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_13),
.B(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_13),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_14),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_15),
.B(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_174),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_173),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_19),
.B(n_113),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_98),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_20),
.A2(n_21),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_35),
.B1(n_36),
.B2(n_54),
.Y(n_22)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_23),
.B(n_36),
.C(n_55),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_25),
.B(n_29),
.Y(n_170)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_28),
.Y(n_167)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_28),
.Y(n_258)
);

NOR2x1_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_30),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_30),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_34),
.Y(n_132)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.C(n_48),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_37),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_182)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_41),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_42),
.B(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_56),
.B(n_62),
.C(n_68),
.Y(n_169)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_59),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_68),
.B2(n_71),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx11_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_70),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_73),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_89),
.B2(n_97),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_83),
.B2(n_88),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_97),
.C(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_87),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

XOR2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_91),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_R g98 ( 
.A(n_99),
.B(n_101),
.C(n_107),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_99),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_99),
.B(n_101),
.C(n_107),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_101),
.A2(n_102),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OR2x2_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

XNOR2x2_ASAP7_75t_L g213 ( 
.A(n_108),
.B(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_149),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_147),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_133),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B(n_125),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_139)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_171),
.B2(n_172),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_168),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_165),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_159),
.Y(n_163)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_269),
.B(n_276),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_215),
.B(n_268),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_201),
.C(n_202),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_178),
.A2(n_201),
.B(n_202),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_196),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_197),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_196),
.C(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.C(n_193),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.C(n_213),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_207),
.B1(n_213),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_234),
.B(n_267),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_231),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.C(n_227),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_219),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_222),
.B(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_261),
.B(n_266),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_246),
.B(n_260),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_259),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_259),
.Y(n_265)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_274),
.Y(n_276)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);


endmodule