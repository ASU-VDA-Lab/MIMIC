module fake_jpeg_917_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_68),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_38),
.B1(n_47),
.B2(n_45),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_38),
.B1(n_43),
.B2(n_49),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_42),
.C(n_37),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_75),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_59),
.B1(n_66),
.B2(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_0),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_95),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_43),
.B(n_59),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_84),
.CON(n_107),
.SN(n_107)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_59),
.B(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_48),
.B1(n_1),
.B2(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_9),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_9),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_0),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_35),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_34),
.B(n_18),
.C(n_19),
.D(n_23),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_10),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_21),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_27),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_20),
.B1(n_33),
.B2(n_30),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_121),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_119),
.B(n_103),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_15),
.B(n_28),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_116),
.B1(n_119),
.B2(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_125),
.B1(n_117),
.B2(n_115),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_131),
.B(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_123),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_124),
.C(n_121),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_109),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_118),
.B(n_24),
.Y(n_139)
);


endmodule