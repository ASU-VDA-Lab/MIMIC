module real_aes_11996_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1595;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1584;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI221xp5_ASAP7_75t_L g1612 ( .A1(n_0), .A2(n_41), .B1(n_705), .B2(n_955), .C(n_960), .Y(n_1612) );
OAI22xp33_ASAP7_75t_L g1617 ( .A1(n_0), .A2(n_276), .B1(n_479), .B2(n_1080), .Y(n_1617) );
XNOR2xp5_ASAP7_75t_L g1578 ( .A(n_1), .B(n_1579), .Y(n_1578) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_2), .Y(n_944) );
XNOR2xp5_ASAP7_75t_L g1035 ( .A(n_3), .B(n_1036), .Y(n_1035) );
AO221x1_ASAP7_75t_L g1284 ( .A1(n_3), .A2(n_154), .B1(n_1285), .B2(n_1291), .C(n_1294), .Y(n_1284) );
CKINVDCx5p33_ASAP7_75t_R g1047 ( .A(n_4), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_5), .A2(n_268), .B1(n_651), .B2(n_912), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_5), .A2(n_268), .B1(n_512), .B2(n_527), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_6), .A2(n_240), .B1(n_416), .B2(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g448 ( .A(n_6), .Y(n_448) );
XNOR2xp5_ASAP7_75t_L g984 ( .A(n_7), .B(n_985), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_8), .Y(n_1233) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_9), .Y(n_963) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_10), .Y(n_294) );
INVx1_ASAP7_75t_L g401 ( .A(n_10), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_10), .B(n_206), .Y(n_545) );
AND2x2_ASAP7_75t_L g553 ( .A(n_10), .B(n_400), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_11), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_12), .A2(n_119), .B1(n_1285), .B2(n_1293), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_13), .A2(n_152), .B1(n_512), .B2(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g593 ( .A(n_13), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_14), .A2(n_187), .B1(n_497), .B2(n_506), .Y(n_1058) );
INVx1_ASAP7_75t_L g1076 ( .A(n_14), .Y(n_1076) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_15), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g1011 ( .A1(n_16), .A2(n_94), .B1(n_802), .B2(n_805), .Y(n_1011) );
INVx1_ASAP7_75t_L g1027 ( .A(n_16), .Y(n_1027) );
INVx1_ASAP7_75t_L g338 ( .A(n_17), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_17), .A2(n_74), .B1(n_438), .B2(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g761 ( .A(n_18), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_18), .A2(n_76), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g997 ( .A(n_19), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g1200 ( .A(n_20), .Y(n_1200) );
AO22x2_ASAP7_75t_L g1130 ( .A1(n_21), .A2(n_1131), .B1(n_1132), .B2(n_1182), .Y(n_1130) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_21), .Y(n_1131) );
AO221x2_ASAP7_75t_L g1377 ( .A1(n_21), .A2(n_174), .B1(n_1291), .B2(n_1378), .C(n_1380), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1074 ( .A1(n_22), .A2(n_231), .B1(n_369), .B2(n_955), .C(n_960), .Y(n_1074) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_22), .A2(n_87), .B1(n_802), .B2(n_805), .Y(n_1081) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_23), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g314 ( .A(n_24), .Y(n_314) );
OR2x2_ASAP7_75t_L g475 ( .A(n_24), .B(n_476), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_25), .A2(n_140), .B1(n_472), .B2(n_479), .Y(n_1095) );
INVx1_ASAP7_75t_L g1114 ( .A(n_25), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_26), .A2(n_101), .B1(n_368), .B2(n_372), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_26), .A2(n_101), .B1(n_408), .B2(n_410), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_27), .Y(n_495) );
BUFx2_ASAP7_75t_L g360 ( .A(n_28), .Y(n_360) );
INVx1_ASAP7_75t_L g397 ( .A(n_28), .Y(n_397) );
BUFx2_ASAP7_75t_L g425 ( .A(n_28), .Y(n_425) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_28), .B(n_545), .Y(n_1209) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_29), .A2(n_196), .B1(n_379), .B2(n_642), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_29), .A2(n_196), .B1(n_713), .B2(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g626 ( .A(n_30), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_30), .A2(n_195), .B1(n_640), .B2(n_642), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g1511 ( .A1(n_31), .A2(n_105), .B1(n_523), .B2(n_718), .C(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1541 ( .A(n_31), .Y(n_1541) );
INVx1_ASAP7_75t_L g1055 ( .A(n_32), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_32), .A2(n_72), .B1(n_771), .B2(n_772), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1521 ( .A1(n_33), .A2(n_157), .B1(n_679), .B2(n_1522), .C(n_1524), .Y(n_1521) );
INVx1_ASAP7_75t_L g1552 ( .A(n_33), .Y(n_1552) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_34), .A2(n_103), .B1(n_630), .B2(n_936), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_34), .A2(n_103), .B1(n_705), .B2(n_955), .C(n_956), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_35), .A2(n_60), .B1(n_295), .B2(n_457), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_35), .A2(n_168), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_36), .A2(n_68), .B1(n_1167), .B2(n_1170), .Y(n_1169) );
INVxp67_ASAP7_75t_SL g1175 ( .A(n_36), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_37), .A2(n_232), .B1(n_630), .B2(n_632), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_37), .A2(n_232), .B1(n_647), .B2(n_654), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_38), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_39), .Y(n_945) );
INVx1_ASAP7_75t_L g1073 ( .A(n_40), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g1079 ( .A1(n_40), .A2(n_231), .B1(n_479), .B2(n_1080), .Y(n_1079) );
OAI22xp33_ASAP7_75t_L g1618 ( .A1(n_41), .A2(n_57), .B1(n_802), .B2(n_805), .Y(n_1618) );
INVx1_ASAP7_75t_L g352 ( .A(n_42), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_42), .A2(n_250), .B1(n_389), .B2(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g754 ( .A(n_43), .Y(n_754) );
OAI211xp5_ASAP7_75t_SL g784 ( .A1(n_43), .A2(n_549), .B(n_785), .C(n_795), .Y(n_784) );
INVx1_ASAP7_75t_L g853 ( .A(n_44), .Y(n_853) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_44), .A2(n_78), .B1(n_802), .B2(n_805), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_45), .A2(n_277), .B1(n_491), .B2(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g949 ( .A(n_45), .Y(n_949) );
INVx1_ASAP7_75t_L g1300 ( .A(n_46), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g1515 ( .A(n_47), .Y(n_1515) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_48), .A2(n_234), .B1(n_619), .B2(n_620), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_48), .A2(n_234), .B1(n_665), .B2(n_666), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_49), .A2(n_158), .B1(n_600), .B2(n_602), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_49), .A2(n_158), .B1(n_1125), .B2(n_1127), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_50), .Y(n_746) );
INVx1_ASAP7_75t_L g1090 ( .A(n_51), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g794 ( .A1(n_52), .A2(n_278), .B1(n_374), .B2(n_569), .C(n_705), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g801 ( .A1(n_52), .A2(n_56), .B1(n_802), .B2(n_805), .Y(n_801) );
INVx1_ASAP7_75t_L g1060 ( .A(n_53), .Y(n_1060) );
INVx1_ASAP7_75t_L g485 ( .A(n_54), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_54), .A2(n_58), .B1(n_565), .B2(n_566), .C(n_569), .Y(n_564) );
INVx1_ASAP7_75t_L g826 ( .A(n_55), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_55), .A2(n_64), .B1(n_771), .B2(n_772), .Y(n_831) );
INVx1_ASAP7_75t_L g789 ( .A(n_56), .Y(n_789) );
INVx1_ASAP7_75t_L g1610 ( .A(n_57), .Y(n_1610) );
INVx1_ASAP7_75t_L g477 ( .A(n_58), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g1594 ( .A1(n_59), .A2(n_270), .B1(n_739), .B2(n_1595), .Y(n_1594) );
OAI22xp5_ASAP7_75t_L g1598 ( .A1(n_59), .A2(n_270), .B1(n_600), .B2(n_602), .Y(n_1598) );
OAI22xp33_ASAP7_75t_L g687 ( .A1(n_60), .A2(n_230), .B1(n_688), .B2(n_691), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g1155 ( .A1(n_61), .A2(n_116), .B1(n_374), .B2(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_61), .A2(n_116), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
INVx1_ASAP7_75t_L g793 ( .A(n_62), .Y(n_793) );
OAI22xp33_ASAP7_75t_L g800 ( .A1(n_62), .A2(n_278), .B1(n_472), .B2(n_479), .Y(n_800) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_63), .A2(n_307), .B1(n_459), .B2(n_460), .Y(n_306) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_63), .Y(n_459) );
INVx1_ASAP7_75t_L g825 ( .A(n_64), .Y(n_825) );
AO221x1_ASAP7_75t_L g959 ( .A1(n_65), .A2(n_86), .B1(n_369), .B2(n_655), .C(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g974 ( .A(n_65), .Y(n_974) );
OAI221xp5_ASAP7_75t_L g1099 ( .A1(n_66), .A2(n_578), .B1(n_783), .B2(n_1100), .C(n_1104), .Y(n_1099) );
AOI22xp33_ASAP7_75t_SL g1123 ( .A1(n_66), .A2(n_212), .B1(n_419), .B2(n_718), .Y(n_1123) );
INVx1_ASAP7_75t_L g891 ( .A(n_67), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_67), .A2(n_135), .B1(n_527), .B2(n_923), .Y(n_922) );
INVxp33_ASAP7_75t_L g1181 ( .A(n_68), .Y(n_1181) );
INVx1_ASAP7_75t_L g1193 ( .A(n_69), .Y(n_1193) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_69), .A2(n_134), .B1(n_414), .B2(n_1252), .C(n_1253), .Y(n_1251) );
INVx1_ASAP7_75t_L g1301 ( .A(n_70), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_71), .A2(n_185), .B1(n_1127), .B2(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1539 ( .A(n_71), .Y(n_1539) );
INVx1_ASAP7_75t_L g1056 ( .A(n_72), .Y(n_1056) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_73), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g1160 ( .A1(n_73), .A2(n_108), .B1(n_372), .B2(n_1156), .Y(n_1160) );
INVx1_ASAP7_75t_L g344 ( .A(n_74), .Y(n_344) );
INVx1_ASAP7_75t_L g894 ( .A(n_75), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_75), .A2(n_209), .B1(n_632), .B2(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g758 ( .A(n_76), .Y(n_758) );
INVx1_ASAP7_75t_L g1103 ( .A(n_77), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_77), .A2(n_213), .B1(n_1121), .B2(n_1122), .Y(n_1120) );
INVx1_ASAP7_75t_L g850 ( .A(n_78), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_79), .A2(n_123), .B1(n_685), .B2(n_686), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_79), .A2(n_123), .B1(n_642), .B2(n_651), .Y(n_709) );
INVx1_ASAP7_75t_L g886 ( .A(n_80), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_80), .A2(n_128), .B1(n_640), .B2(n_778), .Y(n_909) );
AO221x1_ASAP7_75t_L g1331 ( .A1(n_81), .A2(n_126), .B1(n_1285), .B2(n_1293), .C(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g682 ( .A(n_82), .Y(n_682) );
OAI222xp33_ASAP7_75t_L g695 ( .A1(n_82), .A2(n_168), .B1(n_188), .B2(n_441), .C1(n_696), .C2(n_697), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_83), .A2(n_118), .B1(n_422), .B2(n_723), .Y(n_1172) );
INVxp33_ASAP7_75t_SL g1178 ( .A(n_83), .Y(n_1178) );
INVx1_ASAP7_75t_L g1383 ( .A(n_84), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_85), .A2(n_160), .B1(n_526), .B2(n_527), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_85), .A2(n_160), .B1(n_600), .B2(n_602), .Y(n_599) );
INVx1_ASAP7_75t_L g976 ( .A(n_86), .Y(n_976) );
INVx1_ASAP7_75t_L g1071 ( .A(n_87), .Y(n_1071) );
OAI222xp33_ASAP7_75t_L g875 ( .A1(n_88), .A2(n_181), .B1(n_224), .B2(n_620), .C1(n_876), .C2(n_879), .Y(n_875) );
INVx1_ASAP7_75t_L g896 ( .A(n_88), .Y(n_896) );
AO22x2_ASAP7_75t_L g870 ( .A1(n_89), .A2(n_871), .B1(n_872), .B2(n_926), .Y(n_870) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_89), .Y(n_871) );
AO221x1_ASAP7_75t_L g1326 ( .A1(n_89), .A2(n_165), .B1(n_1285), .B2(n_1293), .C(n_1327), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_90), .A2(n_106), .B1(n_565), .B2(n_566), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_90), .A2(n_106), .B1(n_630), .B2(n_632), .Y(n_917) );
INVx1_ASAP7_75t_L g358 ( .A(n_91), .Y(n_358) );
INVx1_ASAP7_75t_L g476 ( .A(n_91), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_92), .A2(n_155), .B1(n_632), .B2(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g671 ( .A(n_92), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_93), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_94), .A2(n_215), .B1(n_955), .B2(n_960), .C(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1219 ( .A(n_95), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_95), .A2(n_274), .B1(n_1266), .B2(n_1268), .Y(n_1265) );
INVx1_ASAP7_75t_L g1329 ( .A(n_96), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_97), .Y(n_1528) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_98), .A2(n_136), .B1(n_513), .B2(n_526), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_98), .A2(n_136), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22x1_ASAP7_75t_L g928 ( .A1(n_99), .A2(n_929), .B1(n_930), .B2(n_977), .Y(n_928) );
INVxp67_ASAP7_75t_SL g977 ( .A(n_99), .Y(n_977) );
INVx1_ASAP7_75t_L g999 ( .A(n_100), .Y(n_999) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_100), .A2(n_578), .B1(n_597), .B2(n_1017), .C(n_1020), .Y(n_1016) );
INVx1_ASAP7_75t_L g882 ( .A(n_102), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_102), .A2(n_224), .B1(n_566), .B2(n_654), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_104), .A2(n_225), .B1(n_1285), .B2(n_1293), .Y(n_1342) );
INVx1_ASAP7_75t_L g1543 ( .A(n_105), .Y(n_1543) );
INVx1_ASAP7_75t_L g616 ( .A(n_107), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_107), .A2(n_193), .B1(n_374), .B2(n_647), .Y(n_646) );
INVxp33_ASAP7_75t_SL g1135 ( .A(n_108), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_109), .Y(n_749) );
INVx1_ASAP7_75t_L g819 ( .A(n_110), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_111), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_112), .A2(n_182), .B1(n_632), .B2(n_938), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_112), .A2(n_549), .B1(n_959), .B2(n_961), .C(n_964), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_113), .A2(n_220), .B1(n_527), .B2(n_660), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_113), .A2(n_220), .B1(n_386), .B2(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_114), .A2(n_245), .B1(n_379), .B2(n_384), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_114), .A2(n_245), .B1(n_414), .B2(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g753 ( .A(n_115), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_115), .A2(n_578), .B1(n_774), .B2(n_780), .C(n_783), .Y(n_773) );
INVx1_ASAP7_75t_L g286 ( .A(n_117), .Y(n_286) );
INVxp67_ASAP7_75t_SL g1179 ( .A(n_118), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_120), .Y(n_623) );
INVx1_ASAP7_75t_L g1334 ( .A(n_121), .Y(n_1334) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_122), .Y(n_320) );
INVx1_ASAP7_75t_L g1002 ( .A(n_124), .Y(n_1002) );
OAI211xp5_ASAP7_75t_SL g1024 ( .A1(n_124), .A2(n_549), .B(n_1025), .C(n_1031), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_125), .A2(n_207), .B1(n_1310), .B2(n_1313), .Y(n_1318) );
INVx1_ASAP7_75t_L g1333 ( .A(n_127), .Y(n_1333) );
INVx1_ASAP7_75t_L g885 ( .A(n_128), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g1240 ( .A(n_129), .Y(n_1240) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_130), .B(n_465), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g1228 ( .A(n_131), .Y(n_1228) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_132), .A2(n_183), .B1(n_1285), .B2(n_1293), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_133), .A2(n_253), .B1(n_410), .B2(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g455 ( .A(n_133), .Y(n_455) );
INVx1_ASAP7_75t_L g1202 ( .A(n_134), .Y(n_1202) );
INVx1_ASAP7_75t_L g890 ( .A(n_135), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g1231 ( .A(n_137), .Y(n_1231) );
AOI22xp5_ASAP7_75t_L g1343 ( .A1(n_138), .A2(n_279), .B1(n_1310), .B2(n_1313), .Y(n_1343) );
XOR2xp5_ASAP7_75t_L g1086 ( .A(n_139), .B(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1109 ( .A(n_140), .Y(n_1109) );
INVx1_ASAP7_75t_L g1381 ( .A(n_141), .Y(n_1381) );
INVx1_ASAP7_75t_L g829 ( .A(n_142), .Y(n_829) );
INVx1_ASAP7_75t_L g1094 ( .A(n_143), .Y(n_1094) );
INVx1_ASAP7_75t_L g1093 ( .A(n_144), .Y(n_1093) );
INVx1_ASAP7_75t_L g1091 ( .A(n_145), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_146), .A2(n_237), .B1(n_527), .B2(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g668 ( .A(n_146), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_147), .Y(n_993) );
INVx1_ASAP7_75t_L g700 ( .A(n_148), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_148), .A2(n_151), .B1(n_422), .B2(n_723), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_149), .A2(n_226), .B1(n_764), .B2(n_766), .Y(n_1008) );
INVx1_ASAP7_75t_L g1033 ( .A(n_149), .Y(n_1033) );
INVx1_ASAP7_75t_L g1004 ( .A(n_150), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_150), .A2(n_261), .B1(n_771), .B2(n_772), .Y(n_1015) );
INVx1_ASAP7_75t_L g701 ( .A(n_151), .Y(n_701) );
INVx1_ASAP7_75t_L g595 ( .A(n_152), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_153), .A2(n_219), .B1(n_518), .B2(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g585 ( .A(n_153), .Y(n_585) );
INVx1_ASAP7_75t_L g663 ( .A(n_155), .Y(n_663) );
INVx1_ASAP7_75t_L g1105 ( .A(n_156), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_156), .A2(n_190), .B1(n_408), .B2(n_936), .Y(n_1119) );
INVx1_ASAP7_75t_L g1555 ( .A(n_157), .Y(n_1555) );
AOI22x1_ASAP7_75t_SL g673 ( .A1(n_159), .A2(n_674), .B1(n_724), .B2(n_725), .Y(n_673) );
INVx1_ASAP7_75t_L g724 ( .A(n_159), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_161), .Y(n_1040) );
INVxp33_ASAP7_75t_SL g1137 ( .A(n_162), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1157 ( .A1(n_162), .A2(n_205), .B1(n_1152), .B2(n_1158), .Y(n_1157) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_163), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_164), .Y(n_1197) );
INVx1_ASAP7_75t_L g678 ( .A(n_166), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_166), .A2(n_230), .B1(n_368), .B2(n_706), .Y(n_710) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_167), .Y(n_288) );
AND3x2_ASAP7_75t_L g1289 ( .A(n_167), .B(n_286), .C(n_1290), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_167), .B(n_286), .Y(n_1297) );
XNOR2xp5_ASAP7_75t_L g728 ( .A(n_169), .B(n_729), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_170), .Y(n_768) );
INVx1_ASAP7_75t_L g1591 ( .A(n_171), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g1599 ( .A1(n_171), .A2(n_578), .B1(n_783), .B2(n_1600), .C(n_1605), .Y(n_1599) );
INVx1_ASAP7_75t_L g823 ( .A(n_172), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_172), .A2(n_549), .B1(n_844), .B2(n_852), .C(n_858), .Y(n_843) );
INVx2_ASAP7_75t_L g299 ( .A(n_173), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_175), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g1587 ( .A(n_176), .Y(n_1587) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_177), .A2(n_178), .B1(n_764), .B2(n_766), .Y(n_827) );
INVx1_ASAP7_75t_L g859 ( .A(n_177), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_178), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_179), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_180), .A2(n_215), .B1(n_472), .B2(n_479), .Y(n_1010) );
INVx1_ASAP7_75t_L g1028 ( .A(n_180), .Y(n_1028) );
INVx1_ASAP7_75t_L g898 ( .A(n_181), .Y(n_898) );
INVx1_ASAP7_75t_L g957 ( .A(n_182), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_184), .A2(n_228), .B1(n_408), .B2(n_1006), .Y(n_1526) );
INVx1_ASAP7_75t_L g1550 ( .A(n_184), .Y(n_1550) );
INVx1_ASAP7_75t_L g1544 ( .A(n_185), .Y(n_1544) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_186), .A2(n_210), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_186), .A2(n_210), .B1(n_1163), .B2(n_1164), .Y(n_1162) );
INVx1_ASAP7_75t_L g1077 ( .A(n_187), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_188), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g807 ( .A(n_189), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g1106 ( .A(n_190), .Y(n_1106) );
INVx1_ASAP7_75t_L g1290 ( .A(n_191), .Y(n_1290) );
INVx1_ASAP7_75t_L g535 ( .A(n_192), .Y(n_535) );
INVx1_ASAP7_75t_L g622 ( .A(n_193), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g1596 ( .A1(n_194), .A2(n_199), .B1(n_764), .B2(n_766), .Y(n_1596) );
INVx1_ASAP7_75t_L g1615 ( .A(n_194), .Y(n_1615) );
INVx1_ASAP7_75t_L g625 ( .A(n_195), .Y(n_625) );
INVx1_ASAP7_75t_L g1049 ( .A(n_197), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_197), .A2(n_578), .B1(n_783), .B2(n_1064), .C(n_1066), .Y(n_1063) );
INVx1_ASAP7_75t_L g1051 ( .A(n_198), .Y(n_1051) );
OAI211xp5_ASAP7_75t_L g1068 ( .A1(n_198), .A2(n_549), .B(n_1069), .C(n_1075), .Y(n_1068) );
INVx1_ASAP7_75t_L g1614 ( .A(n_199), .Y(n_1614) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_200), .A2(n_246), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_200), .A2(n_246), .B1(n_419), .B2(n_718), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g1516 ( .A1(n_201), .A2(n_203), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
OAI221xp5_ASAP7_75t_L g1546 ( .A1(n_201), .A2(n_203), .B1(n_1210), .B2(n_1213), .C(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1222 ( .A(n_202), .Y(n_1222) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_202), .A2(n_271), .B1(n_414), .B2(n_1262), .C(n_1264), .Y(n_1261) );
INVx1_ASAP7_75t_L g1582 ( .A(n_204), .Y(n_1582) );
INVxp33_ASAP7_75t_L g1140 ( .A(n_205), .Y(n_1140) );
INVx1_ASAP7_75t_L g301 ( .A(n_206), .Y(n_301) );
INVx2_ASAP7_75t_L g400 ( .A(n_206), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g1322 ( .A1(n_208), .A2(n_227), .B1(n_1310), .B2(n_1313), .Y(n_1322) );
INVx1_ASAP7_75t_L g903 ( .A(n_209), .Y(n_903) );
INVx1_ASAP7_75t_L g822 ( .A(n_211), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_211), .A2(n_578), .B1(n_783), .B2(n_833), .C(n_839), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g1107 ( .A1(n_212), .A2(n_549), .B1(n_1108), .B2(n_1110), .C(n_1115), .Y(n_1107) );
INVx1_ASAP7_75t_L g1101 ( .A(n_213), .Y(n_1101) );
INVx1_ASAP7_75t_L g1328 ( .A(n_214), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_216), .Y(n_743) );
XNOR2x1_ASAP7_75t_L g1188 ( .A(n_217), .B(n_1189), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_218), .A2(n_275), .B1(n_757), .B2(n_1006), .Y(n_1588) );
INVx1_ASAP7_75t_L g1601 ( .A(n_218), .Y(n_1601) );
INVx1_ASAP7_75t_L g589 ( .A(n_219), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g1044 ( .A(n_221), .Y(n_1044) );
INVx1_ASAP7_75t_L g989 ( .A(n_222), .Y(n_989) );
INVx1_ASAP7_75t_L g348 ( .A(n_223), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_223), .A2(n_233), .B1(n_368), .B2(n_372), .Y(n_393) );
INVx1_ASAP7_75t_L g1032 ( .A(n_226), .Y(n_1032) );
INVx1_ASAP7_75t_L g1559 ( .A(n_228), .Y(n_1559) );
INVx1_ASAP7_75t_L g1534 ( .A(n_229), .Y(n_1534) );
INVx1_ASAP7_75t_L g335 ( .A(n_233), .Y(n_335) );
INVx1_ASAP7_75t_L g1586 ( .A(n_235), .Y(n_1586) );
AOI21xp33_ASAP7_75t_L g1606 ( .A1(n_235), .A2(n_956), .B(n_1030), .Y(n_1606) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_236), .Y(n_815) );
INVx1_ASAP7_75t_L g669 ( .A(n_237), .Y(n_669) );
INVx1_ASAP7_75t_L g991 ( .A(n_238), .Y(n_991) );
INVx1_ASAP7_75t_L g1288 ( .A(n_239), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_239), .B(n_1299), .Y(n_1304) );
INVx1_ASAP7_75t_L g452 ( .A(n_240), .Y(n_452) );
INVx1_ASAP7_75t_L g1143 ( .A(n_241), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_241), .A2(n_262), .B1(n_441), .B2(n_665), .Y(n_1176) );
INVx1_ASAP7_75t_L g1097 ( .A(n_242), .Y(n_1097) );
INVx1_ASAP7_75t_L g1139 ( .A(n_243), .Y(n_1139) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_244), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_247), .A2(n_249), .B1(n_764), .B2(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g796 ( .A(n_247), .Y(n_796) );
INVx1_ASAP7_75t_L g1593 ( .A(n_248), .Y(n_1593) );
OAI211xp5_ASAP7_75t_SL g1607 ( .A1(n_248), .A2(n_549), .B(n_1608), .C(n_1613), .Y(n_1607) );
INVx1_ASAP7_75t_L g797 ( .A(n_249), .Y(n_797) );
INVx1_ASAP7_75t_L g327 ( .A(n_250), .Y(n_327) );
AO22x1_ASAP7_75t_L g1307 ( .A1(n_251), .A2(n_264), .B1(n_1293), .B2(n_1308), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g1533 ( .A(n_252), .Y(n_1533) );
INVx1_ASAP7_75t_L g430 ( .A(n_253), .Y(n_430) );
INVx2_ASAP7_75t_L g298 ( .A(n_254), .Y(n_298) );
AO22x1_ASAP7_75t_L g1309 ( .A1(n_255), .A2(n_269), .B1(n_1310), .B2(n_1313), .Y(n_1309) );
INVx1_ASAP7_75t_L g1567 ( .A(n_255), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_255), .A2(n_1573), .B1(n_1577), .B2(n_1619), .Y(n_1572) );
INVx1_ASAP7_75t_L g847 ( .A(n_256), .Y(n_847) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_256), .A2(n_267), .B1(n_472), .B2(n_479), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g1204 ( .A1(n_257), .A2(n_263), .B1(n_1205), .B2(n_1210), .C(n_1213), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_257), .A2(n_263), .B1(n_1246), .B2(n_1249), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_258), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_259), .A2(n_260), .B1(n_519), .B2(n_523), .Y(n_522) );
OAI211xp5_ASAP7_75t_SL g548 ( .A1(n_259), .A2(n_549), .B(n_554), .C(n_571), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g577 ( .A1(n_260), .A2(n_578), .B1(n_580), .B2(n_592), .C(n_597), .Y(n_577) );
INVx1_ASAP7_75t_L g1007 ( .A(n_261), .Y(n_1007) );
INVx1_ASAP7_75t_L g1144 ( .A(n_262), .Y(n_1144) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_265), .Y(n_1532) );
INVx1_ASAP7_75t_L g813 ( .A(n_266), .Y(n_813) );
INVx1_ASAP7_75t_L g854 ( .A(n_267), .Y(n_854) );
INVx1_ASAP7_75t_L g1224 ( .A(n_271), .Y(n_1224) );
BUFx3_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
INVx1_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
BUFx3_ASAP7_75t_L g318 ( .A(n_273), .Y(n_318) );
INVx1_ASAP7_75t_L g355 ( .A(n_273), .Y(n_355) );
INVx1_ASAP7_75t_L g1226 ( .A(n_274), .Y(n_1226) );
INVx1_ASAP7_75t_L g1604 ( .A(n_275), .Y(n_1604) );
INVx1_ASAP7_75t_L g1611 ( .A(n_276), .Y(n_1611) );
INVx1_ASAP7_75t_L g950 ( .A(n_277), .Y(n_950) );
INVx1_ASAP7_75t_L g1013 ( .A(n_280), .Y(n_1013) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_302), .B(n_1278), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
AND2x4_ASAP7_75t_L g1571 ( .A(n_284), .B(n_290), .Y(n_1571) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g1576 ( .A(n_285), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_285), .B(n_287), .Y(n_1620) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_287), .B(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g458 ( .A(n_292), .B(n_425), .Y(n_458) );
OR2x6_ASAP7_75t_L g672 ( .A(n_292), .B(n_425), .Y(n_672) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g366 ( .A(n_293), .B(n_301), .Y(n_366) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g956 ( .A(n_294), .B(n_447), .Y(n_956) );
INVx8_ASAP7_75t_L g454 ( .A(n_295), .Y(n_454) );
OR2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
OR2x6_ASAP7_75t_L g457 ( .A(n_296), .B(n_446), .Y(n_457) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_296), .Y(n_588) );
INVx2_ASAP7_75t_SL g842 ( .A(n_296), .Y(n_842) );
INVx1_ASAP7_75t_L g849 ( .A(n_296), .Y(n_849) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_296), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_296), .B(n_1209), .Y(n_1238) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g371 ( .A(n_298), .B(n_299), .Y(n_371) );
INVx1_ASAP7_75t_L g376 ( .A(n_298), .Y(n_376) );
INVx2_ASAP7_75t_L g381 ( .A(n_298), .Y(n_381) );
AND2x4_ASAP7_75t_L g387 ( .A(n_298), .B(n_377), .Y(n_387) );
INVx1_ASAP7_75t_L g443 ( .A(n_298), .Y(n_443) );
INVx2_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
INVx1_ASAP7_75t_L g383 ( .A(n_299), .Y(n_383) );
INVx1_ASAP7_75t_L g440 ( .A(n_299), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_299), .B(n_381), .Y(n_558) );
INVx1_ASAP7_75t_L g584 ( .A(n_299), .Y(n_584) );
AND2x4_ASAP7_75t_L g439 ( .A(n_300), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g441 ( .A(n_301), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g666 ( .A(n_301), .B(n_442), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_978), .B2(n_979), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
XNOR2x1_ASAP7_75t_L g304 ( .A(n_305), .B(n_609), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_461), .B1(n_607), .B2(n_608), .Y(n_305) );
INVx2_ASAP7_75t_L g607 ( .A(n_306), .Y(n_607) );
INVx1_ASAP7_75t_L g460 ( .A(n_307), .Y(n_460) );
AOI211x1_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_356), .B(n_361), .C(n_428), .Y(n_307) );
NAND4xp25_ASAP7_75t_L g308 ( .A(n_309), .B(n_319), .C(n_334), .D(n_347), .Y(n_308) );
NAND4xp25_ASAP7_75t_L g1133 ( .A(n_309), .B(n_1134), .C(n_1138), .D(n_1141), .Y(n_1133) );
INVx5_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_310), .A2(n_616), .B(n_617), .C(n_618), .Y(n_615) );
CKINVDCx8_ASAP7_75t_R g683 ( .A(n_310), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_310), .B(n_875), .Y(n_874) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_315), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x6_ASAP7_75t_L g353 ( .A(n_312), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g689 ( .A(n_312), .Y(n_689) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x6_ASAP7_75t_L g345 ( .A(n_313), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_314), .Y(n_323) );
INVx1_ASAP7_75t_L g330 ( .A(n_314), .Y(n_330) );
AND2x2_ASAP7_75t_L g406 ( .A(n_314), .B(n_358), .Y(n_406) );
INVx2_ASAP7_75t_L g427 ( .A(n_314), .Y(n_427) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_315), .Y(n_337) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_315), .Y(n_412) );
INVx2_ASAP7_75t_L g633 ( .A(n_315), .Y(n_633) );
INVx1_ASAP7_75t_L g734 ( .A(n_315), .Y(n_734) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_316), .Y(n_521) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g325 ( .A(n_317), .Y(n_325) );
AND2x4_ASAP7_75t_L g354 ( .A(n_317), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g326 ( .A(n_318), .Y(n_326) );
AND2x4_ASAP7_75t_L g332 ( .A(n_318), .B(n_333), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B1(n_327), .B2(n_328), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_320), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_321), .A2(n_349), .B1(n_622), .B2(n_623), .Y(n_621) );
INVx4_ASAP7_75t_L g691 ( .A(n_321), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_321), .A2(n_349), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_321), .A2(n_328), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
AND2x4_ASAP7_75t_L g340 ( .A(n_322), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx6_ASAP7_75t_L g351 ( .A(n_324), .Y(n_351) );
INVx2_ASAP7_75t_L g420 ( .A(n_324), .Y(n_420) );
BUFx2_ASAP7_75t_L g518 ( .A(n_324), .Y(n_518) );
AND2x2_ASAP7_75t_L g538 ( .A(n_324), .B(n_502), .Y(n_538) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g346 ( .A(n_325), .Y(n_346) );
INVx1_ASAP7_75t_L g343 ( .A(n_326), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_328), .A2(n_353), .B1(n_625), .B2(n_626), .Y(n_624) );
INVx4_ASAP7_75t_L g686 ( .A(n_328), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_328), .A2(n_353), .B1(n_885), .B2(n_886), .Y(n_884) );
AND2x6_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
AND2x4_ASAP7_75t_L g349 ( .A(n_329), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g1136 ( .A(n_329), .B(n_350), .Y(n_1136) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g877 ( .A(n_330), .B(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_331), .Y(n_942) );
BUFx6f_ASAP7_75t_L g1006 ( .A(n_331), .Y(n_1006) );
INVx2_ASAP7_75t_L g1128 ( .A(n_331), .Y(n_1128) );
INVx1_ASAP7_75t_L g1165 ( .A(n_331), .Y(n_1165) );
BUFx6f_ASAP7_75t_L g1595 ( .A(n_331), .Y(n_1595) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_332), .Y(n_417) );
INVx1_ASAP7_75t_L g473 ( .A(n_332), .Y(n_473) );
INVx2_ASAP7_75t_L g516 ( .A(n_332), .Y(n_516) );
INVx1_ASAP7_75t_L g716 ( .A(n_332), .Y(n_716) );
INVx1_ASAP7_75t_L g482 ( .A(n_333), .Y(n_482) );
AOI222xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_338), .B2(n_339), .C1(n_344), .C2(n_345), .Y(n_334) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_337), .Y(n_617) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_337), .Y(n_1168) );
BUFx4f_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g619 ( .A(n_340), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_340), .A2(n_345), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI222xp33_ASAP7_75t_L g1141 ( .A1(n_340), .A2(n_345), .B1(n_718), .B2(n_1142), .C1(n_1143), .C2(n_1144), .Y(n_1141) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g878 ( .A(n_342), .Y(n_878) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g499 ( .A(n_343), .Y(n_499) );
INVx3_ASAP7_75t_L g620 ( .A(n_345), .Y(n_620) );
BUFx3_ASAP7_75t_L g508 ( .A(n_346), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_352), .B2(n_353), .Y(n_347) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_351), .Y(n_524) );
INVx2_ASAP7_75t_L g631 ( .A(n_351), .Y(n_631) );
INVx1_ASAP7_75t_L g921 ( .A(n_351), .Y(n_921) );
INVx2_ASAP7_75t_SL g940 ( .A(n_351), .Y(n_940) );
CKINVDCx6p67_ASAP7_75t_R g685 ( .A(n_353), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_353), .A2(n_1135), .B1(n_1136), .B2(n_1137), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_354), .Y(n_415) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_354), .Y(n_423) );
INVx2_ASAP7_75t_SL g492 ( .A(n_354), .Y(n_492) );
BUFx2_ASAP7_75t_L g512 ( .A(n_354), .Y(n_512) );
BUFx3_ASAP7_75t_L g739 ( .A(n_354), .Y(n_739) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_354), .Y(n_757) );
BUFx2_ASAP7_75t_L g923 ( .A(n_354), .Y(n_923) );
BUFx6f_ASAP7_75t_L g1054 ( .A(n_354), .Y(n_1054) );
INVx1_ASAP7_75t_L g483 ( .A(n_355), .Y(n_483) );
AO211x2_ASAP7_75t_L g613 ( .A1(n_356), .A2(n_614), .B(n_627), .C(n_661), .Y(n_613) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_356), .Y(n_887) );
INVx1_ASAP7_75t_L g1146 ( .A(n_356), .Y(n_1146) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AND2x4_ASAP7_75t_L g692 ( .A(n_357), .B(n_359), .Y(n_692) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g426 ( .A(n_358), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g972 ( .A(n_359), .Y(n_972) );
BUFx2_ASAP7_75t_L g1277 ( .A(n_359), .Y(n_1277) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g365 ( .A(n_360), .Y(n_365) );
OR2x6_ASAP7_75t_L g1216 ( .A(n_360), .B(n_956), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_402), .Y(n_361) );
AOI33xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .A3(n_378), .B1(n_388), .B2(n_393), .B3(n_394), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_364), .B(n_650), .C(n_653), .Y(n_649) );
INVx2_ASAP7_75t_L g1150 ( .A(n_364), .Y(n_1150) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
OR2x6_ASAP7_75t_L g404 ( .A(n_365), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g540 ( .A(n_365), .Y(n_540) );
BUFx2_ASAP7_75t_L g606 ( .A(n_365), .Y(n_606) );
OR2x2_ASAP7_75t_L g636 ( .A(n_365), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g703 ( .A(n_365), .B(n_366), .Y(n_703) );
OR2x2_ASAP7_75t_L g736 ( .A(n_365), .B(n_405), .Y(n_736) );
INVx1_ASAP7_75t_L g591 ( .A(n_366), .Y(n_591) );
BUFx2_ASAP7_75t_SL g1067 ( .A(n_366), .Y(n_1067) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g546 ( .A(n_370), .Y(n_546) );
INVx2_ASAP7_75t_SL g1030 ( .A(n_370), .Y(n_1030) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_371), .Y(n_568) );
AOI211xp5_ASAP7_75t_L g662 ( .A1(n_372), .A2(n_434), .B(n_663), .C(n_664), .Y(n_662) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g895 ( .A(n_373), .Y(n_895) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx3_ASAP7_75t_L g433 ( .A(n_375), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_375), .B(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_375), .Y(n_655) );
BUFx3_ASAP7_75t_L g955 ( .A(n_375), .Y(n_955) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_380), .Y(n_391) );
AND2x4_ASAP7_75t_L g445 ( .A(n_380), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g601 ( .A(n_380), .B(n_553), .Y(n_601) );
INVx1_ASAP7_75t_L g641 ( .A(n_380), .Y(n_641) );
BUFx2_ASAP7_75t_L g651 ( .A(n_380), .Y(n_651) );
BUFx6f_ASAP7_75t_L g953 ( .A(n_380), .Y(n_953) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g576 ( .A(n_381), .Y(n_576) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_385), .A2(n_1026), .B1(n_1027), .B2(n_1028), .C(n_1029), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_385), .A2(n_1040), .B1(n_1042), .B2(n_1065), .Y(n_1064) );
OAI221xp5_ASAP7_75t_L g1608 ( .A1(n_385), .A2(n_1609), .B1(n_1610), .B2(n_1611), .C(n_1612), .Y(n_1608) );
INVx4_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g392 ( .A(n_386), .Y(n_392) );
INVx2_ASAP7_75t_SL g1072 ( .A(n_386), .Y(n_1072) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_386), .Y(n_1102) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_386), .Y(n_1159) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g451 ( .A(n_387), .Y(n_451) );
INVx1_ASAP7_75t_L g563 ( .A(n_387), .Y(n_563) );
INVx3_ASAP7_75t_L g645 ( .A(n_387), .Y(n_645) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_391), .B(n_1196), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_391), .B(n_1196), .Y(n_1545) );
INVx1_ASAP7_75t_L g1560 ( .A(n_392), .Y(n_1560) );
AOI33xp33_ASAP7_75t_L g702 ( .A1(n_394), .A2(n_703), .A3(n_704), .B1(n_708), .B2(n_709), .B3(n_710), .Y(n_702) );
INVx2_ASAP7_75t_L g1234 ( .A(n_394), .Y(n_1234) );
INVx6_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx5_ASAP7_75t_L g648 ( .A(n_395), .Y(n_648) );
OR2x6_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_396), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g474 ( .A(n_397), .B(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_397), .B(n_553), .Y(n_1196) );
INVx2_ASAP7_75t_L g570 ( .A(n_398), .Y(n_570) );
BUFx2_ASAP7_75t_L g960 ( .A(n_398), .Y(n_960) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
AOI33xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_407), .A3(n_413), .B1(n_418), .B2(n_421), .B3(n_424), .Y(n_402) );
AOI33xp33_ASAP7_75t_L g711 ( .A1(n_403), .A2(n_424), .A3(n_712), .B1(n_717), .B2(n_719), .B3(n_722), .Y(n_711) );
AOI33xp33_ASAP7_75t_L g1161 ( .A1(n_403), .A2(n_424), .A3(n_1162), .B1(n_1166), .B2(n_1169), .B3(n_1172), .Y(n_1161) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g510 ( .A(n_404), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g1118 ( .A(n_404), .Y(n_1118) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g637 ( .A(n_406), .Y(n_637) );
INVx2_ASAP7_75t_SL g1264 ( .A(n_406), .Y(n_1264) );
BUFx3_ASAP7_75t_L g1525 ( .A(n_406), .Y(n_1525) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_409), .Y(n_720) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_412), .Y(n_721) );
AND2x4_ASAP7_75t_L g1269 ( .A(n_412), .B(n_1270), .Y(n_1269) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g714 ( .A(n_415), .Y(n_714) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_415), .B(n_1244), .Y(n_1243) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g814 ( .A(n_417), .Y(n_814) );
INVx1_ASAP7_75t_L g990 ( .A(n_417), .Y(n_990) );
INVx1_ASAP7_75t_L g1041 ( .A(n_417), .Y(n_1041) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g487 ( .A(n_420), .Y(n_487) );
BUFx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx4f_ASAP7_75t_L g526 ( .A(n_423), .Y(n_526) );
INVx1_ASAP7_75t_L g806 ( .A(n_423), .Y(n_806) );
INVx4_ASAP7_75t_L g762 ( .A(n_424), .Y(n_762) );
BUFx4f_ASAP7_75t_L g1129 ( .A(n_424), .Y(n_1129) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AND2x4_ASAP7_75t_L g528 ( .A(n_425), .B(n_426), .Y(n_528) );
AND2x4_ASAP7_75t_L g537 ( .A(n_425), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g1256 ( .A(n_426), .Y(n_1256) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_426), .Y(n_1512) );
AND2x4_ASAP7_75t_L g502 ( .A(n_427), .B(n_503), .Y(n_502) );
AOI31xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_444), .A3(n_453), .B(n_458), .Y(n_428) );
AOI211xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_434), .C(n_437), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g1174 ( .A1(n_431), .A2(n_434), .B(n_1175), .C(n_1176), .Y(n_1174) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g565 ( .A(n_432), .Y(n_565) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g550 ( .A(n_433), .B(n_551), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_434), .B(n_695), .C(n_698), .Y(n_694) );
CKINVDCx11_ASAP7_75t_R g904 ( .A(n_434), .Y(n_904) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g901 ( .A(n_436), .Y(n_901) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g665 ( .A(n_439), .Y(n_665) );
INVx2_ASAP7_75t_L g696 ( .A(n_439), .Y(n_696) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_440), .Y(n_573) );
INVx1_ASAP7_75t_L g969 ( .A(n_440), .Y(n_969) );
INVx1_ASAP7_75t_L g900 ( .A(n_442), .Y(n_900) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g583 ( .A(n_443), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_443), .B(n_584), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_448), .B1(n_449), .B2(n_452), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_445), .A2(n_449), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_445), .A2(n_449), .B1(n_700), .B2(n_701), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_445), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g1177 ( .A1(n_445), .A2(n_892), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AND2x4_ASAP7_75t_L g449 ( .A(n_446), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g892 ( .A(n_446), .B(n_450), .Y(n_892) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_451), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_454), .A2(n_456), .B1(n_623), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_454), .A2(n_456), .B1(n_883), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g1180 ( .A1(n_454), .A2(n_456), .B1(n_1139), .B2(n_1181), .Y(n_1180) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI31xp33_ASAP7_75t_L g1173 ( .A1(n_458), .A2(n_1174), .A3(n_1177), .B(n_1180), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g608 ( .A(n_464), .Y(n_608) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_534), .C(n_547), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_493), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_484), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_477), .B2(n_478), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_470), .A2(n_489), .B1(n_555), .B2(n_559), .C(n_564), .Y(n_554) );
AOI222xp33_ASAP7_75t_L g973 ( .A1(n_471), .A2(n_486), .B1(n_537), .B2(n_962), .C1(n_965), .C2(n_974), .Y(n_973) );
CKINVDCx6p67_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_473), .A2(n_738), .B1(n_825), .B2(n_826), .Y(n_824) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_473), .B(n_474), .Y(n_1080) );
INVx2_ASAP7_75t_L g1268 ( .A(n_473), .Y(n_1268) );
OR2x6_ASAP7_75t_L g479 ( .A(n_474), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g488 ( .A(n_474), .Y(n_488) );
OR2x2_ASAP7_75t_L g802 ( .A(n_474), .B(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g805 ( .A(n_474), .B(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g1244 ( .A(n_475), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_475), .B(n_690), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_475), .B(n_516), .Y(n_1275) );
INVx1_ASAP7_75t_L g503 ( .A(n_476), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_478), .A2(n_490), .B1(n_963), .B2(n_976), .Y(n_975) );
CKINVDCx6p67_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_480), .A2(n_751), .B1(n_753), .B2(n_754), .Y(n_750) );
BUFx3_ASAP7_75t_L g818 ( .A(n_480), .Y(n_818) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g748 ( .A(n_481), .Y(n_748) );
INVx1_ASAP7_75t_L g996 ( .A(n_481), .Y(n_996) );
BUFx4f_ASAP7_75t_L g1001 ( .A(n_481), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_481), .Y(n_1046) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OR2x2_ASAP7_75t_L g690 ( .A(n_482), .B(n_483), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_489), .B2(n_490), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_486), .A2(n_490), .B1(n_1093), .B2(n_1094), .C(n_1095), .Y(n_1092) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
BUFx2_ASAP7_75t_L g1167 ( .A(n_487), .Y(n_1167) );
AND2x2_ASAP7_75t_L g490 ( .A(n_488), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g660 ( .A(n_492), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_509), .C(n_529), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_504), .B2(n_505), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_495), .A2(n_504), .B1(n_572), .B2(n_574), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g1089 ( .A1(n_496), .A2(n_505), .B1(n_732), .B2(n_1090), .C(n_1091), .Y(n_1089) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g765 ( .A(n_497), .Y(n_765) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g1248 ( .A(n_499), .Y(n_1248) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x6_ASAP7_75t_L g506 ( .A(n_501), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g533 ( .A(n_501), .Y(n_533) );
OR2x2_ASAP7_75t_L g766 ( .A(n_501), .B(n_507), .Y(n_766) );
AND2x4_ASAP7_75t_L g1247 ( .A(n_502), .B(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1250 ( .A(n_502), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_502), .B(n_508), .Y(n_1519) );
BUFx2_ASAP7_75t_L g1530 ( .A(n_502), .Y(n_1530) );
AOI221xp5_ASAP7_75t_L g943 ( .A1(n_505), .A2(n_732), .B1(n_765), .B2(n_944), .C(n_945), .Y(n_943) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_507), .B(n_1250), .Y(n_1249) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI33xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .A3(n_517), .B1(n_522), .B2(n_525), .B3(n_528), .Y(n_509) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g527 ( .A(n_514), .Y(n_527) );
INVx2_ASAP7_75t_SL g742 ( .A(n_514), .Y(n_742) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g679 ( .A(n_520), .Y(n_679) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_521), .Y(n_532) );
BUFx3_ASAP7_75t_L g718 ( .A(n_521), .Y(n_718) );
BUFx4f_ASAP7_75t_L g936 ( .A(n_521), .Y(n_936) );
AND2x4_ASAP7_75t_L g1260 ( .A(n_521), .B(n_1244), .Y(n_1260) );
INVx1_ASAP7_75t_L g1263 ( .A(n_521), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1529 ( .A(n_521), .B(n_1530), .Y(n_1529) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g658 ( .A(n_524), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_528), .B(n_657), .C(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g925 ( .A(n_528), .Y(n_925) );
AOI33xp33_ASAP7_75t_L g932 ( .A1(n_528), .A2(n_933), .A3(n_934), .B1(n_935), .B2(n_937), .B3(n_941), .Y(n_932) );
INVx1_ASAP7_75t_L g1057 ( .A(n_528), .Y(n_1057) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g1171 ( .A(n_532), .Y(n_1171) );
AND2x2_ASAP7_75t_L g732 ( .A(n_533), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_536), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_536), .B(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_536), .B(n_1013), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_536), .B(n_1060), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_536), .B(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_536), .B(n_1582), .Y(n_1581) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g1239 ( .A(n_537), .Y(n_1239) );
NOR2xp67_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g798 ( .A(n_540), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
AND2x2_ASAP7_75t_L g572 ( .A(n_542), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g860 ( .A(n_542), .B(n_573), .Y(n_860) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x6_ASAP7_75t_L g575 ( .A(n_543), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g597 ( .A(n_543), .B(n_598), .Y(n_597) );
OR2x6_ASAP7_75t_L g783 ( .A(n_543), .B(n_598), .Y(n_783) );
INVx1_ASAP7_75t_L g970 ( .A(n_543), .Y(n_970) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g647 ( .A(n_546), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_577), .A3(n_599), .B(n_604), .Y(n_547) );
INVx8_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g603 ( .A(n_551), .B(n_562), .Y(n_603) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g579 ( .A(n_553), .B(n_568), .Y(n_579) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_556), .Y(n_1111) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g594 ( .A(n_557), .Y(n_594) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_557), .Y(n_776) );
INVx1_ASAP7_75t_L g1070 ( .A(n_557), .Y(n_1070) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g788 ( .A(n_558), .Y(n_788) );
INVx1_ASAP7_75t_L g836 ( .A(n_558), .Y(n_836) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g652 ( .A(n_561), .Y(n_652) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g964 ( .A1(n_566), .A2(n_965), .B(n_966), .C(n_970), .Y(n_964) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_568), .Y(n_705) );
INVx1_ASAP7_75t_L g851 ( .A(n_569), .Y(n_851) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_572), .A2(n_574), .B1(n_796), .B2(n_797), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g1115 ( .A1(n_572), .A2(n_574), .B1(n_1090), .B2(n_1091), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_572), .A2(n_574), .B1(n_1614), .B2(n_1615), .Y(n_1613) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_574), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_574), .A2(n_860), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_574), .A2(n_860), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
CKINVDCx11_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g1212 ( .A(n_576), .Y(n_1212) );
CKINVDCx6p67_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g951 ( .A1(n_579), .A2(n_952), .B1(n_954), .B2(n_957), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B1(n_586), .B2(n_589), .C(n_590), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g598 ( .A(n_583), .Y(n_598) );
INVx2_ASAP7_75t_L g697 ( .A(n_583), .Y(n_697) );
INVx3_ASAP7_75t_L g840 ( .A(n_583), .Y(n_840) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_588), .A2(n_590), .B1(n_746), .B2(n_749), .C(n_781), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_588), .A2(n_781), .B1(n_1067), .B2(n_1105), .C(n_1106), .Y(n_1104) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_588), .A2(n_840), .B1(n_851), .B2(n_1094), .C(n_1109), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1566 ( .A(n_588), .Y(n_1566) );
OAI221xp5_ASAP7_75t_L g839 ( .A1(n_590), .A2(n_817), .B1(n_819), .B2(n_840), .C(n_841), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g1020 ( .A1(n_590), .A2(n_840), .B1(n_993), .B2(n_997), .C(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_594), .A2(n_643), .B1(n_962), .B2(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g838 ( .A(n_596), .Y(n_838) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx3_ASAP7_75t_L g771 ( .A(n_601), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_601), .A2(n_603), .B1(n_949), .B2(n_950), .Y(n_948) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx3_ASAP7_75t_L g772 ( .A(n_603), .Y(n_772) );
OAI31xp33_ASAP7_75t_L g830 ( .A1(n_604), .A2(n_831), .A3(n_832), .B(n_843), .Y(n_830) );
OAI31xp33_ASAP7_75t_L g1014 ( .A1(n_604), .A2(n_1015), .A3(n_1016), .B(n_1024), .Y(n_1014) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
CKINVDCx8_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
XNOR2x1_ASAP7_75t_L g609 ( .A(n_610), .B(n_866), .Y(n_609) );
XNOR2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_726), .Y(n_610) );
XNOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_673), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_621), .C(n_624), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_638), .C(n_649), .D(n_656), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_634), .C(n_635), .Y(n_628) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g1267 ( .A(n_631), .Y(n_1267) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_635), .B(n_917), .C(n_918), .Y(n_916) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_646), .C(n_648), .Y(n_638) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g1019 ( .A(n_643), .Y(n_1019) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g779 ( .A(n_644), .Y(n_779) );
INVx2_ASAP7_75t_L g857 ( .A(n_644), .Y(n_857) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_645), .Y(n_792) );
INVx3_ASAP7_75t_L g914 ( .A(n_645), .Y(n_914) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_648), .B(n_908), .C(n_909), .Y(n_907) );
AOI33xp33_ASAP7_75t_L g1148 ( .A1(n_648), .A2(n_1149), .A3(n_1151), .B1(n_1155), .B2(n_1157), .B3(n_1160), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g707 ( .A(n_655), .Y(n_707) );
AOI31xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_667), .A3(n_670), .B(n_672), .Y(n_661) );
INVx1_ASAP7_75t_L g897 ( .A(n_665), .Y(n_897) );
AO21x1_ASAP7_75t_SL g693 ( .A1(n_672), .A2(n_694), .B(n_699), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g905 ( .A(n_672), .Y(n_905) );
AND4x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_693), .C(n_702), .D(n_711), .Y(n_674) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_675), .B(n_693), .C(n_702), .D(n_711), .Y(n_725) );
OAI31xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_684), .A3(n_687), .B(n_692), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .C(n_683), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
BUFx2_ASAP7_75t_L g745 ( .A(n_690), .Y(n_745) );
INVx1_ASAP7_75t_L g752 ( .A(n_690), .Y(n_752) );
INVx2_ASAP7_75t_L g804 ( .A(n_690), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_703), .B(n_911), .C(n_915), .Y(n_910) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_714), .A2(n_1004), .B1(n_1005), .B2(n_1007), .Y(n_1003) );
INVx1_ASAP7_75t_L g1121 ( .A(n_714), .Y(n_1121) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g723 ( .A(n_716), .Y(n_723) );
INVx1_ASAP7_75t_L g760 ( .A(n_716), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_807), .B2(n_865), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND4x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_767), .C(n_769), .D(n_799), .Y(n_729) );
NOR3xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .C(n_763), .Y(n_730) );
NOR3xp33_ASAP7_75t_SL g809 ( .A(n_731), .B(n_810), .C(n_827), .Y(n_809) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR3xp33_ASAP7_75t_SL g986 ( .A(n_732), .B(n_987), .C(n_1008), .Y(n_986) );
NOR3xp33_ASAP7_75t_L g1037 ( .A(n_732), .B(n_1038), .C(n_1058), .Y(n_1037) );
NOR3xp33_ASAP7_75t_SL g1583 ( .A(n_732), .B(n_1584), .C(n_1596), .Y(n_1583) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI33xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .A3(n_744), .B1(n_750), .B2(n_755), .B3(n_762), .Y(n_735) );
OAI33xp33_ASAP7_75t_L g810 ( .A1(n_736), .A2(n_762), .A3(n_811), .B1(n_816), .B2(n_820), .B3(n_824), .Y(n_810) );
INVx1_ASAP7_75t_SL g933 ( .A(n_736), .Y(n_933) );
OAI33xp33_ASAP7_75t_L g987 ( .A1(n_736), .A2(n_762), .A3(n_988), .B1(n_992), .B2(n_998), .B3(n_1003), .Y(n_987) );
OAI33xp33_ASAP7_75t_L g1038 ( .A1(n_736), .A2(n_1039), .A3(n_1043), .B1(n_1048), .B2(n_1052), .B3(n_1057), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1584 ( .A1(n_736), .A2(n_1585), .B1(n_1589), .B2(n_1590), .Y(n_1584) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B1(n_741), .B2(n_743), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g1039 ( .A1(n_738), .A2(n_1040), .B1(n_1041), .B2(n_1042), .Y(n_1039) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_739), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_740), .A2(n_743), .B1(n_775), .B2(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_749), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g816 ( .A1(n_745), .A2(n_817), .B1(n_818), .B2(n_819), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_745), .A2(n_1197), .B1(n_1200), .B2(n_1254), .C(n_1255), .Y(n_1253) );
OAI221xp5_ASAP7_75t_L g1585 ( .A1(n_745), .A2(n_1000), .B1(n_1586), .B2(n_1587), .C(n_1588), .Y(n_1585) );
OAI221xp5_ASAP7_75t_L g1590 ( .A1(n_745), .A2(n_1591), .B1(n_1592), .B2(n_1593), .C(n_1594), .Y(n_1590) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g880 ( .A(n_748), .Y(n_880) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .B1(n_759), .B2(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g812 ( .A(n_757), .Y(n_812) );
BUFx3_ASAP7_75t_L g1514 ( .A(n_757), .Y(n_1514) );
INVx2_ASAP7_75t_L g1523 ( .A(n_757), .Y(n_1523) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI31xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_773), .A3(n_784), .B(n_798), .Y(n_769) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g846 ( .A(n_781), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_781), .B(n_967), .Y(n_966) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_781), .A2(n_848), .B1(n_1044), .B2(n_1047), .C(n_1067), .Y(n_1066) );
BUFx3_ASAP7_75t_L g1553 ( .A(n_781), .Y(n_1553) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_789), .B1(n_790), .B2(n_793), .C(n_794), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_788), .Y(n_1225) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx3_ASAP7_75t_L g1113 ( .A(n_792), .Y(n_1113) );
INVx2_ASAP7_75t_L g1154 ( .A(n_792), .Y(n_1154) );
INVx2_ASAP7_75t_L g1603 ( .A(n_792), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g821 ( .A(n_804), .Y(n_821) );
INVx1_ASAP7_75t_L g865 ( .A(n_807), .Y(n_865) );
AND4x1_ASAP7_75t_L g808 ( .A(n_809), .B(n_828), .C(n_830), .D(n_862), .Y(n_808) );
OAI22xp33_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g988 ( .A1(n_812), .A2(n_989), .B1(n_990), .B2(n_991), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_813), .A2(n_815), .B1(n_834), .B2(n_837), .Y(n_833) );
INVx1_ASAP7_75t_L g1122 ( .A(n_814), .Y(n_1122) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_818), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_821), .A2(n_993), .B1(n_994), .B2(n_997), .Y(n_992) );
OAI22xp33_ASAP7_75t_L g998 ( .A1(n_821), .A2(n_999), .B1(n_1000), .B2(n_1002), .Y(n_998) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_821), .A2(n_1044), .B1(n_1045), .B2(n_1047), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_821), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1048) );
OAI22xp5_ASAP7_75t_SL g852 ( .A1(n_834), .A2(n_853), .B1(n_854), .B2(n_855), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_834), .A2(n_989), .B1(n_991), .B2(n_1018), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1600 ( .A1(n_834), .A2(n_1601), .B1(n_1602), .B2(n_1604), .Y(n_1600) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g1026 ( .A(n_835), .Y(n_1026) );
INVx2_ASAP7_75t_SL g1065 ( .A(n_835), .Y(n_1065) );
INVx2_ASAP7_75t_L g1609 ( .A(n_835), .Y(n_1609) );
BUFx3_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g1558 ( .A(n_836), .Y(n_1558) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g1221 ( .A(n_840), .Y(n_1221) );
BUFx2_ASAP7_75t_L g1218 ( .A(n_841), .Y(n_1218) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_847), .B1(n_848), .B2(n_850), .C(n_851), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1551 ( .A(n_849), .Y(n_1551) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OAI22x1_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B1(n_927), .B2(n_928), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g926 ( .A(n_872), .Y(n_926) );
AOI221x1_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_887), .B1(n_888), .B2(n_905), .C(n_906), .Y(n_872) );
NAND3xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_881), .C(n_884), .Y(n_873) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NAND4xp25_ASAP7_75t_SL g888 ( .A(n_889), .B(n_893), .C(n_902), .D(n_904), .Y(n_888) );
AOI222xp33_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_896), .B2(n_897), .C1(n_898), .C2(n_899), .Y(n_893) );
AND2x4_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_900), .A2(n_944), .B1(n_945), .B2(n_968), .Y(n_967) );
NAND4xp25_ASAP7_75t_L g906 ( .A(n_907), .B(n_910), .C(n_916), .D(n_919), .Y(n_906) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AND2x4_ASAP7_75t_L g1195 ( .A(n_914), .B(n_1196), .Y(n_1195) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_922), .C(n_924), .Y(n_919) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_SL g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NAND4xp75_ASAP7_75t_L g930 ( .A(n_931), .B(n_946), .C(n_973), .D(n_975), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_932), .B(n_943), .Y(n_931) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
OAI21xp5_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_958), .B(n_971), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_951), .Y(n_947) );
BUFx3_ASAP7_75t_L g1152 ( .A(n_953), .Y(n_1152) );
AND2x6_ASAP7_75t_L g1198 ( .A(n_955), .B(n_1196), .Y(n_1198) );
NAND2x1p5_ASAP7_75t_L g1214 ( .A(n_955), .B(n_1208), .Y(n_1214) );
NAND2x1_ASAP7_75t_SL g1207 ( .A(n_968), .B(n_1208), .Y(n_1207) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
OAI31xp33_ASAP7_75t_L g1061 ( .A1(n_971), .A2(n_1062), .A3(n_1063), .B(n_1068), .Y(n_1061) );
OAI31xp33_ASAP7_75t_L g1098 ( .A1(n_971), .A2(n_1099), .A3(n_1107), .B(n_1116), .Y(n_1098) );
OAI31xp33_ASAP7_75t_L g1597 ( .A1(n_971), .A2(n_1598), .A3(n_1599), .B(n_1607), .Y(n_1597) );
BUFx8_ASAP7_75t_SL g971 ( .A(n_972), .Y(n_971) );
INVx2_ASAP7_75t_L g1508 ( .A(n_972), .Y(n_1508) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
XNOR2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_1187), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1084), .B1(n_1185), .B2(n_1186), .Y(n_980) );
INVx1_ASAP7_75t_L g1185 ( .A(n_981), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_1034), .B1(n_1082), .B2(n_1083), .Y(n_981) );
INVx1_ASAP7_75t_L g1083 ( .A(n_982), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AND4x1_ASAP7_75t_L g985 ( .A(n_986), .B(n_1009), .C(n_1012), .D(n_1014), .Y(n_985) );
INVx1_ASAP7_75t_L g1252 ( .A(n_990), .Y(n_1252) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
BUFx2_ASAP7_75t_L g1592 ( .A(n_996), .Y(n_1592) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1001), .Y(n_1050) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1001), .Y(n_1254) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_1005), .A2(n_1053), .B1(n_1055), .B2(n_1056), .Y(n_1052) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_1006), .Y(n_1005) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1021 ( .A(n_1022), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_1023), .Y(n_1022) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_1030), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1201 ( .A(n_1030), .B(n_1196), .Y(n_1201) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1034), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
AND4x1_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1059), .C(n_1061), .D(n_1078), .Y(n_1036) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1054), .Y(n_1126) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_1065), .A2(n_1101), .B1(n_1102), .B2(n_1103), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1071), .B1(n_1072), .B2(n_1073), .C(n_1074), .Y(n_1069) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1070), .Y(n_1563) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_1072), .A2(n_1224), .B1(n_1225), .B2(n_1226), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1081), .Y(n_1078) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1084), .Y(n_1186) );
AO22x1_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1130), .B1(n_1183), .B2(n_1184), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1086), .Y(n_1184) );
NAND4xp75_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1096), .C(n_1098), .D(n_1117), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1092), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_1093), .A2(n_1111), .B1(n_1112), .B2(n_1114), .Y(n_1110) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1113), .Y(n_1564) );
AOI33xp33_ASAP7_75t_L g1117 ( .A1(n_1118), .A2(n_1119), .A3(n_1120), .B1(n_1123), .B2(n_1124), .B3(n_1129), .Y(n_1117) );
INVx2_ASAP7_75t_SL g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1589 ( .A(n_1129), .Y(n_1589) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1130), .Y(n_1183) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1132), .Y(n_1182) );
AOI211x1_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1145), .B(n_1147), .C(n_1173), .Y(n_1132) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1161), .Y(n_1147) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_1159), .A2(n_1225), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx3_ASAP7_75t_SL g1187 ( .A(n_1188), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1235), .Y(n_1189) );
NOR3xp33_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1204), .C(n_1215), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1199), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1194), .B1(n_1197), .B2(n_1198), .Y(n_1192) );
BUFx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1540 ( .A(n_1195), .Y(n_1540) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_1198), .A2(n_1539), .B1(n_1540), .B2(n_1541), .Y(n_1538) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_1200), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1542 ( .A1(n_1201), .A2(n_1543), .B1(n_1544), .B2(n_1545), .Y(n_1542) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx2_ASAP7_75t_SL g1547 ( .A(n_1206), .Y(n_1547) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
NAND2x1p5_ASAP7_75t_L g1211 ( .A(n_1208), .B(n_1212), .Y(n_1211) );
INVx3_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
BUFx4f_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
BUFx2_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
OAI33xp33_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1217), .A3(n_1223), .B1(n_1227), .B2(n_1230), .B3(n_1234), .Y(n_1215) );
OAI33xp33_ASAP7_75t_L g1548 ( .A1(n_1216), .A2(n_1234), .A3(n_1549), .B1(n_1554), .B2(n_1561), .B3(n_1565), .Y(n_1548) );
OAI22xp33_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1219), .B1(n_1220), .B2(n_1222), .Y(n_1217) );
OAI22xp33_ASAP7_75t_L g1230 ( .A1(n_1218), .A2(n_1231), .B1(n_1232), .B2(n_1233), .Y(n_1230) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1221), .Y(n_1232) );
AOI211xp5_ASAP7_75t_L g1242 ( .A1(n_1228), .A2(n_1243), .B(n_1245), .C(n_1251), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_1229), .A2(n_1231), .B1(n_1272), .B2(n_1274), .Y(n_1271) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_1233), .A2(n_1258), .B1(n_1261), .B2(n_1265), .C(n_1269), .Y(n_1257) );
AOI21xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1240), .B(n_1241), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1237), .Y(n_1535) );
AND2x4_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
AOI31xp33_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1257), .A3(n_1271), .B(n_1276), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1510 ( .A1(n_1243), .A2(n_1511), .B1(n_1513), .B2(n_1515), .C(n_1516), .Y(n_1510) );
INVx2_ASAP7_75t_SL g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1247), .Y(n_1517) );
INVx1_ASAP7_75t_SL g1270 ( .A(n_1250), .Y(n_1270) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
BUFx6f_ASAP7_75t_L g1527 ( .A(n_1260), .Y(n_1527) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_1272), .A2(n_1274), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
INVx6_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx4_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
OAI221xp5_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1502), .B1(n_1504), .B2(n_1568), .C(n_1572), .Y(n_1278) );
AND4x1_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1415), .C(n_1450), .D(n_1480), .Y(n_1279) );
A2O1A1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1367), .B(n_1368), .C(n_1399), .Y(n_1280) );
OAI211xp5_ASAP7_75t_SL g1281 ( .A1(n_1282), .A2(n_1315), .B(n_1346), .C(n_1349), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1305), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1283), .B(n_1364), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1283), .B(n_1306), .Y(n_1396) );
AND2x4_ASAP7_75t_SL g1491 ( .A(n_1283), .B(n_1305), .Y(n_1491) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_1284), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1284), .B(n_1305), .Y(n_1362) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1284), .Y(n_1367) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1285), .Y(n_1379) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1289), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1286), .B(n_1289), .Y(n_1308) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1287), .B(n_1289), .Y(n_1293) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1288), .B(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1290), .Y(n_1299) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1294 ( .A1(n_1295), .A2(n_1300), .B1(n_1301), .B2(n_1302), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g1327 ( .A1(n_1295), .A2(n_1303), .B1(n_1328), .B2(n_1329), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_1295), .A2(n_1303), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
BUFx3_ASAP7_75t_L g1382 ( .A(n_1295), .Y(n_1382) );
BUFx6f_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1297), .B(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1297), .Y(n_1312) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1298), .Y(n_1311) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1303), .Y(n_1385) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1304), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1305), .B(n_1341), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1305), .B(n_1365), .Y(n_1404) );
OAI221xp5_ASAP7_75t_L g1451 ( .A1(n_1305), .A2(n_1433), .B1(n_1452), .B2(n_1454), .C(n_1456), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1305), .B(n_1417), .Y(n_1459) );
CKINVDCx6p67_ASAP7_75t_R g1305 ( .A(n_1306), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1306), .B(n_1375), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1306), .B(n_1341), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1306), .B(n_1421), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g1467 ( .A1(n_1306), .A2(n_1347), .B1(n_1468), .B2(n_1471), .C(n_1473), .Y(n_1467) );
A2O1A1Ixp33_ASAP7_75t_L g1481 ( .A1(n_1306), .A2(n_1435), .B(n_1482), .C(n_1483), .Y(n_1481) );
AOI221xp5_ASAP7_75t_L g1483 ( .A1(n_1306), .A2(n_1374), .B1(n_1427), .B2(n_1484), .C(n_1485), .Y(n_1483) );
OR2x6_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1309), .Y(n_1306) );
AND2x4_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1312), .Y(n_1310) );
OAI21xp33_ASAP7_75t_SL g1619 ( .A1(n_1311), .A2(n_1576), .B(n_1620), .Y(n_1619) );
AND2x4_ASAP7_75t_L g1313 ( .A(n_1312), .B(n_1314), .Y(n_1313) );
AOI211xp5_ASAP7_75t_L g1315 ( .A1(n_1316), .A2(n_1324), .B(n_1335), .C(n_1339), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1316), .B(n_1394), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1316), .B(n_1337), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1316), .B(n_1325), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1320), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1317), .B(n_1337), .Y(n_1336) );
INVx4_ASAP7_75t_L g1344 ( .A(n_1317), .Y(n_1344) );
INVx3_ASAP7_75t_L g1357 ( .A(n_1317), .Y(n_1357) );
NOR2xp67_ASAP7_75t_SL g1409 ( .A(n_1317), .B(n_1410), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g1443 ( .A(n_1317), .B(n_1444), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1317), .B(n_1325), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1317), .B(n_1341), .Y(n_1493) );
AND2x4_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1320), .B(n_1348), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1320), .B(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1320), .B(n_1330), .Y(n_1410) );
NOR2xp33_ASAP7_75t_L g1418 ( .A(n_1320), .B(n_1330), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1464 ( .A(n_1320), .B(n_1465), .Y(n_1464) );
BUFx3_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1321), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1321), .B(n_1359), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1321), .B(n_1337), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1321), .B(n_1325), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1321), .B(n_1394), .Y(n_1431) );
OR2x2_ASAP7_75t_L g1479 ( .A(n_1321), .B(n_1448), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
AOI21xp33_ASAP7_75t_L g1412 ( .A1(n_1324), .A2(n_1413), .B(n_1414), .Y(n_1412) );
AOI21xp5_ASAP7_75t_L g1478 ( .A1(n_1324), .A2(n_1414), .B(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1325), .B(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1325), .B(n_1357), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1330), .Y(n_1325) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1326), .Y(n_1338) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1326), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1326), .B(n_1331), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1330), .B(n_1338), .Y(n_1345) );
INVx2_ASAP7_75t_L g1353 ( .A(n_1330), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1330), .B(n_1373), .Y(n_1477) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1331), .B(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1337), .B(n_1344), .Y(n_1348) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1337), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1337), .B(n_1372), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1345), .Y(n_1339) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1340), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1344), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g1365 ( .A(n_1341), .Y(n_1365) );
INVx1_ASAP7_75t_SL g1375 ( .A(n_1341), .Y(n_1375) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1341), .Y(n_1411) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1341), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1344), .B(n_1352), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1344), .B(n_1373), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1344), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1344), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1344), .B(n_1428), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1344), .B(n_1374), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1344), .B(n_1388), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1345), .B(n_1373), .Y(n_1434) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1345), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1345), .B(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_1348), .A2(n_1352), .B1(n_1402), .B2(n_1404), .C(n_1405), .Y(n_1401) );
A2O1A1Ixp33_ASAP7_75t_L g1349 ( .A1(n_1350), .A2(n_1353), .B(n_1354), .C(n_1360), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1352), .B(n_1393), .Y(n_1406) );
A2O1A1Ixp33_ASAP7_75t_L g1474 ( .A1(n_1352), .A2(n_1376), .B(n_1475), .C(n_1478), .Y(n_1474) );
INVxp67_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1358), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1356), .B(n_1404), .Y(n_1414) );
A2O1A1Ixp33_ASAP7_75t_L g1495 ( .A1(n_1356), .A2(n_1496), .B(n_1497), .C(n_1498), .Y(n_1495) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1357), .B(n_1425), .Y(n_1424) );
OR2x2_ASAP7_75t_L g1433 ( .A(n_1357), .B(n_1434), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1357), .B(n_1418), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1357), .B(n_1477), .Y(n_1476) );
NOR2x1_ASAP7_75t_L g1403 ( .A(n_1359), .B(n_1373), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1359), .B(n_1373), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1363), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1366), .Y(n_1363) );
AOI321xp33_ASAP7_75t_L g1415 ( .A1(n_1364), .A2(n_1374), .A3(n_1416), .B1(n_1419), .B2(n_1422), .C(n_1432), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1364), .B(n_1436), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1454 ( .A(n_1364), .B(n_1455), .Y(n_1454) );
INVx3_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1452 ( .A(n_1365), .B(n_1453), .Y(n_1452) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1365), .B(n_1491), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1366), .B(n_1377), .Y(n_1386) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_1366), .B(n_1377), .Y(n_1400) );
AOI21xp5_ASAP7_75t_SL g1480 ( .A1(n_1366), .A2(n_1481), .B(n_1489), .Y(n_1480) );
NOR3xp33_ASAP7_75t_L g1492 ( .A(n_1366), .B(n_1493), .C(n_1494), .Y(n_1492) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1367), .B(n_1388), .Y(n_1387) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1367), .Y(n_1430) );
INVxp67_ASAP7_75t_SL g1368 ( .A(n_1369), .Y(n_1368) );
OAI211xp5_ASAP7_75t_L g1399 ( .A1(n_1369), .A2(n_1400), .B(n_1401), .C(n_1407), .Y(n_1399) );
AOI221xp5_ASAP7_75t_L g1369 ( .A1(n_1370), .A2(n_1386), .B1(n_1387), .B2(n_1389), .C(n_1390), .Y(n_1369) );
OAI21xp33_ASAP7_75t_SL g1370 ( .A1(n_1371), .A2(n_1374), .B(n_1376), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1373), .B(n_1394), .Y(n_1428) );
OR2x2_ASAP7_75t_L g1469 ( .A(n_1373), .B(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1374), .Y(n_1461) );
A2O1A1Ixp33_ASAP7_75t_L g1422 ( .A1(n_1376), .A2(n_1423), .B(n_1426), .C(n_1429), .Y(n_1422) );
INVx2_ASAP7_75t_L g1445 ( .A(n_1376), .Y(n_1445) );
BUFx3_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1377), .Y(n_1421) );
AOI21xp5_ASAP7_75t_L g1437 ( .A1(n_1377), .A2(n_1438), .B(n_1439), .Y(n_1437) );
AOI31xp33_ASAP7_75t_L g1489 ( .A1(n_1377), .A2(n_1490), .A3(n_1495), .B(n_1499), .Y(n_1489) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
OAI22xp33_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1382), .B1(n_1383), .B2(n_1384), .Y(n_1380) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1382), .Y(n_1503) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1386), .Y(n_1462) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1387), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1387), .B(n_1398), .Y(n_1473) );
AOI21xp33_ASAP7_75t_L g1442 ( .A1(n_1388), .A2(n_1443), .B(n_1445), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1389), .B(n_1488), .Y(n_1487) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_1391), .A2(n_1392), .B1(n_1395), .B2(n_1397), .Y(n_1390) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1391), .Y(n_1498) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1394), .Y(n_1444) );
NAND2xp5_ASAP7_75t_SL g1471 ( .A(n_1395), .B(n_1472), .Y(n_1471) );
INVx2_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
AOI221xp5_ASAP7_75t_L g1490 ( .A1(n_1396), .A2(n_1408), .B1(n_1409), .B2(n_1491), .C(n_1492), .Y(n_1490) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
OAI21xp5_ASAP7_75t_L g1441 ( .A1(n_1402), .A2(n_1404), .B(n_1409), .Y(n_1441) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1403), .Y(n_1425) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
O2A1O1Ixp33_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1409), .B(n_1411), .C(n_1412), .Y(n_1407) );
NAND2xp5_ASAP7_75t_SL g1457 ( .A(n_1410), .B(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1411), .Y(n_1472) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1413), .Y(n_1496) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
AOI331xp33_ASAP7_75t_L g1432 ( .A1(n_1419), .A2(n_1433), .A3(n_1435), .B1(n_1437), .B2(n_1441), .B3(n_1442), .C1(n_1446), .Y(n_1432) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVxp67_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1428), .Y(n_1458) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1431), .Y(n_1429) );
NOR2xp33_ASAP7_75t_L g1460 ( .A(n_1434), .B(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
NOR2xp33_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1449), .Y(n_1447) );
AOI21xp5_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1462), .B(n_1463), .Y(n_1450) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1453), .Y(n_1482) );
AOI21xp5_ASAP7_75t_SL g1456 ( .A1(n_1457), .A2(n_1459), .B(n_1460), .Y(n_1456) );
OAI21xp33_ASAP7_75t_L g1485 ( .A1(n_1458), .A2(n_1486), .B(n_1487), .Y(n_1485) );
OAI211xp5_ASAP7_75t_SL g1463 ( .A1(n_1464), .A2(n_1466), .B(n_1467), .C(n_1474), .Y(n_1463) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1464), .Y(n_1484) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1479), .Y(n_1497) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_1503), .Y(n_1502) );
INVx2_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
XNOR2x1_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1567), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1536), .Y(n_1506) );
AOI22xp5_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1509), .B1(n_1534), .B2(n_1535), .Y(n_1507) );
NAND3xp33_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1520), .C(n_1531), .Y(n_1509) );
OAI22xp5_ASAP7_75t_L g1561 ( .A1(n_1515), .A2(n_1533), .B1(n_1562), .B2(n_1564), .Y(n_1561) );
INVx3_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
AOI221xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1526), .B1(n_1527), .B2(n_1528), .C(n_1529), .Y(n_1520) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
INVx3_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_1528), .A2(n_1532), .B1(n_1553), .B2(n_1566), .Y(n_1565) );
NOR3xp33_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1546), .C(n_1548), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1542), .Y(n_1537) );
OAI22xp33_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1551), .B1(n_1552), .B2(n_1553), .Y(n_1549) );
OAI21xp33_ASAP7_75t_L g1605 ( .A1(n_1553), .A2(n_1587), .B(n_1606), .Y(n_1605) );
OAI22xp5_ASAP7_75t_SL g1554 ( .A1(n_1555), .A2(n_1556), .B1(n_1559), .B2(n_1560), .Y(n_1554) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
INVx2_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
CKINVDCx5p33_ASAP7_75t_R g1574 ( .A(n_1575), .Y(n_1574) );
INVxp33_ASAP7_75t_SL g1577 ( .A(n_1578), .Y(n_1577) );
HB1xp67_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
AND4x1_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1583), .C(n_1597), .D(n_1616), .Y(n_1580) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1618), .Y(n_1616) );
endmodule