module fake_jpeg_11608_n_165 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_5),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_47),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_26),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_26),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_53),
.Y(n_74)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_14),
.Y(n_82)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_26),
.B1(n_24),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_67),
.B1(n_72),
.B2(n_66),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_60),
.B(n_73),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_27),
.B(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_12),
.B(n_14),
.C(n_6),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_12),
.B1(n_14),
.B2(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_7),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_12),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_14),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_76),
.Y(n_100)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_91),
.Y(n_106)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_34),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_69),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_75),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_60),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_73),
.B1(n_72),
.B2(n_66),
.Y(n_107)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_70),
.C(n_58),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_91),
.C(n_96),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_104),
.C(n_119),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_132),
.B(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_126),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_83),
.B1(n_100),
.B2(n_90),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_104),
.B(n_102),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_83),
.B(n_88),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_111),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_115),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_87),
.B(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_134),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_106),
.A3(n_108),
.B1(n_118),
.B2(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_136),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_108),
.A3(n_79),
.B1(n_85),
.B2(n_98),
.C1(n_111),
.C2(n_119),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_127),
.B(n_125),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_122),
.C(n_127),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_123),
.B(n_121),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_105),
.B1(n_61),
.B2(n_84),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_128),
.B1(n_105),
.B2(n_102),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_128),
.C(n_136),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_150),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_153),
.B1(n_142),
.B2(n_54),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_148),
.B1(n_71),
.B2(n_54),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_114),
.B1(n_103),
.B2(n_94),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_147),
.C(n_145),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_152),
.B(n_145),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_149),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_64),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_157),
.B(n_98),
.C(n_71),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_160),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_56),
.B(n_65),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_65),
.Y(n_165)
);


endmodule