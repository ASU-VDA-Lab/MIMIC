module fake_jpeg_13619_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_0),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_80),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_56),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_50),
.B1(n_24),
.B2(n_25),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_69),
.B1(n_62),
.B2(n_74),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_2),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_64),
.B(n_65),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_55),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_73),
.B1(n_62),
.B2(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_98),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_53),
.B1(n_69),
.B2(n_68),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_63),
.B(n_61),
.C(n_51),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_72),
.B(n_4),
.C(n_5),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_68),
.B1(n_61),
.B2(n_52),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_83),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_80),
.B1(n_55),
.B2(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_31),
.B1(n_46),
.B2(n_45),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_114),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_4),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_79),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_71),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_119),
.B(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_21),
.Y(n_128)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_3),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_5),
.B(n_6),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_85),
.B(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_140),
.B(n_14),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_72),
.A3(n_27),
.B1(n_29),
.B2(n_49),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_126),
.B1(n_130),
.B2(n_16),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_38),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_129),
.Y(n_146)
);

OAI22x1_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_112),
.B1(n_106),
.B2(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_136),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_15),
.B(n_16),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_7),
.B(n_10),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_144),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_149),
.B(n_150),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_152),
.B(n_137),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_122),
.A3(n_139),
.B1(n_140),
.B2(n_121),
.C1(n_47),
.C2(n_44),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_30),
.B(n_34),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_153),
.C(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_36),
.B(n_37),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_123),
.A3(n_121),
.B1(n_127),
.B2(n_133),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_143),
.B1(n_151),
.B2(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_163),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_141),
.B(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_156),
.C(n_154),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_158),
.B1(n_159),
.B2(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_165),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_41),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_43),
.B(n_133),
.Y(n_170)
);


endmodule