module fake_jpeg_20061_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_6),
.B(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_54),
.B1(n_65),
.B2(n_44),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_19),
.B(n_15),
.C(n_17),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_32),
.B1(n_18),
.B2(n_27),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_24),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_38),
.B(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_72),
.B1(n_95),
.B2(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_96),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_29),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_75),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_41),
.B1(n_40),
.B2(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_80),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_43),
.B1(n_20),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_97),
.B1(n_61),
.B2(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_85),
.Y(n_117)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_83),
.B(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_54),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_29),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_88),
.Y(n_125)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_38),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_0),
.B(n_1),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_98),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_42),
.B1(n_39),
.B2(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_38),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_51),
.B(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_22),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_22),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_1),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.C(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_62),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_105),
.B(n_131),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_61),
.B1(n_56),
.B2(n_4),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_79),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_112),
.A2(n_122),
.B1(n_123),
.B2(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_61),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_2),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_82),
.B1(n_13),
.B2(n_74),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_68),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_83),
.B1(n_101),
.B2(n_82),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_135),
.B1(n_97),
.B2(n_91),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_72),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_12),
.B1(n_13),
.B2(n_102),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_144),
.B1(n_155),
.B2(n_156),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_147),
.B(n_124),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_92),
.B1(n_88),
.B2(n_94),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_104),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_160),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_109),
.B(n_134),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_145),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_78),
.C(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_124),
.C(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_136),
.B1(n_118),
.B2(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_118),
.B1(n_111),
.B2(n_116),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_116),
.B1(n_130),
.B2(n_121),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_107),
.B1(n_163),
.B2(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_170),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_178),
.C(n_144),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_184),
.B(n_138),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_108),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_186),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_106),
.C(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_107),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_185),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_156),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_143),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_163),
.B1(n_141),
.B2(n_155),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_195),
.B1(n_184),
.B2(n_165),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_147),
.B(n_148),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_203),
.B(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_149),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_181),
.B1(n_173),
.B2(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_165),
.B1(n_178),
.B2(n_168),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_138),
.B(n_142),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_164),
.B(n_170),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_205),
.C(n_166),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_140),
.B(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_140),
.C(n_161),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_216),
.C(n_220),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_221),
.B1(n_196),
.B2(n_197),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_176),
.C(n_168),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_199),
.C(n_200),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_191),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_199),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_195),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_188),
.B1(n_194),
.B2(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_233),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_189),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_215),
.B1(n_209),
.B2(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_221),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_222),
.C(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_218),
.B1(n_213),
.B2(n_192),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_227),
.B(n_213),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_236),
.B(n_201),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_237),
.C(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_252),
.A2(n_244),
.B(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_238),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_259),
.B(n_256),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_237),
.Y(n_262)
);


endmodule