module fake_jpeg_1912_n_294 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_44),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_45),
.B(n_48),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_7),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_10),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_10),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_5),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_11),
.C(n_14),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_84),
.Y(n_109)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_25),
.B1(n_38),
.B2(n_27),
.Y(n_98)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_2),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_26),
.B1(n_33),
.B2(n_39),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_91),
.A2(n_122),
.B1(n_128),
.B2(n_101),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_106),
.B1(n_115),
.B2(n_124),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_19),
.B1(n_39),
.B2(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_33),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_38),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_126),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_52),
.A2(n_33),
.B1(n_73),
.B2(n_80),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_130),
.B1(n_89),
.B2(n_93),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_47),
.B(n_13),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_95),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_1),
.B1(n_13),
.B2(n_14),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_59),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_15),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_74),
.A2(n_63),
.B1(n_82),
.B2(n_44),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_111),
.B1(n_120),
.B2(n_132),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_94),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_142),
.Y(n_183)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_57),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_94),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_143),
.B(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_151),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_105),
.B(n_102),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_146),
.B(n_163),
.Y(n_200)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_51),
.B1(n_56),
.B2(n_62),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_166),
.B1(n_171),
.B2(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_57),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_88),
.A2(n_75),
.B(n_79),
.C(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_87),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_79),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_159),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_85),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_162),
.Y(n_197)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_123),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_110),
.A2(n_128),
.B(n_108),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_176),
.Y(n_206)
);

NAND2x1_ASAP7_75t_SL g170 ( 
.A(n_93),
.B(n_118),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_130),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_141),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_132),
.B1(n_116),
.B2(n_96),
.Y(n_177)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_178),
.B1(n_182),
.B2(n_205),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_87),
.B1(n_96),
.B2(n_107),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_186),
.A2(n_139),
.B1(n_138),
.B2(n_148),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_192),
.C(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_140),
.B(n_96),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_203),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_107),
.B1(n_147),
.B2(n_155),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_149),
.B1(n_154),
.B2(n_162),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_136),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_140),
.B(n_107),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_146),
.B1(n_172),
.B2(n_141),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_152),
.B1(n_159),
.B2(n_157),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_205),
.B1(n_188),
.B2(n_194),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_143),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_211),
.B(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_219),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_150),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_174),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_227),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_175),
.C(n_149),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_204),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_149),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_145),
.B(n_161),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_185),
.B(n_199),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_207),
.B1(n_194),
.B2(n_190),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_196),
.A2(n_186),
.B1(n_187),
.B2(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_200),
.C(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_224),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_201),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_182),
.C(n_183),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_183),
.B(n_195),
.C(n_177),
.D(n_185),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_239),
.B(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_181),
.B1(n_198),
.B2(n_195),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_236),
.B1(n_204),
.B2(n_223),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_181),
.B1(n_198),
.B2(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_215),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_228),
.A3(n_224),
.B1(n_210),
.B2(n_222),
.C1(n_209),
.C2(n_225),
.Y(n_245)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_180),
.B1(n_231),
.B2(n_247),
.C(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_226),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_212),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_217),
.B1(n_219),
.B2(n_230),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_234),
.B1(n_245),
.B2(n_242),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_239),
.B(n_238),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_259),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_180),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.C(n_260),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_180),
.C(n_247),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_231),
.C(n_234),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_240),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_257),
.C(n_260),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_252),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_264),
.Y(n_281)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_246),
.B1(n_236),
.B2(n_238),
.Y(n_275)
);

OAI321xp33_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_262),
.A3(n_251),
.B1(n_255),
.B2(n_246),
.C(n_253),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_277),
.A2(n_261),
.B1(n_262),
.B2(n_254),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_232),
.B(n_276),
.Y(n_285)
);

AOI221xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_277),
.B1(n_255),
.B2(n_239),
.C(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_276),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_285),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_286),
.A2(n_278),
.B(n_232),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_265),
.B(n_266),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_290),
.A2(n_291),
.B1(n_289),
.B2(n_282),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_293),
.CI(n_285),
.CON(n_294),
.SN(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_289),
.C(n_236),
.Y(n_293)
);


endmodule