module fake_aes_12001_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx4_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVxp33_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_12), .B(n_2), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_12), .B(n_2), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_13), .B(n_3), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
OAI21x1_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_16), .B(n_14), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_21), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
AOI31xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_13), .A3(n_22), .B(n_20), .Y(n_27) );
AOI21xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_23), .B(n_17), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_15), .B1(n_16), .B2(n_14), .Y(n_29) );
A2O1A1Ixp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_27), .B(n_23), .C(n_12), .Y(n_30) );
AO221x1_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_27), .B1(n_12), .B2(n_5), .C(n_6), .Y(n_31) );
OAI221xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_23), .B1(n_4), .B2(n_6), .C(n_7), .Y(n_32) );
AND2x4_ASAP7_75t_L g33 ( .A(n_30), .B(n_9), .Y(n_33) );
NAND2x1p5_ASAP7_75t_L g34 ( .A(n_31), .B(n_3), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_32), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_35), .B(n_7), .Y(n_36) );
NOR3xp33_ASAP7_75t_L g37 ( .A(n_33), .B(n_8), .C(n_10), .Y(n_37) );
OAI31xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_34), .A3(n_33), .B(n_8), .Y(n_38) );
AOI22xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_33), .B1(n_34), .B2(n_36), .Y(n_39) );
endmodule