module fake_netlist_6_760_n_1661 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1661);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1661;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_25),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_74),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_9),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_27),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_75),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_41),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_67),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_64),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_9),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_42),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_22),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_21),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_43),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_21),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_30),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_104),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_27),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_19),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_58),
.Y(n_195)
);

BUFx8_ASAP7_75t_SL g196 ( 
.A(n_50),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_40),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_131),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_16),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_85),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_14),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_47),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_26),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_44),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_103),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_51),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_59),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_12),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_12),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_62),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_35),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_48),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_63),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_88),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_87),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_51),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_125),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_108),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_35),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_28),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_73),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_83),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_25),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_81),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_55),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_52),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_31),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_55),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_80),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_78),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_127),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_13),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_110),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_0),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_0),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_24),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_23),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_48),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_39),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_45),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_82),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_90),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_68),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_56),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_146),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_20),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_116),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_84),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_86),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_124),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_19),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_121),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_57),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_16),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_54),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_8),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_130),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_61),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_42),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_34),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_91),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_41),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_105),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_29),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_10),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_148),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_139),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_65),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_93),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_23),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_17),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_71),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_4),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_53),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_11),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_1),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_30),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_203),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_196),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_203),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_173),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_153),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_176),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_161),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_1),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_203),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_156),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_159),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_232),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_166),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_170),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_158),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_2),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_172),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_158),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_177),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_158),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_197),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_197),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_197),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_224),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_224),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_157),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_163),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_157),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_171),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_171),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_212),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_217),
.B(n_2),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_276),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_186),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_173),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_189),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_181),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_181),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_288),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_192),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_182),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_182),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_183),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_194),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_183),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_162),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_206),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_190),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_190),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_193),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_208),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_210),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_193),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_276),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_214),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_198),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_221),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_276),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_225),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_228),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_240),
.B(n_3),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_230),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_236),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_240),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_358),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_176),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

BUFx8_ASAP7_75t_L g384 ( 
.A(n_322),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_311),
.B(n_176),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_306),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_306),
.B(n_234),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_312),
.B(n_175),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_338),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_313),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_314),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_314),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_238),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_234),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_341),
.B(n_304),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_348),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_322),
.B(n_234),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_346),
.A2(n_184),
.B1(n_258),
.B2(n_301),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_325),
.B(n_327),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_325),
.B(n_247),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_320),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g431 ( 
.A(n_329),
.B(n_250),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_329),
.B(n_248),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_345),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_330),
.B(n_250),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_351),
.B(n_261),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_400),
.A2(n_280),
.B1(n_368),
.B2(n_216),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_250),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_415),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_331),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_400),
.B(n_310),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_415),
.B(n_315),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_422),
.B(n_316),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_422),
.B(n_319),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_321),
.Y(n_464)
);

OAI21xp33_ASAP7_75t_SL g465 ( 
.A1(n_411),
.A2(n_368),
.B(n_249),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_403),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_410),
.A2(n_222),
.B1(n_249),
.B2(n_253),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_435),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

OAI21xp33_ASAP7_75t_SL g472 ( 
.A1(n_411),
.A2(n_253),
.B(n_222),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_403),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_435),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_410),
.B(n_331),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_378),
.A2(n_255),
.B1(n_256),
.B2(n_259),
.Y(n_482)
);

CKINVDCx6p67_ASAP7_75t_R g483 ( 
.A(n_386),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_324),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_427),
.B(n_326),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_328),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_382),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_382),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_386),
.Y(n_494)
);

OR2x2_ASAP7_75t_SL g495 ( 
.A(n_378),
.B(n_255),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_343),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_433),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_441),
.B(n_355),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_425),
.B(n_154),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_390),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_381),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_439),
.A2(n_267),
.B1(n_256),
.B2(n_259),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_388),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_379),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_359),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_390),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_418),
.B(n_364),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_381),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_418),
.B(n_367),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_420),
.B(n_369),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_388),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_397),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_420),
.B(n_373),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_426),
.B(n_376),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_426),
.B(n_375),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_L g519 ( 
.A(n_390),
.B(n_333),
.C(n_332),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_381),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_426),
.B(n_350),
.Y(n_521)
);

BUFx6f_ASAP7_75t_SL g522 ( 
.A(n_439),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_382),
.B(n_162),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_393),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_397),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_418),
.B(n_188),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_381),
.B(n_209),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_384),
.B(n_356),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_396),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_397),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_384),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_403),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_381),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_379),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_398),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_403),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_403),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_398),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_399),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_439),
.B(n_154),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_384),
.B(n_372),
.Y(n_545)
);

CKINVDCx6p67_ASAP7_75t_R g546 ( 
.A(n_439),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_407),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_439),
.B(n_332),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_421),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_399),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_421),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_402),
.B(n_363),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_407),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_384),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_384),
.B(n_307),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_380),
.Y(n_558)
);

BUFx8_ASAP7_75t_SL g559 ( 
.A(n_392),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_404),
.B(n_334),
.C(n_333),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_385),
.B(n_294),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_405),
.B(n_406),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_405),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_407),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_385),
.B(n_334),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_392),
.A2(n_263),
.B1(n_267),
.B2(n_277),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_406),
.B(n_360),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_408),
.B(n_413),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_407),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_392),
.A2(n_205),
.B1(n_160),
.B2(n_246),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_408),
.A2(n_207),
.B1(n_223),
.B2(n_219),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_385),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_407),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_413),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_382),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_392),
.A2(n_263),
.B1(n_277),
.B2(n_281),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_407),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_392),
.A2(n_281),
.B1(n_302),
.B2(n_297),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_414),
.A2(n_285),
.B1(n_290),
.B2(n_297),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_414),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_416),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_440),
.B(n_252),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_416),
.B(n_419),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_382),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_419),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_430),
.A2(n_285),
.B1(n_290),
.B2(n_302),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_R g589 ( 
.A(n_475),
.B(n_336),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_499),
.B(n_453),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_499),
.B(n_440),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_447),
.A2(n_431),
.B1(n_440),
.B2(n_227),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_570),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_449),
.B(n_162),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_484),
.B(n_440),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_483),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_570),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_502),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_464),
.B(n_440),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_451),
.B(n_340),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_563),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_451),
.B(n_430),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_585),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_488),
.B(n_440),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_447),
.A2(n_431),
.B1(n_440),
.B2(n_284),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_585),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_489),
.B(n_180),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_496),
.B(n_394),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_508),
.A2(n_273),
.B1(n_265),
.B2(n_266),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_483),
.B(n_261),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_449),
.B(n_162),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_465),
.A2(n_282),
.B1(n_268),
.B2(n_271),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_502),
.B(n_436),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_452),
.B(n_394),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_449),
.B(n_450),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_516),
.B(n_164),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_452),
.B(n_394),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_449),
.B(n_162),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_509),
.B(n_436),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_450),
.B(n_162),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_568),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_477),
.B(n_394),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_477),
.B(n_394),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_510),
.B(n_512),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_509),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_448),
.B(n_437),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_448),
.B(n_437),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_447),
.A2(n_431),
.B1(n_284),
.B2(n_211),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_456),
.B(n_437),
.Y(n_633)
);

BUFx5_ASAP7_75t_L g634 ( 
.A(n_492),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_456),
.B(n_437),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_554),
.B(n_168),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_506),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_514),
.Y(n_639)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_522),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_549),
.B(n_438),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_514),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_458),
.B(n_431),
.Y(n_643)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_465),
.A2(n_211),
.B(n_292),
.C(n_274),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_445),
.B(n_185),
.C(n_174),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_450),
.B(n_220),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_517),
.B(n_187),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_458),
.B(n_431),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_470),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_525),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_459),
.B(n_191),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_553),
.B(n_220),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_478),
.B(n_220),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_469),
.B(n_431),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_469),
.B(n_431),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_471),
.B(n_431),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_460),
.B(n_195),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_478),
.B(n_220),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_462),
.B(n_200),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_497),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_471),
.B(n_473),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_478),
.B(n_220),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_513),
.B(n_202),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_519),
.B(n_218),
.C(n_305),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_478),
.B(n_272),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_495),
.B(n_438),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_524),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_560),
.B(n_261),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_498),
.B(n_287),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_447),
.A2(n_431),
.B1(n_274),
.B2(n_270),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_360),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_560),
.B(n_213),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_498),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_534),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_524),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_473),
.B(n_431),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_494),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_530),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_476),
.B(n_431),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_472),
.A2(n_500),
.B1(n_526),
.B2(n_546),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_455),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_476),
.B(n_385),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_505),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_530),
.B(n_155),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_564),
.B(n_261),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_531),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_531),
.B(n_533),
.Y(n_687)
);

AO22x2_ASAP7_75t_L g688 ( 
.A1(n_528),
.A2(n_179),
.B1(n_155),
.B2(n_165),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_472),
.B(n_289),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_573),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_533),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_455),
.B(n_295),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_546),
.A2(n_296),
.B1(n_300),
.B2(n_237),
.Y(n_693)
);

NOR3xp33_ASAP7_75t_L g694 ( 
.A(n_518),
.B(n_254),
.C(n_215),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_539),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_539),
.B(n_165),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_542),
.B(n_380),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_542),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_535),
.B(n_382),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_543),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_167),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_551),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_229),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_552),
.B(n_380),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_552),
.B(n_167),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_482),
.A2(n_169),
.B1(n_179),
.B2(n_201),
.C(n_204),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_447),
.A2(n_169),
.B1(n_201),
.B2(n_292),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_576),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_549),
.A2(n_204),
.B1(n_226),
.B2(n_270),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_576),
.B(n_226),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_521),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_503),
.Y(n_713)
);

NOR2x1p5_ASAP7_75t_L g714 ( 
.A(n_515),
.B(n_233),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_582),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_582),
.B(n_227),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_583),
.B(n_231),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_583),
.B(n_231),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_494),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_587),
.B(n_237),
.Y(n_720)
);

AND2x4_ASAP7_75t_SL g721 ( 
.A(n_494),
.B(n_535),
.Y(n_721)
);

AOI22x1_ASAP7_75t_L g722 ( 
.A1(n_511),
.A2(n_262),
.B1(n_362),
.B2(n_365),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_587),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_494),
.B(n_298),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_501),
.A2(n_262),
.B1(n_387),
.B2(n_382),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_550),
.B(n_235),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_SL g727 ( 
.A(n_467),
.B(n_239),
.Y(n_727)
);

BUFx5_ASAP7_75t_L g728 ( 
.A(n_503),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_503),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_527),
.B(n_387),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_562),
.B(n_380),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_501),
.A2(n_387),
.B1(n_382),
.B2(n_423),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_520),
.B(n_537),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_544),
.B(n_361),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_520),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_572),
.B(n_298),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_572),
.B(n_241),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_520),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_490),
.B(n_380),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_553),
.B(n_557),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_545),
.B(n_361),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_561),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_537),
.B(n_387),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_537),
.B(n_387),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_490),
.B(n_380),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_501),
.B(n_298),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_574),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_574),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_566),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_574),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_544),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_559),
.B(n_242),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_556),
.A2(n_303),
.B1(n_244),
.B2(n_245),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_463),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_490),
.B(n_380),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_628),
.A2(n_556),
.B1(n_501),
.B2(n_522),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_601),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_668),
.B(n_501),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_652),
.B(n_490),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_652),
.B(n_680),
.Y(n_760)
);

CKINVDCx6p67_ASAP7_75t_R g761 ( 
.A(n_603),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_629),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_619),
.A2(n_595),
.B(n_602),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_590),
.B(n_490),
.Y(n_764)
);

NOR2x1p5_ASAP7_75t_L g765 ( 
.A(n_736),
.B(n_243),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_598),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_607),
.A2(n_457),
.B(n_443),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_637),
.B(n_257),
.C(n_251),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_590),
.A2(n_522),
.B1(n_544),
.B2(n_504),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_620),
.B(n_544),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_611),
.B(n_490),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_650),
.B(n_544),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_712),
.B(n_584),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_610),
.A2(n_567),
.B(n_578),
.C(n_580),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_591),
.A2(n_479),
.B(n_538),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_634),
.B(n_491),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_733),
.A2(n_479),
.B(n_538),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_644),
.A2(n_523),
.B(n_581),
.C(n_588),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_647),
.B(n_468),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_605),
.B(n_468),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_740),
.A2(n_474),
.B(n_466),
.C(n_575),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_599),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_644),
.A2(n_536),
.B(n_579),
.C(n_529),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_589),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_731),
.A2(n_538),
.B(n_457),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_616),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_731),
.A2(n_538),
.B(n_457),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_636),
.B(n_468),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_649),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_690),
.B(n_522),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_617),
.A2(n_457),
.B(n_538),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_638),
.B(n_468),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_639),
.B(n_480),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_621),
.A2(n_538),
.B(n_457),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_642),
.B(n_480),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_600),
.B(n_362),
.Y(n_796)
);

AO21x1_ASAP7_75t_L g797 ( 
.A1(n_689),
.A2(n_669),
.B(n_661),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_726),
.B(n_480),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_589),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_626),
.A2(n_443),
.B(n_479),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_634),
.B(n_491),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_627),
.A2(n_443),
.B(n_479),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_685),
.B(n_298),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_640),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_665),
.A2(n_443),
.B(n_479),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_480),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_675),
.B(n_481),
.Y(n_807)
);

AO21x2_ASAP7_75t_L g808 ( 
.A1(n_665),
.A2(n_540),
.B(n_579),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_730),
.A2(n_443),
.B(n_479),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_737),
.A2(n_663),
.B(n_657),
.C(n_659),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_594),
.A2(n_481),
.B(n_507),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_682),
.A2(n_558),
.B(n_443),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_707),
.A2(n_529),
.B(n_579),
.C(n_532),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_594),
.A2(n_481),
.B(n_507),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_678),
.B(n_481),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_695),
.B(n_507),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_614),
.A2(n_507),
.B(n_442),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_672),
.B(n_260),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_709),
.B(n_558),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_687),
.A2(n_558),
.B(n_577),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_715),
.B(n_558),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_SL g822 ( 
.A1(n_643),
.A2(n_529),
.B(n_565),
.C(n_555),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_SL g823 ( 
.A(n_596),
.B(n_269),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_614),
.A2(n_558),
.B(n_577),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_704),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_622),
.A2(n_586),
.B(n_577),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_624),
.A2(n_586),
.B(n_577),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_604),
.A2(n_569),
.B1(n_444),
.B2(n_487),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_641),
.A2(n_569),
.B1(n_463),
.B2(n_575),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_624),
.A2(n_586),
.B(n_577),
.Y(n_830)
);

O2A1O1Ixp5_ASAP7_75t_L g831 ( 
.A1(n_669),
.A2(n_444),
.B(n_442),
.C(n_446),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_641),
.B(n_442),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_646),
.A2(n_658),
.B(n_653),
.Y(n_833)
);

AO21x1_ASAP7_75t_L g834 ( 
.A1(n_689),
.A2(n_571),
.B(n_466),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_599),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_641),
.B(n_444),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_606),
.B(n_365),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_623),
.B(n_446),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_609),
.B(n_446),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_686),
.B(n_454),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_686),
.B(n_454),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_651),
.A2(n_666),
.B(n_618),
.C(n_625),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_691),
.B(n_454),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_660),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_653),
.A2(n_491),
.B(n_461),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_658),
.A2(n_487),
.B(n_461),
.Y(n_846)
);

AO21x1_ASAP7_75t_L g847 ( 
.A1(n_662),
.A2(n_696),
.B(n_684),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_599),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_662),
.A2(n_487),
.B(n_461),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_749),
.A2(n_486),
.B(n_493),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_697),
.A2(n_486),
.B(n_493),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_640),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_SL g853 ( 
.A(n_596),
.B(n_275),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_673),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_593),
.A2(n_569),
.B1(n_486),
.B2(n_493),
.Y(n_855)
);

O2A1O1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_597),
.A2(n_541),
.B(n_532),
.C(n_565),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_699),
.A2(n_571),
.B(n_474),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_671),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_734),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_691),
.A2(n_569),
.B1(n_547),
.B2(n_548),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_683),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_719),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_699),
.A2(n_547),
.B(n_548),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_742),
.A2(n_717),
.B(n_720),
.C(n_718),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_724),
.B(n_278),
.Y(n_865)
);

NOR2x1_ASAP7_75t_L g866 ( 
.A(n_714),
.B(n_532),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_640),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_751),
.A2(n_565),
.B1(n_555),
.B2(n_541),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_698),
.A2(n_555),
.B1(n_541),
.B2(n_540),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_677),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_630),
.A2(n_540),
.B(n_536),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_698),
.B(n_536),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_702),
.A2(n_371),
.B(n_377),
.C(n_412),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_631),
.A2(n_383),
.B(n_380),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_674),
.B(n_279),
.C(n_283),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_633),
.A2(n_635),
.B(n_743),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_734),
.B(n_371),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_407),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_744),
.A2(n_383),
.B(n_377),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_746),
.B(n_286),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_729),
.A2(n_383),
.B(n_377),
.Y(n_881)
);

NOR2x1_ASAP7_75t_L g882 ( 
.A(n_664),
.B(n_391),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_701),
.A2(n_291),
.B1(n_293),
.B2(n_299),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_734),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_683),
.Y(n_885)
);

BUFx4f_ASAP7_75t_L g886 ( 
.A(n_741),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_741),
.B(n_5),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_634),
.B(n_383),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_701),
.B(n_417),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_612),
.B(n_69),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_729),
.A2(n_383),
.B(n_424),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_752),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_735),
.A2(n_748),
.B(n_747),
.Y(n_893)
);

AOI21x1_ASAP7_75t_L g894 ( 
.A1(n_697),
.A2(n_428),
.B(n_424),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_735),
.A2(n_428),
.B(n_424),
.Y(n_895)
);

AO21x1_ASAP7_75t_L g896 ( 
.A1(n_706),
.A2(n_428),
.B(n_424),
.Y(n_896)
);

NOR2x1_ASAP7_75t_R g897 ( 
.A(n_613),
.B(n_423),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_738),
.A2(n_428),
.B(n_391),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_694),
.B(n_412),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_615),
.A2(n_412),
.B(n_401),
.C(n_395),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_5),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_723),
.B(n_423),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_738),
.A2(n_412),
.B(n_401),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_747),
.A2(n_401),
.B(n_395),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_748),
.A2(n_401),
.B(n_395),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_634),
.B(n_423),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_648),
.A2(n_387),
.B(n_395),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_741),
.B(n_11),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_654),
.A2(n_391),
.B(n_417),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_723),
.B(n_423),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_599),
.B(n_423),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_708),
.A2(n_681),
.B1(n_750),
.B2(n_693),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_681),
.B(n_423),
.Y(n_914)
);

AOI33xp33_ASAP7_75t_L g915 ( 
.A1(n_710),
.A2(n_391),
.A3(n_15),
.B1(n_17),
.B2(n_20),
.B3(n_22),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_681),
.B(n_417),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_727),
.A2(n_417),
.B(n_387),
.C(n_26),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_681),
.B(n_66),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_713),
.B(n_417),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_713),
.A2(n_417),
.B1(n_387),
.B2(n_76),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_754),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_640),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_692),
.A2(n_387),
.B1(n_417),
.B2(n_152),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_810),
.B(n_645),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_763),
.A2(n_713),
.B(n_692),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_770),
.B(n_728),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_818),
.A2(n_727),
.B(n_721),
.C(n_711),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_757),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_818),
.A2(n_753),
.B(n_688),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_762),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_770),
.A2(n_721),
.B(n_716),
.C(n_679),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_786),
.B(n_688),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_760),
.A2(n_705),
.B(n_656),
.C(n_655),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_786),
.B(n_688),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_773),
.A2(n_676),
.B(n_754),
.C(n_705),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_760),
.A2(n_713),
.B1(n_608),
.B2(n_592),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_825),
.B(n_728),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_766),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_842),
.A2(n_632),
.B(n_670),
.C(n_739),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_773),
.B(n_728),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_774),
.A2(n_725),
.B(n_732),
.C(n_739),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_887),
.A2(n_755),
.B(n_745),
.C(n_722),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_779),
.A2(n_755),
.B(n_745),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_758),
.B(n_798),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_865),
.A2(n_14),
.B(n_24),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_859),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_858),
.B(n_880),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_798),
.B(n_728),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_835),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_759),
.A2(n_728),
.B1(n_92),
.B2(n_97),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_880),
.A2(n_790),
.B(n_864),
.C(n_865),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_799),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_833),
.A2(n_728),
.B(n_387),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_797),
.B(n_728),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_877),
.B(n_151),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_766),
.Y(n_957)
);

NAND2x1_ASAP7_75t_L g958 ( 
.A(n_922),
.B(n_387),
.Y(n_958)
);

AOI222xp33_ASAP7_75t_L g959 ( 
.A1(n_887),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_790),
.B(n_149),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_902),
.A2(n_32),
.B(n_34),
.C(n_36),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_767),
.A2(n_98),
.B(n_145),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_902),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_909),
.A2(n_38),
.B(n_43),
.C(n_45),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_909),
.A2(n_46),
.B(n_47),
.C(n_49),
.Y(n_965)
);

AO22x1_ASAP7_75t_L g966 ( 
.A1(n_768),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_966)
);

O2A1O1Ixp5_ASAP7_75t_L g967 ( 
.A1(n_896),
.A2(n_109),
.B(n_129),
.C(n_126),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_777),
.A2(n_876),
.B(n_805),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_L g969 ( 
.A(n_892),
.B(n_100),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_886),
.B(n_101),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_886),
.B(n_99),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_838),
.A2(n_111),
.B(n_117),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_918),
.B(n_832),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_803),
.B(n_52),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_789),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_877),
.B(n_796),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_856),
.A2(n_114),
.B(n_115),
.C(n_147),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_862),
.B(n_784),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_796),
.B(n_837),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_859),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_844),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_917),
.A2(n_60),
.B(n_759),
.C(n_875),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_809),
.A2(n_60),
.B(n_791),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_847),
.A2(n_834),
.B(n_756),
.C(n_781),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_794),
.A2(n_800),
.B(n_802),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_883),
.A2(n_913),
.B(n_772),
.C(n_839),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_837),
.B(n_780),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_761),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_884),
.B(n_898),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_775),
.A2(n_801),
.B(n_776),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_SL g991 ( 
.A(n_823),
.B(n_853),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_804),
.B(n_852),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_804),
.Y(n_993)
);

AO32x1_ASAP7_75t_L g994 ( 
.A1(n_855),
.A2(n_869),
.A3(n_828),
.B1(n_860),
.B2(n_900),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_884),
.Y(n_995)
);

AO21x2_ASAP7_75t_L g996 ( 
.A1(n_822),
.A2(n_808),
.B(n_787),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_835),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_L g998 ( 
.A1(n_769),
.A2(n_836),
.B(n_897),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_890),
.A2(n_854),
.B1(n_885),
.B2(n_861),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_921),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_870),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_764),
.B(n_788),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_SL g1003 ( 
.A1(n_918),
.A2(n_765),
.B1(n_866),
.B2(n_782),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_848),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_893),
.A2(n_783),
.B(n_831),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_804),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_829),
.A2(n_821),
.B1(n_819),
.B2(n_868),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_776),
.A2(n_801),
.B(n_888),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_848),
.B(n_840),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_764),
.B(n_792),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_851),
.A2(n_771),
.B(n_914),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_804),
.B(n_852),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_882),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_922),
.A2(n_807),
.B1(n_816),
.B2(n_815),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_923),
.A2(n_852),
.B1(n_867),
.B2(n_915),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_888),
.A2(n_771),
.B(n_916),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_793),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_795),
.A2(n_806),
.B1(n_852),
.B2(n_867),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_778),
.A2(n_813),
.B(n_850),
.C(n_871),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_846),
.A2(n_857),
.B(n_863),
.C(n_817),
.Y(n_1021)
);

AO32x1_ASAP7_75t_L g1022 ( 
.A1(n_920),
.A2(n_822),
.A3(n_901),
.B1(n_808),
.B2(n_873),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_912),
.A2(n_812),
.B(n_811),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_867),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_841),
.B(n_843),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_867),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_878),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_820),
.B(n_824),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_814),
.A2(n_785),
.B(n_907),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_919),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_894),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_849),
.B(n_908),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_879),
.A2(n_895),
.B1(n_906),
.B2(n_905),
.C(n_904),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_889),
.B(n_911),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_914),
.A2(n_919),
.B(n_907),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_903),
.A2(n_910),
.B(n_881),
.C(n_899),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_874),
.A2(n_891),
.B(n_845),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_SL g1038 ( 
.A(n_826),
.B(n_827),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_830),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_763),
.A2(n_619),
.B(n_595),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_810),
.B(n_628),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_SL g1042 ( 
.A(n_810),
.B(n_475),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_810),
.A2(n_760),
.B1(n_770),
.B2(n_652),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_810),
.A2(n_833),
.B(n_781),
.Y(n_1044)
);

AOI222xp33_ASAP7_75t_L g1045 ( 
.A1(n_818),
.A2(n_553),
.B1(n_421),
.B2(n_737),
.C1(n_736),
.C2(n_550),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_799),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_763),
.A2(n_619),
.B(n_595),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_810),
.A2(n_590),
.B(n_818),
.C(n_760),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_810),
.B(n_770),
.Y(n_1049)
);

AOI22x1_ASAP7_75t_L g1050 ( 
.A1(n_900),
.A2(n_833),
.B1(n_850),
.B2(n_876),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_786),
.B(n_858),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_SL g1052 ( 
.A1(n_760),
.A2(n_411),
.B(n_590),
.C(n_689),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_1043),
.A2(n_1020),
.A3(n_1021),
.B(n_931),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_1041),
.A2(n_952),
.B1(n_945),
.B2(n_999),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_948),
.B(n_1045),
.Y(n_1056)
);

AO31x2_ASAP7_75t_L g1057 ( 
.A1(n_983),
.A2(n_924),
.A3(n_1040),
.B(n_1047),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_949),
.A2(n_1049),
.B(n_1044),
.Y(n_1058)
);

AOI221x1_ASAP7_75t_L g1059 ( 
.A1(n_929),
.A2(n_924),
.B1(n_946),
.B2(n_998),
.C(n_961),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_948),
.A2(n_974),
.B1(n_1042),
.B2(n_959),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1049),
.A2(n_925),
.B(n_926),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_1037),
.A2(n_1012),
.B(n_954),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_978),
.B(n_930),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_SL g1064 ( 
.A1(n_927),
.A2(n_1048),
.B(n_960),
.C(n_971),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_937),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_937),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_974),
.A2(n_980),
.B1(n_960),
.B2(n_970),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_932),
.A2(n_934),
.B1(n_955),
.B2(n_971),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_926),
.A2(n_941),
.B(n_1023),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1017),
.A2(n_1005),
.B(n_1050),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_1036),
.A2(n_1029),
.B(n_1008),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_1007),
.A2(n_1002),
.A3(n_1010),
.B(n_936),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_975),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_1002),
.A2(n_1010),
.A3(n_1015),
.B(n_935),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_986),
.A2(n_987),
.B(n_973),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1052),
.A2(n_943),
.B(n_942),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_940),
.B(n_991),
.C(n_963),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_956),
.B(n_1051),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_956),
.B(n_1001),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_928),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1011),
.B(n_1018),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1025),
.A2(n_955),
.B(n_1032),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_984),
.A2(n_944),
.B(n_933),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_1024),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_947),
.B(n_995),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_953),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_964),
.B(n_965),
.C(n_966),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_988),
.Y(n_1088)
);

BUFx8_ASAP7_75t_L g1089 ( 
.A(n_939),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_967),
.A2(n_1032),
.B(n_1033),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_957),
.B(n_1046),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_1004),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1026),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_970),
.A2(n_977),
.B(n_973),
.C(n_938),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_993),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_999),
.A2(n_1014),
.B(n_1009),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_1031),
.A2(n_1039),
.A3(n_951),
.B(n_1019),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1030),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1027),
.A2(n_989),
.B(n_1000),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_993),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_969),
.B(n_972),
.C(n_962),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_1038),
.A2(n_977),
.B(n_1013),
.C(n_1035),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_958),
.A2(n_1013),
.B(n_950),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1003),
.B(n_981),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_997),
.B(n_950),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_997),
.A2(n_1016),
.B1(n_1006),
.B2(n_1028),
.Y(n_1106)
);

AO22x2_ASAP7_75t_L g1107 ( 
.A1(n_994),
.A2(n_1022),
.B1(n_1006),
.B2(n_996),
.Y(n_1107)
);

BUFx10_ASAP7_75t_L g1108 ( 
.A(n_1028),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_996),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_1022),
.A2(n_994),
.A3(n_1028),
.B(n_1034),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_994),
.Y(n_1111)
);

AOI221x1_ASAP7_75t_L g1112 ( 
.A1(n_1022),
.A2(n_992),
.B1(n_1034),
.B2(n_810),
.C(n_1043),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1043),
.A2(n_896),
.A3(n_834),
.B(n_1020),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1043),
.A2(n_896),
.A3(n_834),
.B(n_1020),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_978),
.B(n_858),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1048),
.A2(n_810),
.B(n_1043),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_984),
.A2(n_1044),
.B(n_1005),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1045),
.A2(n_810),
.B1(n_740),
.B2(n_1043),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_991),
.A2(n_613),
.B1(n_508),
.B2(n_553),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1048),
.A2(n_810),
.B(n_924),
.C(n_1041),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1041),
.B(n_453),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_952),
.A2(n_810),
.B(n_818),
.C(n_637),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_810),
.B1(n_1043),
.B2(n_952),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1051),
.B(n_803),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1045),
.A2(n_810),
.B1(n_740),
.B2(n_1043),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1048),
.A2(n_810),
.B(n_1043),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1043),
.A2(n_896),
.A3(n_834),
.B(n_1020),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1041),
.B(n_453),
.Y(n_1130)
);

INVx8_ASAP7_75t_L g1131 ( 
.A(n_1024),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1041),
.B(n_453),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_1043),
.A2(n_1049),
.B(n_1048),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_930),
.Y(n_1136)
);

INVx6_ASAP7_75t_SL g1137 ( 
.A(n_956),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_978),
.B(n_858),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_930),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1045),
.B(n_810),
.C(n_818),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_952),
.A2(n_810),
.B(n_818),
.C(n_637),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_974),
.A2(n_553),
.B1(n_737),
.B2(n_550),
.C(n_726),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1048),
.A2(n_810),
.B(n_924),
.C(n_1041),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1048),
.A2(n_810),
.B(n_924),
.C(n_1041),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1048),
.A2(n_810),
.B(n_1043),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1041),
.B(n_453),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_991),
.A2(n_613),
.B1(n_508),
.B2(n_553),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1043),
.A2(n_896),
.A3(n_834),
.B(n_1020),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1045),
.A2(n_810),
.B1(n_740),
.B2(n_1043),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1041),
.B(n_453),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_937),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_948),
.B(n_825),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_953),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_948),
.B(n_825),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_928),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1048),
.A2(n_810),
.B(n_1043),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_952),
.A2(n_810),
.B(n_818),
.C(n_637),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_993),
.B(n_1006),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_952),
.A2(n_810),
.B(n_818),
.C(n_637),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1041),
.B(n_453),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_1046),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1041),
.B(n_453),
.Y(n_1170)
);

BUFx2_ASAP7_75t_R g1171 ( 
.A(n_975),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_979),
.B(n_976),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1044),
.A2(n_955),
.B(n_1049),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_930),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_930),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_SL g1179 ( 
.A1(n_986),
.A2(n_1048),
.B(n_797),
.Y(n_1179)
);

BUFx4f_ASAP7_75t_L g1180 ( 
.A(n_978),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_SL g1181 ( 
.A1(n_986),
.A2(n_1048),
.B(n_797),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1043),
.A2(n_896),
.A3(n_834),
.B(n_1020),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_990),
.A2(n_985),
.B(n_968),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_L g1184 ( 
.A(n_1045),
.B(n_810),
.C(n_818),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_988),
.B(n_789),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1048),
.A2(n_810),
.B(n_1043),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1161),
.Y(n_1188)
);

INVx8_ASAP7_75t_L g1189 ( 
.A(n_1131),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1086),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1081),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1100),
.Y(n_1192)
);

INVx8_ASAP7_75t_L g1193 ( 
.A(n_1131),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1060),
.A2(n_1118),
.B1(n_1126),
.B2(n_1152),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1122),
.B(n_1130),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1060),
.A2(n_1126),
.B1(n_1118),
.B2(n_1152),
.Y(n_1196)
);

BUFx8_ASAP7_75t_SL g1197 ( 
.A(n_1157),
.Y(n_1197)
);

CKINVDCx6p67_ASAP7_75t_R g1198 ( 
.A(n_1168),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1119),
.A2(n_1149),
.B1(n_1087),
.B2(n_1186),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1125),
.B(n_1078),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1168),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1133),
.A2(n_1148),
.B1(n_1166),
.B2(n_1170),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1089),
.Y(n_1203)
);

BUFx4f_ASAP7_75t_SL g1204 ( 
.A(n_1137),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1085),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1116),
.A2(n_1147),
.B1(n_1162),
.B2(n_1127),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1089),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1067),
.A2(n_1124),
.B1(n_1154),
.B2(n_1134),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1055),
.A2(n_1158),
.B1(n_1156),
.B2(n_1075),
.Y(n_1209)
);

INVx6_ASAP7_75t_L g1210 ( 
.A(n_1084),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1095),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1084),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1084),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1078),
.Y(n_1214)
);

INVx8_ASAP7_75t_L g1215 ( 
.A(n_1185),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1059),
.A2(n_1180),
.B1(n_1112),
.B2(n_1098),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1173),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1179),
.A2(n_1181),
.B1(n_1117),
.B2(n_1058),
.Y(n_1218)
);

OAI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1077),
.A2(n_1146),
.B(n_1145),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1117),
.A2(n_1180),
.B1(n_1104),
.B2(n_1068),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1121),
.A2(n_1123),
.B1(n_1142),
.B2(n_1163),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1140),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1068),
.A2(n_1106),
.B1(n_1172),
.B2(n_1093),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1105),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1079),
.B(n_1115),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1165),
.A2(n_1139),
.B1(n_1063),
.B2(n_1137),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1076),
.A2(n_1083),
.B1(n_1099),
.B2(n_1065),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1101),
.A2(n_1155),
.B1(n_1066),
.B2(n_1136),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1090),
.A2(n_1096),
.B1(n_1082),
.B2(n_1178),
.Y(n_1229)
);

INVx6_ASAP7_75t_L g1230 ( 
.A(n_1185),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1090),
.A2(n_1175),
.B1(n_1091),
.B2(n_1061),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1171),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1073),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1164),
.B(n_1103),
.Y(n_1234)
);

INVx8_ASAP7_75t_L g1235 ( 
.A(n_1164),
.Y(n_1235)
);

INVx8_ASAP7_75t_L g1236 ( 
.A(n_1088),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1092),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1108),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1120),
.A2(n_1160),
.B1(n_1176),
.B2(n_1132),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1111),
.A2(n_1108),
.B1(n_1069),
.B2(n_1138),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1109),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1135),
.A2(n_1151),
.B(n_1153),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1109),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1064),
.A2(n_1107),
.B1(n_1070),
.B2(n_1111),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1107),
.A2(n_1094),
.B1(n_1072),
.B2(n_1074),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1072),
.A2(n_1054),
.B1(n_1074),
.B2(n_1129),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1071),
.A2(n_1072),
.B1(n_1128),
.B2(n_1183),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1053),
.A2(n_1174),
.B1(n_1143),
.B2(n_1159),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1057),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1074),
.A2(n_1054),
.B1(n_1102),
.B2(n_1097),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1062),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1054),
.A2(n_1177),
.B1(n_1169),
.B2(n_1167),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_L g1253 ( 
.A(n_1113),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1113),
.A2(n_1114),
.B1(n_1129),
.B2(n_1150),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1114),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1114),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1110),
.A2(n_1129),
.B1(n_1150),
.B2(n_1182),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1110),
.A2(n_1149),
.B1(n_1119),
.B2(n_1056),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1150),
.B(n_1110),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1141),
.A2(n_810),
.B1(n_1184),
.B2(n_1060),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1140),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1141),
.A2(n_810),
.B(n_1184),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1084),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1168),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1086),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1042),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1056),
.A2(n_1126),
.B1(n_1152),
.B2(n_1118),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1125),
.B(n_1078),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1141),
.A2(n_810),
.B1(n_1184),
.B2(n_1060),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1080),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1086),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1122),
.B(n_1130),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1131),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1141),
.A2(n_1184),
.B1(n_1056),
.B2(n_1144),
.Y(n_1279)
);

BUFx4_ASAP7_75t_SL g1280 ( 
.A(n_1086),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1084),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1056),
.A2(n_1126),
.B1(n_1152),
.B2(n_1118),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1086),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1084),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1131),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1080),
.Y(n_1286)
);

OAI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1144),
.A2(n_818),
.B(n_637),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1056),
.A2(n_1126),
.B1(n_1152),
.B2(n_1118),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1086),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1241),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1217),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1251),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1257),
.B(n_1254),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1253),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1239),
.A2(n_1248),
.B(n_1247),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1253),
.B(n_1206),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1256),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1249),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1256),
.B(n_1259),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1287),
.A2(n_1219),
.B(n_1196),
.C(n_1194),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1243),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1255),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1187),
.A2(n_1274),
.B1(n_1273),
.B2(n_1262),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1234),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1248),
.A2(n_1247),
.B(n_1250),
.Y(n_1306)
);

OAI211xp5_ASAP7_75t_L g1307 ( 
.A1(n_1199),
.A2(n_1187),
.B(n_1277),
.C(n_1273),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1260),
.A2(n_1271),
.B1(n_1263),
.B2(n_1221),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1244),
.B(n_1218),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1246),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1224),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1242),
.A2(n_1234),
.B(n_1240),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1218),
.B(n_1208),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1208),
.B(n_1240),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1229),
.A2(n_1231),
.B(n_1227),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1205),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1258),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1227),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1220),
.B(n_1229),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1188),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1238),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1272),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1262),
.A2(n_1267),
.B1(n_1279),
.B2(n_1277),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1220),
.B(n_1268),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1269),
.A2(n_1282),
.B(n_1288),
.C(n_1202),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1231),
.A2(n_1228),
.B(n_1209),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1228),
.A2(n_1209),
.B(n_1199),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1216),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1216),
.B(n_1282),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1269),
.A2(n_1288),
.B(n_1202),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1286),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1197),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1223),
.B(n_1252),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1215),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1267),
.B(n_1279),
.Y(n_1335)
);

BUFx2_ASAP7_75t_SL g1336 ( 
.A(n_1201),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1274),
.B(n_1191),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1195),
.B(n_1276),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1200),
.B(n_1270),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1226),
.B(n_1214),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1222),
.A2(n_1261),
.A3(n_1278),
.B(n_1211),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1225),
.A2(n_1213),
.B(n_1237),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1235),
.Y(n_1343)
);

CKINVDCx9p33_ASAP7_75t_R g1344 ( 
.A(n_1280),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1235),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1341),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1323),
.A2(n_1230),
.B1(n_1198),
.B2(n_1203),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1295),
.A2(n_1215),
.B(n_1230),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1325),
.A2(n_1284),
.B(n_1281),
.C(n_1189),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1300),
.A2(n_1207),
.B(n_1230),
.C(n_1212),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1290),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1290),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1301),
.B(n_1316),
.Y(n_1353)
);

OAI211xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1323),
.A2(n_1289),
.B(n_1283),
.C(n_1275),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1303),
.A2(n_1233),
.B1(n_1265),
.B2(n_1232),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1303),
.B(n_1284),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1316),
.B(n_1285),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1308),
.B(n_1192),
.C(n_1190),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1308),
.A2(n_1192),
.B(n_1266),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1300),
.A2(n_1192),
.B(n_1278),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1338),
.B(n_1311),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1307),
.B(n_1210),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1293),
.B(n_1210),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1294),
.B(n_1192),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1344),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1320),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1296),
.B(n_1264),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1296),
.B(n_1339),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1307),
.A2(n_1203),
.B1(n_1236),
.B2(n_1189),
.C(n_1193),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_SL g1370 ( 
.A1(n_1325),
.A2(n_1189),
.B(n_1193),
.C(n_1204),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1335),
.B(n_1210),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1327),
.A2(n_1236),
.B(n_1204),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1335),
.B(n_1193),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1296),
.B(n_1236),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1306),
.A2(n_1315),
.B(n_1295),
.Y(n_1375)
);

INVx3_ASAP7_75t_SL g1376 ( 
.A(n_1332),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1317),
.A2(n_1329),
.B1(n_1328),
.B2(n_1318),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1306),
.A2(n_1295),
.B(n_1315),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1306),
.A2(n_1315),
.B(n_1312),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1290),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1293),
.B(n_1299),
.Y(n_1381)
);

NOR3xp33_ASAP7_75t_SL g1382 ( 
.A(n_1340),
.B(n_1345),
.C(n_1343),
.Y(n_1382)
);

NOR2x1_ASAP7_75t_L g1383 ( 
.A(n_1334),
.B(n_1298),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1299),
.B(n_1319),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1317),
.A2(n_1330),
.B1(n_1324),
.B2(n_1318),
.Y(n_1385)
);

AO32x2_ASAP7_75t_L g1386 ( 
.A1(n_1304),
.A2(n_1292),
.A3(n_1321),
.B1(n_1328),
.B2(n_1291),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1339),
.B(n_1342),
.Y(n_1387)
);

AO32x2_ASAP7_75t_L g1388 ( 
.A1(n_1304),
.A2(n_1292),
.A3(n_1321),
.B1(n_1328),
.B2(n_1291),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1317),
.A2(n_1330),
.B1(n_1324),
.B2(n_1340),
.Y(n_1389)
);

NOR2x1_ASAP7_75t_SL g1390 ( 
.A(n_1330),
.B(n_1294),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1294),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1312),
.A2(n_1326),
.B(n_1327),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1319),
.B(n_1310),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1391),
.B(n_1304),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1389),
.A2(n_1329),
.B1(n_1324),
.B2(n_1302),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1384),
.B(n_1305),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1387),
.B(n_1310),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1355),
.B(n_1336),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1386),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1351),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1358),
.A2(n_1330),
.B1(n_1329),
.B2(n_1356),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1365),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1386),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1351),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1361),
.B(n_1305),
.Y(n_1405)
);

OAI211xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1385),
.A2(n_1321),
.B(n_1322),
.C(n_1331),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1352),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1357),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1362),
.A2(n_1330),
.B1(n_1356),
.B2(n_1314),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1377),
.A2(n_1314),
.B1(n_1327),
.B2(n_1302),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1353),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1380),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1392),
.B(n_1312),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1366),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1381),
.B(n_1319),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1386),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1386),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1381),
.B(n_1309),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1388),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1393),
.B(n_1309),
.Y(n_1420)
);

NOR2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1364),
.B(n_1302),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1388),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1392),
.B(n_1297),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1364),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1392),
.B(n_1379),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1407),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1397),
.B(n_1393),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1412),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1411),
.B(n_1368),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1399),
.B(n_1378),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1425),
.A2(n_1378),
.B(n_1390),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1399),
.B(n_1388),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1409),
.A2(n_1302),
.B1(n_1359),
.B2(n_1314),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1395),
.A2(n_1354),
.B1(n_1313),
.B2(n_1337),
.Y(n_1434)
);

OAI321xp33_ASAP7_75t_L g1435 ( 
.A1(n_1409),
.A2(n_1360),
.A3(n_1372),
.B1(n_1362),
.B2(n_1347),
.C(n_1337),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1395),
.A2(n_1401),
.B1(n_1410),
.B2(n_1333),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1403),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1403),
.B(n_1388),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1423),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1394),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1410),
.A2(n_1313),
.B1(n_1326),
.B2(n_1333),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1416),
.B(n_1346),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1425),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1400),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1411),
.B(n_1367),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1400),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1424),
.Y(n_1447)
);

NAND5xp2_ASAP7_75t_L g1448 ( 
.A(n_1398),
.B(n_1369),
.C(n_1350),
.D(n_1370),
.E(n_1373),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1404),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1413),
.A2(n_1348),
.B(n_1379),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1394),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1408),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1415),
.B(n_1375),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1443),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1430),
.B(n_1396),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1447),
.B(n_1421),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1444),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1444),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1452),
.B(n_1414),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1444),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1440),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1440),
.B(n_1418),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1452),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1446),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1447),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1440),
.B(n_1418),
.Y(n_1466)
);

NOR3xp33_ASAP7_75t_SL g1467 ( 
.A(n_1448),
.B(n_1406),
.C(n_1349),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1446),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1430),
.B(n_1396),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1447),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1445),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1445),
.B(n_1376),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1440),
.B(n_1451),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1446),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1429),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1449),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1449),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1447),
.B(n_1421),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1426),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1451),
.B(n_1408),
.Y(n_1480)
);

AND2x2_ASAP7_75t_SL g1481 ( 
.A(n_1441),
.B(n_1342),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1447),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1428),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1430),
.B(n_1405),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1451),
.B(n_1437),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1442),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1451),
.B(n_1424),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1443),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1484),
.B(n_1437),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1457),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1457),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1456),
.B(n_1453),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1488),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1488),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1486),
.B(n_1432),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1486),
.B(n_1432),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1458),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1475),
.B(n_1432),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1463),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1458),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1471),
.B(n_1429),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1456),
.B(n_1439),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1438),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1467),
.A2(n_1436),
.B1(n_1441),
.B2(n_1434),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1454),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1460),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1460),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1488),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1454),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1459),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1484),
.B(n_1442),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1456),
.Y(n_1513)
);

NAND2x1_ASAP7_75t_L g1514 ( 
.A(n_1478),
.B(n_1438),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1464),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1454),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1485),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1464),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1459),
.B(n_1438),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1478),
.B(n_1453),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1453),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1468),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1468),
.Y(n_1523)
);

NOR2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1478),
.B(n_1334),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1485),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1480),
.B(n_1420),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1473),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1420),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1465),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1499),
.B(n_1455),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1505),
.B(n_1462),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1491),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1491),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1524),
.B(n_1465),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1492),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1499),
.B(n_1455),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1530),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1505),
.B(n_1462),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1514),
.A2(n_1436),
.B1(n_1433),
.B2(n_1435),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1530),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1500),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1502),
.B(n_1376),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1492),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1524),
.B(n_1470),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1498),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1433),
.C(n_1434),
.Y(n_1549)
);

INVxp33_ASAP7_75t_SL g1550 ( 
.A(n_1525),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1504),
.B(n_1427),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1514),
.B(n_1383),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1504),
.B(n_1427),
.Y(n_1553)
);

NAND2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1517),
.B(n_1365),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1498),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1529),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1490),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1494),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1513),
.B(n_1470),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1494),
.A2(n_1482),
.B(n_1479),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1466),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1501),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1513),
.B(n_1482),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1513),
.B(n_1473),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1466),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1533),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1544),
.B(n_1472),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1554),
.B(n_1481),
.Y(n_1568)
);

OAI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1554),
.A2(n_1517),
.B1(n_1513),
.B2(n_1497),
.C(n_1496),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1541),
.B(n_1481),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1534),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1536),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1549),
.A2(n_1481),
.B(n_1435),
.C(n_1496),
.Y(n_1573)
);

AOI321xp33_ASAP7_75t_L g1574 ( 
.A1(n_1532),
.A2(n_1490),
.A3(n_1521),
.B1(n_1520),
.B2(n_1493),
.C(n_1503),
.Y(n_1574)
);

OAI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1540),
.A2(n_1497),
.B1(n_1489),
.B2(n_1461),
.C(n_1512),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1550),
.Y(n_1576)
);

AOI322xp5_ASAP7_75t_L g1577 ( 
.A1(n_1557),
.A2(n_1422),
.A3(n_1419),
.B1(n_1417),
.B2(n_1416),
.C1(n_1520),
.C2(n_1493),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1538),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1550),
.B(n_1521),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1547),
.A2(n_1489),
.B(n_1382),
.C(n_1406),
.Y(n_1580)
);

NAND2x1_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1503),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1538),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1542),
.A2(n_1448),
.B1(n_1333),
.B2(n_1431),
.Y(n_1583)
);

NAND4xp25_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1373),
.C(n_1350),
.D(n_1371),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1547),
.A2(n_1503),
.B1(n_1487),
.B2(n_1461),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1535),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1561),
.B(n_1349),
.C(n_1371),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1556),
.A2(n_1431),
.B1(n_1309),
.B2(n_1313),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1535),
.A2(n_1503),
.B(n_1487),
.C(n_1450),
.Y(n_1589)
);

AND3x1_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1374),
.C(n_1363),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1586),
.B(n_1564),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1566),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1571),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1578),
.B(n_1565),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1572),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1576),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1570),
.A2(n_1552),
.B(n_1559),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1582),
.B(n_1559),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1583),
.A2(n_1568),
.B1(n_1569),
.B2(n_1573),
.Y(n_1599)
);

OAI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1583),
.A2(n_1537),
.B(n_1531),
.Y(n_1600)
);

NOR2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1579),
.B(n_1551),
.Y(n_1601)
);

AOI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1575),
.A2(n_1563),
.B(n_1562),
.C(n_1548),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1588),
.A2(n_1545),
.B1(n_1555),
.B2(n_1563),
.C(n_1537),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1587),
.B(n_1551),
.Y(n_1604)
);

AOI221x1_ASAP7_75t_L g1605 ( 
.A1(n_1580),
.A2(n_1558),
.B1(n_1507),
.B2(n_1518),
.C(n_1501),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1581),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1585),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1574),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1567),
.B(n_1552),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1588),
.B(n_1402),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1591),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1608),
.B(n_1577),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1605),
.A2(n_1589),
.B(n_1558),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1606),
.B(n_1590),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1610),
.A2(n_1584),
.B(n_1560),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1607),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1607),
.B(n_1553),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1599),
.A2(n_1495),
.B(n_1494),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1598),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1610),
.A2(n_1560),
.B(n_1531),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1616),
.B(n_1596),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1617),
.Y(n_1622)
);

NOR3xp33_ASAP7_75t_L g1623 ( 
.A(n_1619),
.B(n_1594),
.C(n_1603),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1617),
.B(n_1601),
.Y(n_1624)
);

AOI21xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1613),
.A2(n_1609),
.B(n_1604),
.Y(n_1625)
);

AOI211x1_ASAP7_75t_L g1626 ( 
.A1(n_1620),
.A2(n_1597),
.B(n_1609),
.C(n_1600),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1614),
.B(n_1619),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1613),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1625),
.A2(n_1612),
.B1(n_1615),
.B2(n_1602),
.C(n_1611),
.Y(n_1630)
);

AOI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1628),
.A2(n_1611),
.B(n_1593),
.C(n_1595),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_SL g1632 ( 
.A(n_1623),
.B(n_1624),
.C(n_1622),
.Y(n_1632)
);

AOI21xp33_ASAP7_75t_L g1633 ( 
.A1(n_1629),
.A2(n_1618),
.B(n_1614),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1621),
.A2(n_1618),
.B(n_1560),
.Y(n_1634)
);

AND4x2_ASAP7_75t_L g1635 ( 
.A(n_1630),
.B(n_1626),
.C(n_1618),
.D(n_1627),
.Y(n_1635)
);

OAI321xp33_ASAP7_75t_L g1636 ( 
.A1(n_1632),
.A2(n_1631),
.A3(n_1634),
.B1(n_1633),
.B2(n_1546),
.C(n_1539),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1630),
.A2(n_1553),
.B1(n_1546),
.B2(n_1539),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1631),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1633),
.A2(n_1370),
.B(n_1344),
.C(n_1512),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1634),
.B(n_1487),
.Y(n_1640)
);

AO22x2_ASAP7_75t_L g1641 ( 
.A1(n_1638),
.A2(n_1336),
.B1(n_1523),
.B2(n_1522),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1637),
.B(n_1507),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1636),
.A2(n_1506),
.B(n_1495),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_L g1644 ( 
.A(n_1639),
.B(n_1506),
.C(n_1495),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1640),
.A2(n_1527),
.B1(n_1523),
.B2(n_1522),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1644),
.A2(n_1635),
.B1(n_1527),
.B2(n_1518),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1641),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1642),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1647),
.B(n_1643),
.C(n_1645),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1649),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1650),
.A2(n_1648),
.B1(n_1646),
.B2(n_1516),
.Y(n_1651)
);

OAI22x1_ASAP7_75t_SL g1652 ( 
.A1(n_1651),
.A2(n_1515),
.B1(n_1508),
.B2(n_1510),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1652),
.A2(n_1509),
.B(n_1506),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1653),
.A2(n_1510),
.B(n_1509),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1653),
.A2(n_1516),
.B1(n_1510),
.B2(n_1509),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1654),
.B(n_1516),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1655),
.B(n_1508),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1656),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1657),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1515),
.B1(n_1477),
.B2(n_1476),
.C(n_1474),
.Y(n_1660)
);

AOI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1660),
.A2(n_1659),
.B(n_1334),
.C(n_1364),
.Y(n_1661)
);


endmodule