module fake_netlist_1_3955_n_32 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_11), .Y(n_15) );
OAI22xp5_ASAP7_75t_SL g16 ( .A1(n_5), .A2(n_12), .B1(n_4), .B2(n_8), .Y(n_16) );
OAI22xp5_ASAP7_75t_SL g17 ( .A1(n_7), .A2(n_10), .B1(n_2), .B2(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
INVx5_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_14), .B(n_0), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_21), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_18), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_15), .Y(n_24) );
NAND4xp25_ASAP7_75t_L g25 ( .A(n_24), .B(n_23), .C(n_19), .D(n_16), .Y(n_25) );
AO21x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_24), .B(n_17), .Y(n_26) );
XNOR2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_15), .Y(n_27) );
NAND2xp5_ASAP7_75t_SL g28 ( .A(n_27), .B(n_14), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AOI222xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_26), .B1(n_20), .B2(n_4), .C1(n_5), .C2(n_1), .Y(n_30) );
OAI22x1_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_29), .B1(n_20), .B2(n_6), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_3), .B1(n_9), .B2(n_13), .Y(n_32) );
endmodule