module real_aes_11318_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_1404;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_0), .A2(n_81), .B1(n_704), .B2(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1082 ( .A(n_0), .Y(n_1082) );
INVxp33_ASAP7_75t_L g395 ( .A(n_1), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_1), .A2(n_498), .B(n_501), .Y(n_497) );
INVxp67_ASAP7_75t_SL g1255 ( .A(n_2), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_2), .A2(n_10), .B1(n_612), .B2(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1488 ( .A(n_3), .Y(n_1488) );
INVx1_ASAP7_75t_L g571 ( .A(n_4), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g1105 ( .A1(n_5), .A2(n_16), .B1(n_536), .B2(n_1106), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g1128 ( .A(n_5), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_6), .A2(n_165), .B1(n_1184), .B2(n_1226), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_6), .A2(n_165), .B1(n_1235), .B2(n_1239), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_7), .A2(n_228), .B1(n_682), .B2(n_1061), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_7), .A2(n_228), .B1(n_1226), .B2(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1249 ( .A(n_8), .Y(n_1249) );
INVx1_ASAP7_75t_L g1053 ( .A(n_9), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_9), .A2(n_255), .B1(n_612), .B2(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1254 ( .A(n_10), .Y(n_1254) );
INVxp67_ASAP7_75t_SL g922 ( .A(n_11), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_11), .A2(n_58), .B1(n_553), .B2(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g1579 ( .A(n_12), .Y(n_1579) );
INVxp33_ASAP7_75t_SL g1100 ( .A(n_13), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_13), .A2(n_318), .B1(n_1030), .B2(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g864 ( .A(n_14), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_14), .A2(n_207), .B1(n_534), .B2(n_776), .Y(n_881) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_15), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_15), .A2(n_216), .B1(n_591), .B2(n_960), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1129 ( .A(n_16), .Y(n_1129) );
INVx1_ASAP7_75t_L g1248 ( .A(n_17), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_17), .A2(n_55), .B1(n_614), .B2(n_1231), .Y(n_1273) );
AO221x2_ASAP7_75t_L g1577 ( .A1(n_18), .A2(n_267), .B1(n_1534), .B2(n_1555), .C(n_1578), .Y(n_1577) );
INVxp33_ASAP7_75t_L g963 ( .A(n_19), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_19), .A2(n_34), .B1(n_635), .B2(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1343 ( .A(n_20), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_20), .A2(n_323), .B1(n_1015), .B2(n_1194), .Y(n_1357) );
CKINVDCx16_ASAP7_75t_R g1586 ( .A(n_21), .Y(n_1586) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_22), .A2(n_353), .B1(n_661), .B2(n_1070), .Y(n_1073) );
INVx1_ASAP7_75t_L g1079 ( .A(n_22), .Y(n_1079) );
XOR2x2_ASAP7_75t_L g1087 ( .A(n_23), .B(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1384 ( .A(n_24), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_25), .A2(n_69), .B1(n_677), .B2(n_1162), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_25), .A2(n_69), .B1(n_1174), .B2(n_1177), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_26), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_26), .A2(n_212), .B1(n_534), .B2(n_536), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g1767 ( .A1(n_27), .A2(n_549), .B(n_579), .C(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1783 ( .A(n_27), .Y(n_1783) );
OAI222xp33_ASAP7_75t_L g847 ( .A1(n_28), .A2(n_74), .B1(n_223), .B2(n_848), .C1(n_851), .C2(n_854), .Y(n_847) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_28), .A2(n_186), .B1(n_753), .B2(n_754), .Y(n_887) );
INVx1_ASAP7_75t_L g1145 ( .A(n_29), .Y(n_1145) );
INVx1_ASAP7_75t_L g1304 ( .A(n_30), .Y(n_1304) );
AOI22xp33_ASAP7_75t_SL g1318 ( .A1(n_30), .A2(n_197), .B1(n_1184), .B2(n_1185), .Y(n_1318) );
CKINVDCx5p33_ASAP7_75t_R g1428 ( .A(n_31), .Y(n_1428) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_32), .A2(n_85), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_32), .A2(n_85), .B1(n_534), .B2(n_553), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g1788 ( .A(n_33), .Y(n_1788) );
INVx1_ASAP7_75t_L g957 ( .A(n_34), .Y(n_957) );
INVx1_ASAP7_75t_L g1378 ( .A(n_35), .Y(n_1378) );
INVx1_ASAP7_75t_L g860 ( .A(n_36), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_36), .A2(n_179), .B1(n_749), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_37), .A2(n_78), .B1(n_488), .B2(n_612), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_37), .A2(n_78), .B1(n_830), .B2(n_938), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_38), .A2(n_111), .B1(n_452), .B2(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_38), .A2(n_111), .B1(n_534), .B2(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g366 ( .A(n_39), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g1204 ( .A1(n_40), .A2(n_233), .B1(n_685), .B2(n_749), .C(n_1205), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_40), .A2(n_233), .B1(n_1184), .B2(n_1185), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_41), .A2(n_224), .B1(n_750), .B2(n_757), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_41), .A2(n_224), .B1(n_534), .B2(n_938), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_42), .A2(n_114), .B1(n_1015), .B2(n_1017), .Y(n_1014) );
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_42), .A2(n_114), .B1(n_672), .B2(n_1030), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_43), .A2(n_343), .B1(n_757), .B2(n_889), .Y(n_1028) );
AOI22xp33_ASAP7_75t_SL g1038 ( .A1(n_43), .A2(n_234), .B1(n_695), .B2(n_1039), .Y(n_1038) );
INVxp33_ASAP7_75t_L g745 ( .A(n_44), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_44), .A2(n_291), .B1(n_768), .B2(n_773), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g1429 ( .A(n_45), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_46), .A2(n_192), .B1(n_1231), .B2(n_1309), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_46), .A2(n_192), .B1(n_661), .B2(n_1070), .Y(n_1314) );
INVxp33_ASAP7_75t_SL g572 ( .A(n_47), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_47), .A2(n_195), .B1(n_488), .B2(n_612), .Y(n_611) );
INVxp33_ASAP7_75t_SL g603 ( .A(n_48), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_48), .A2(n_66), .B1(n_633), .B2(n_635), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g1591 ( .A1(n_49), .A2(n_324), .B1(n_1534), .B2(n_1555), .Y(n_1591) );
INVxp67_ASAP7_75t_SL g1141 ( .A(n_50), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_50), .A2(n_64), .B1(n_1182), .B2(n_1185), .Y(n_1181) );
INVxp33_ASAP7_75t_SL g1024 ( .A(n_51), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_51), .A2(n_160), .B1(n_695), .B2(n_1042), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_52), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_52), .A2(n_211), .B1(n_684), .B2(n_685), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_53), .A2(n_105), .B1(n_1235), .B2(n_1239), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_53), .A2(n_97), .B1(n_1473), .B2(n_1474), .Y(n_1472) );
INVx1_ASAP7_75t_L g1223 ( .A(n_54), .Y(n_1223) );
INVx1_ASAP7_75t_L g1251 ( .A(n_55), .Y(n_1251) );
INVx1_ASAP7_75t_L g1258 ( .A(n_56), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_56), .A2(n_249), .B1(n_732), .B2(n_773), .Y(n_1280) );
OAI211xp5_ASAP7_75t_L g1195 ( .A1(n_57), .A2(n_579), .B(n_1196), .C(n_1198), .Y(n_1195) );
INVx1_ASAP7_75t_L g1215 ( .A(n_57), .Y(n_1215) );
INVxp33_ASAP7_75t_SL g923 ( .A(n_58), .Y(n_923) );
AO22x2_ASAP7_75t_L g898 ( .A1(n_59), .A2(n_899), .B1(n_947), .B2(n_948), .Y(n_898) );
CKINVDCx14_ASAP7_75t_R g947 ( .A(n_59), .Y(n_947) );
XNOR2xp5_ASAP7_75t_L g1044 ( .A(n_60), .B(n_1045), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_61), .Y(n_859) );
INVx1_ASAP7_75t_L g1491 ( .A(n_62), .Y(n_1491) );
INVx1_ASAP7_75t_L g1486 ( .A(n_63), .Y(n_1486) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_63), .A2(n_156), .B1(n_536), .B2(n_1157), .Y(n_1508) );
INVxp67_ASAP7_75t_SL g1148 ( .A(n_64), .Y(n_1148) );
INVx1_ASAP7_75t_L g908 ( .A(n_65), .Y(n_908) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_66), .Y(n_584) );
INVx1_ASAP7_75t_L g796 ( .A(n_67), .Y(n_796) );
INVx1_ASAP7_75t_L g1376 ( .A(n_68), .Y(n_1376) );
AO22x2_ASAP7_75t_L g1421 ( .A1(n_70), .A2(n_1422), .B1(n_1423), .B2(n_1476), .Y(n_1421) );
INVxp67_ASAP7_75t_L g1476 ( .A(n_70), .Y(n_1476) );
CKINVDCx5p33_ASAP7_75t_R g1361 ( .A(n_71), .Y(n_1361) );
INVxp33_ASAP7_75t_SL g1498 ( .A(n_72), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_72), .A2(n_146), .B1(n_677), .B2(n_1453), .Y(n_1514) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_73), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_73), .A2(n_302), .B1(n_934), .B2(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g869 ( .A(n_74), .Y(n_869) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_75), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_75), .A2(n_271), .B1(n_534), .B2(n_553), .Y(n_552) );
XOR2xp5_ASAP7_75t_L g999 ( .A(n_76), .B(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1009 ( .A(n_77), .Y(n_1009) );
OAI222xp33_ASAP7_75t_L g1021 ( .A1(n_77), .A2(n_174), .B1(n_269), .B2(n_493), .C1(n_711), .C2(n_740), .Y(n_1021) );
AOI221xp5_ASAP7_75t_L g1784 ( .A1(n_79), .A2(n_256), .B1(n_934), .B2(n_1785), .C(n_1786), .Y(n_1784) );
AOI22xp33_ASAP7_75t_L g1791 ( .A1(n_79), .A2(n_256), .B1(n_1176), .B2(n_1185), .Y(n_1791) );
OAI21xp33_ASAP7_75t_SL g1004 ( .A1(n_80), .A2(n_1005), .B(n_1008), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_80), .A2(n_306), .B1(n_488), .B2(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1083 ( .A(n_81), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_82), .A2(n_90), .B1(n_625), .B2(n_628), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_82), .A2(n_90), .B1(n_633), .B2(n_635), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_83), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1778 ( .A1(n_84), .A2(n_240), .B1(n_1235), .B2(n_1239), .Y(n_1778) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_84), .A2(n_240), .B1(n_1176), .B2(n_1226), .Y(n_1794) );
BUFx2_ASAP7_75t_L g445 ( .A(n_86), .Y(n_445) );
BUFx2_ASAP7_75t_L g558 ( .A(n_86), .Y(n_558) );
INVx1_ASAP7_75t_L g619 ( .A(n_86), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_87), .A2(n_246), .B1(n_575), .B2(n_765), .Y(n_1104) );
INVxp67_ASAP7_75t_SL g1123 ( .A(n_87), .Y(n_1123) );
INVx1_ASAP7_75t_L g574 ( .A(n_88), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_88), .A2(n_109), .B1(n_583), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_89), .A2(n_347), .B1(n_534), .B2(n_1110), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_89), .A2(n_347), .B1(n_1030), .B2(n_1118), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_91), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_91), .A2(n_305), .B1(n_591), .B2(n_740), .Y(n_920) );
AO22x2_ASAP7_75t_L g842 ( .A1(n_92), .A2(n_843), .B1(n_844), .B2(n_895), .Y(n_842) );
INVx1_ASAP7_75t_L g895 ( .A(n_92), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_93), .A2(n_284), .B1(n_575), .B2(n_836), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_93), .A2(n_284), .B1(n_737), .B2(n_823), .Y(n_1120) );
INVx1_ASAP7_75t_L g1290 ( .A(n_94), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_94), .A2(n_351), .B1(n_679), .B2(n_682), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_95), .A2(n_279), .B1(n_612), .B2(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_95), .A2(n_279), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_96), .A2(n_311), .B1(n_583), .B2(n_671), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_96), .A2(n_311), .B1(n_700), .B2(n_794), .Y(n_1172) );
INVx1_ASAP7_75t_L g1432 ( .A(n_97), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g1776 ( .A(n_98), .Y(n_1776) );
OAI22xp33_ASAP7_75t_L g1201 ( .A1(n_99), .A2(n_245), .B1(n_1017), .B2(n_1202), .Y(n_1201) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_99), .A2(n_245), .B1(n_677), .B2(n_1167), .C(n_1211), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_100), .A2(n_234), .B1(n_823), .B2(n_1027), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_100), .A2(n_343), .B1(n_1035), .B2(n_1037), .Y(n_1034) );
INVx1_ASAP7_75t_L g1411 ( .A(n_101), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_102), .A2(n_112), .B1(n_854), .B2(n_1295), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_102), .A2(n_112), .B1(n_591), .B2(n_960), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_103), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_103), .A2(n_232), .B1(n_749), .B2(n_820), .Y(n_819) );
CKINVDCx16_ASAP7_75t_R g1588 ( .A(n_104), .Y(n_1588) );
INVx1_ASAP7_75t_L g1471 ( .A(n_105), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_106), .A2(n_132), .B1(n_1506), .B2(n_1507), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_106), .A2(n_132), .B1(n_867), .B2(n_1453), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_107), .A2(n_260), .B1(n_768), .B2(n_877), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_107), .A2(n_260), .B1(n_762), .B2(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g1206 ( .A(n_108), .Y(n_1206) );
INVxp33_ASAP7_75t_SL g567 ( .A(n_109), .Y(n_567) );
INVx1_ASAP7_75t_L g1405 ( .A(n_110), .Y(n_1405) );
INVxp33_ASAP7_75t_SL g1483 ( .A(n_113), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_113), .A2(n_158), .B1(n_1504), .B2(n_1510), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g1787 ( .A(n_115), .Y(n_1787) );
INVx1_ASAP7_75t_L g1388 ( .A(n_116), .Y(n_1388) );
OAI22xp33_ASAP7_75t_SL g1417 ( .A1(n_116), .A2(n_214), .B1(n_375), .B2(n_1235), .Y(n_1417) );
INVx1_ASAP7_75t_L g1200 ( .A(n_117), .Y(n_1200) );
AOI22xp5_ASAP7_75t_L g1576 ( .A1(n_118), .A2(n_320), .B1(n_1534), .B2(n_1555), .Y(n_1576) );
INVxp33_ASAP7_75t_SL g742 ( .A(n_119), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_119), .A2(n_213), .B1(n_775), .B2(n_776), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_120), .A2(n_252), .B1(n_575), .B2(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_120), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_121), .A2(n_202), .B1(n_694), .B2(n_776), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_121), .A2(n_202), .B1(n_757), .B2(n_889), .Y(n_888) );
XOR2xp5_ASAP7_75t_L g1320 ( .A(n_122), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g964 ( .A(n_123), .Y(n_964) );
INVx1_ASAP7_75t_L g1052 ( .A(n_124), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_124), .A2(n_257), .B1(n_583), .B2(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g662 ( .A(n_125), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_125), .A2(n_303), .B1(n_589), .B2(n_711), .Y(n_710) );
INVxp33_ASAP7_75t_L g1151 ( .A(n_126), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_126), .A2(n_183), .B1(n_671), .B2(n_1170), .Y(n_1169) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_127), .A2(n_299), .B1(n_753), .B2(n_754), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_127), .A2(n_299), .B1(n_765), .B2(n_768), .Y(n_764) );
INVxp33_ASAP7_75t_SL g726 ( .A(n_128), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_128), .A2(n_341), .B1(n_757), .B2(n_759), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g1565 ( .A1(n_129), .A2(n_131), .B1(n_1566), .B2(n_1569), .Y(n_1565) );
INVx1_ASAP7_75t_L g1401 ( .A(n_130), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g1407 ( .A1(n_130), .A2(n_138), .B1(n_1015), .B2(n_1017), .Y(n_1407) );
INVx1_ASAP7_75t_L g1140 ( .A(n_133), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1571 ( .A1(n_134), .A2(n_339), .B1(n_1526), .B2(n_1572), .Y(n_1571) );
INVxp33_ASAP7_75t_L g972 ( .A(n_135), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_135), .A2(n_321), .B1(n_583), .B2(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g1341 ( .A(n_136), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_136), .A2(n_292), .B1(n_1017), .B2(n_1202), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_137), .A2(n_180), .B1(n_375), .B2(n_606), .Y(n_1020) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_137), .A2(n_269), .B1(n_698), .B2(n_1037), .Y(n_1040) );
INVx1_ASAP7_75t_L g1404 ( .A(n_138), .Y(n_1404) );
AO221x2_ASAP7_75t_L g1599 ( .A1(n_139), .A2(n_205), .B1(n_1526), .B2(n_1534), .C(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1531 ( .A(n_140), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_141), .Y(n_1532) );
INVxp33_ASAP7_75t_SL g785 ( .A(n_142), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_142), .A2(n_296), .B1(n_817), .B2(n_823), .Y(n_822) );
INVxp33_ASAP7_75t_SL g653 ( .A(n_143), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_143), .A2(n_188), .B1(n_671), .B2(n_687), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_144), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_145), .A2(n_239), .B1(n_614), .B2(n_918), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_145), .A2(n_239), .B1(n_903), .B2(n_1276), .Y(n_1275) );
INVxp67_ASAP7_75t_SL g1500 ( .A(n_146), .Y(n_1500) );
XNOR2xp5_ASAP7_75t_L g391 ( .A(n_147), .B(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g1590 ( .A1(n_147), .A2(n_350), .B1(n_1566), .B2(n_1569), .Y(n_1590) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_148), .Y(n_1143) );
INVx1_ASAP7_75t_L g733 ( .A(n_149), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_149), .A2(n_286), .B1(n_711), .B2(n_740), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g1436 ( .A1(n_150), .A2(n_579), .B(n_1437), .C(n_1439), .Y(n_1436) );
INVx1_ASAP7_75t_L g1459 ( .A(n_150), .Y(n_1459) );
AO22x2_ASAP7_75t_SL g648 ( .A1(n_151), .A2(n_649), .B1(n_650), .B2(n_718), .Y(n_648) );
CKINVDCx16_ASAP7_75t_R g649 ( .A(n_151), .Y(n_649) );
INVx1_ASAP7_75t_L g1353 ( .A(n_152), .Y(n_1353) );
OAI22xp33_ASAP7_75t_SL g1370 ( .A1(n_152), .A2(n_164), .B1(n_375), .B2(n_1235), .Y(n_1370) );
INVxp33_ASAP7_75t_SL g1091 ( .A(n_153), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_153), .A2(n_162), .B1(n_672), .B2(n_737), .Y(n_1115) );
INVx1_ASAP7_75t_L g1529 ( .A(n_154), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_154), .B(n_1542), .Y(n_1547) );
INVxp33_ASAP7_75t_SL g915 ( .A(n_155), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_155), .A2(n_327), .B1(n_765), .B2(n_942), .Y(n_941) );
INVxp67_ASAP7_75t_SL g1484 ( .A(n_156), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_157), .A2(n_222), .B1(n_675), .B2(n_980), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_157), .A2(n_222), .B1(n_661), .B2(n_1070), .Y(n_1069) );
INVxp33_ASAP7_75t_SL g1490 ( .A(n_158), .Y(n_1490) );
OAI22xp5_ASAP7_75t_L g1765 ( .A1(n_159), .A2(n_173), .B1(n_1015), .B2(n_1017), .Y(n_1765) );
AOI221xp5_ASAP7_75t_L g1780 ( .A1(n_159), .A2(n_307), .B1(n_677), .B2(n_680), .C(n_1781), .Y(n_1780) );
INVxp33_ASAP7_75t_L g1023 ( .A(n_160), .Y(n_1023) );
INVx2_ASAP7_75t_L g378 ( .A(n_161), .Y(n_378) );
INVxp67_ASAP7_75t_SL g1094 ( .A(n_162), .Y(n_1094) );
INVxp33_ASAP7_75t_L g725 ( .A(n_163), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_163), .A2(n_329), .B1(n_675), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_164), .A2(n_285), .B1(n_830), .B2(n_1226), .Y(n_1355) );
BUFx3_ASAP7_75t_L g404 ( .A(n_166), .Y(n_404) );
INVx1_ASAP7_75t_L g422 ( .A(n_166), .Y(n_422) );
INVx1_ASAP7_75t_L g807 ( .A(n_167), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_167), .A2(n_248), .B1(n_425), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g424 ( .A(n_168), .Y(n_424) );
INVx1_ASAP7_75t_L g1601 ( .A(n_169), .Y(n_1601) );
INVx1_ASAP7_75t_L g795 ( .A(n_170), .Y(n_795) );
INVx1_ASAP7_75t_L g414 ( .A(n_171), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g1307 ( .A1(n_172), .A2(n_236), .B1(n_682), .B2(n_1061), .Y(n_1307) );
AOI22xp33_ASAP7_75t_SL g1315 ( .A1(n_172), .A2(n_236), .B1(n_1184), .B2(n_1226), .Y(n_1315) );
INVx1_ASAP7_75t_L g1782 ( .A(n_173), .Y(n_1782) );
INVx1_ASAP7_75t_L g1010 ( .A(n_174), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_175), .A2(n_355), .B1(n_672), .B2(n_817), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_175), .A2(n_355), .B1(n_635), .B2(n_698), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g1442 ( .A1(n_176), .A2(n_336), .B1(n_1015), .B2(n_1017), .Y(n_1442) );
AOI221xp5_ASAP7_75t_L g1452 ( .A1(n_176), .A2(n_336), .B1(n_677), .B2(n_1453), .C(n_1456), .Y(n_1452) );
INVx1_ASAP7_75t_L g1287 ( .A(n_177), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_177), .A2(n_308), .B1(n_1231), .B2(n_1309), .Y(n_1312) );
INVxp33_ASAP7_75t_L g1147 ( .A(n_178), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_178), .A2(n_238), .B1(n_700), .B2(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g857 ( .A(n_179), .Y(n_857) );
INVx1_ASAP7_75t_L g1012 ( .A(n_180), .Y(n_1012) );
INVxp33_ASAP7_75t_L g407 ( .A(n_181), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_181), .A2(n_300), .B1(n_488), .B2(n_490), .C(n_492), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_182), .A2(n_231), .B1(n_677), .B2(n_680), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_182), .A2(n_231), .B1(n_694), .B2(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g1156 ( .A(n_183), .Y(n_1156) );
INVx1_ASAP7_75t_L g1524 ( .A(n_184), .Y(n_1524) );
INVx1_ASAP7_75t_L g788 ( .A(n_185), .Y(n_788) );
INVx1_ASAP7_75t_L g856 ( .A(n_186), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_187), .A2(n_352), .B1(n_671), .B2(n_673), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_187), .A2(n_352), .B1(n_635), .B2(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g659 ( .A(n_188), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_189), .A2(n_288), .B1(n_536), .B2(n_1504), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_189), .A2(n_288), .B1(n_677), .B2(n_1113), .Y(n_1513) );
INVx1_ASAP7_75t_L g958 ( .A(n_190), .Y(n_958) );
INVx1_ASAP7_75t_L g1602 ( .A(n_191), .Y(n_1602) );
XNOR2xp5_ASAP7_75t_L g1762 ( .A(n_191), .B(n_1763), .Y(n_1762) );
AOI22xp33_ASAP7_75t_L g1800 ( .A1(n_191), .A2(n_1801), .B1(n_1805), .B2(n_1809), .Y(n_1800) );
INVx1_ASAP7_75t_L g1389 ( .A(n_193), .Y(n_1389) );
OAI211xp5_ASAP7_75t_SL g1415 ( .A1(n_193), .A2(n_810), .B(n_1367), .C(n_1416), .Y(n_1415) );
AO22x2_ASAP7_75t_L g950 ( .A1(n_194), .A2(n_951), .B1(n_991), .B2(n_992), .Y(n_950) );
INVx1_ASAP7_75t_L g991 ( .A(n_194), .Y(n_991) );
INVxp33_ASAP7_75t_SL g569 ( .A(n_195), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_196), .A2(n_289), .B1(n_1015), .B2(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1233 ( .A(n_196), .Y(n_1233) );
INVx1_ASAP7_75t_L g1302 ( .A(n_197), .Y(n_1302) );
INVx1_ASAP7_75t_L g443 ( .A(n_198), .Y(n_443) );
INVxp33_ASAP7_75t_SL g800 ( .A(n_199), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_199), .A2(n_230), .B1(n_694), .B2(n_839), .Y(n_838) );
INVxp67_ASAP7_75t_L g1264 ( .A(n_200), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_200), .A2(n_294), .B1(n_1184), .B2(n_1185), .Y(n_1281) );
INVx1_ASAP7_75t_L g1057 ( .A(n_201), .Y(n_1057) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_201), .A2(n_326), .B1(n_711), .B2(n_740), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g1336 ( .A(n_203), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_203), .A2(n_328), .B1(n_704), .B2(n_1226), .Y(n_1350) );
INVx1_ASAP7_75t_L g1560 ( .A(n_204), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_206), .A2(n_349), .B1(n_682), .B2(n_1061), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_206), .A2(n_349), .B1(n_638), .B2(n_945), .Y(n_1071) );
INVx1_ASAP7_75t_L g863 ( .A(n_207), .Y(n_863) );
CKINVDCx14_ASAP7_75t_R g1190 ( .A(n_208), .Y(n_1190) );
INVx1_ASAP7_75t_L g1199 ( .A(n_209), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1575 ( .A1(n_210), .A2(n_295), .B1(n_1566), .B2(n_1569), .Y(n_1575) );
INVxp33_ASAP7_75t_SL g654 ( .A(n_211), .Y(n_654) );
INVxp33_ASAP7_75t_L g597 ( .A(n_212), .Y(n_597) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_213), .Y(n_743) );
INVx1_ASAP7_75t_L g1391 ( .A(n_214), .Y(n_1391) );
OAI22xp5_ASAP7_75t_L g1766 ( .A1(n_215), .A2(n_307), .B1(n_1194), .B2(n_1202), .Y(n_1766) );
INVx1_ASAP7_75t_L g1777 ( .A(n_215), .Y(n_1777) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_216), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_217), .Y(n_1448) );
INVxp33_ASAP7_75t_L g954 ( .A(n_218), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_218), .A2(n_312), .B1(n_638), .B2(n_830), .Y(n_990) );
INVxp33_ASAP7_75t_L g971 ( .A(n_219), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_219), .A2(n_278), .B1(n_460), .B2(n_490), .Y(n_978) );
INVx1_ASAP7_75t_L g656 ( .A(n_220), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_221), .A2(n_345), .B1(n_583), .B2(n_614), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_221), .A2(n_345), .B1(n_661), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g868 ( .A(n_223), .Y(n_868) );
INVx1_ASAP7_75t_L g1099 ( .A(n_225), .Y(n_1099) );
INVx1_ASAP7_75t_L g1331 ( .A(n_226), .Y(n_1331) );
INVxp33_ASAP7_75t_SL g911 ( .A(n_227), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_227), .A2(n_241), .B1(n_737), .B2(n_762), .Y(n_932) );
CKINVDCx16_ASAP7_75t_R g1556 ( .A(n_229), .Y(n_1556) );
INVxp33_ASAP7_75t_SL g801 ( .A(n_230), .Y(n_801) );
INVxp33_ASAP7_75t_SL g786 ( .A(n_232), .Y(n_786) );
INVx1_ASAP7_75t_L g1208 ( .A(n_235), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_237), .A2(n_243), .B1(n_1194), .B2(n_1202), .Y(n_1441) );
INVx1_ASAP7_75t_L g1457 ( .A(n_237), .Y(n_1457) );
INVxp67_ASAP7_75t_SL g1144 ( .A(n_238), .Y(n_1144) );
INVx1_ASAP7_75t_L g902 ( .A(n_241), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_242), .Y(n_482) );
INVx1_ASAP7_75t_L g1433 ( .A(n_243), .Y(n_1433) );
INVx1_ASAP7_75t_L g1496 ( .A(n_244), .Y(n_1496) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_244), .A2(n_293), .B1(n_675), .B2(n_685), .Y(n_1515) );
INVxp67_ASAP7_75t_SL g1126 ( .A(n_246), .Y(n_1126) );
INVx1_ASAP7_75t_L g1392 ( .A(n_247), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_247), .A2(n_258), .B1(n_606), .B2(n_1239), .Y(n_1414) );
INVxp33_ASAP7_75t_SL g809 ( .A(n_248), .Y(n_809) );
INVxp33_ASAP7_75t_L g1261 ( .A(n_249), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1774 ( .A(n_250), .Y(n_1774) );
INVx1_ASAP7_75t_L g1487 ( .A(n_251), .Y(n_1487) );
INVxp33_ASAP7_75t_L g717 ( .A(n_252), .Y(n_717) );
BUFx3_ASAP7_75t_L g406 ( .A(n_253), .Y(n_406) );
INVx1_ASAP7_75t_L g412 ( .A(n_253), .Y(n_412) );
INVx1_ASAP7_75t_L g1224 ( .A(n_254), .Y(n_1224) );
INVx1_ASAP7_75t_L g1050 ( .A(n_255), .Y(n_1050) );
INVx1_ASAP7_75t_L g1055 ( .A(n_257), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_258), .A2(n_266), .B1(n_1194), .B2(n_1202), .Y(n_1408) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_259), .Y(n_374) );
AND2x2_ASAP7_75t_L g450 ( .A(n_259), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_259), .B(n_334), .Y(n_473) );
INVx1_ASAP7_75t_L g505 ( .A(n_259), .Y(n_505) );
INVx1_ASAP7_75t_L g433 ( .A(n_261), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_261), .A2(n_358), .B1(n_466), .B2(n_474), .C(n_476), .Y(n_465) );
AOI221xp5_ASAP7_75t_SL g1445 ( .A1(n_262), .A2(n_276), .B1(n_1113), .B2(n_1446), .C(n_1447), .Y(n_1445) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_262), .A2(n_276), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
AO22x2_ASAP7_75t_L g781 ( .A1(n_263), .A2(n_782), .B1(n_840), .B2(n_841), .Y(n_781) );
INVx1_ASAP7_75t_L g840 ( .A(n_263), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_264), .A2(n_309), .B1(n_762), .B2(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_264), .A2(n_309), .B1(n_768), .B2(n_877), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_265), .Y(n_1362) );
INVx1_ASAP7_75t_L g1402 ( .A(n_266), .Y(n_1402) );
XNOR2xp5_ASAP7_75t_L g1371 ( .A(n_268), .B(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1561 ( .A(n_268), .Y(n_1561) );
INVx2_ASAP7_75t_L g399 ( .A(n_270), .Y(n_399) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_271), .Y(n_456) );
INVx1_ASAP7_75t_L g1244 ( .A(n_272), .Y(n_1244) );
INVx1_ASAP7_75t_L g1536 ( .A(n_273), .Y(n_1536) );
INVx1_ASAP7_75t_L g872 ( .A(n_274), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_274), .A2(n_283), .B1(n_877), .B2(n_879), .Y(n_876) );
INVx1_ASAP7_75t_L g728 ( .A(n_275), .Y(n_728) );
INVx1_ASAP7_75t_L g578 ( .A(n_277), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_277), .A2(n_314), .B1(n_589), .B2(n_591), .Y(n_588) );
INVxp33_ASAP7_75t_L g969 ( .A(n_278), .Y(n_969) );
INVx1_ASAP7_75t_L g1412 ( .A(n_280), .Y(n_1412) );
CKINVDCx16_ASAP7_75t_R g1558 ( .A(n_281), .Y(n_1558) );
AOI22xp5_ASAP7_75t_L g1806 ( .A1(n_282), .A2(n_1763), .B1(n_1807), .B2(n_1808), .Y(n_1806) );
CKINVDCx5p33_ASAP7_75t_R g1807 ( .A(n_282), .Y(n_1807) );
INVx1_ASAP7_75t_L g866 ( .A(n_283), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_285), .A2(n_323), .B1(n_606), .B2(n_1239), .Y(n_1365) );
INVx1_ASAP7_75t_L g734 ( .A(n_286), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_287), .Y(n_1449) );
INVx1_ASAP7_75t_L g1212 ( .A(n_289), .Y(n_1212) );
INVx1_ASAP7_75t_L g1584 ( .A(n_290), .Y(n_1584) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_291), .Y(n_738) );
INVx1_ASAP7_75t_L g1339 ( .A(n_292), .Y(n_1339) );
INVxp33_ASAP7_75t_SL g1494 ( .A(n_293), .Y(n_1494) );
INVx1_ASAP7_75t_L g1262 ( .A(n_294), .Y(n_1262) );
INVx1_ASAP7_75t_L g791 ( .A(n_296), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_297), .A2(n_333), .B1(n_749), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_297), .A2(n_333), .B1(n_828), .B2(n_831), .Y(n_827) );
INVx1_ASAP7_75t_L g1354 ( .A(n_298), .Y(n_1354) );
OAI211xp5_ASAP7_75t_SL g1366 ( .A1(n_298), .A2(n_810), .B(n_1367), .C(n_1369), .Y(n_1366) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_300), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_301), .A2(n_331), .B1(n_848), .B2(n_854), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_301), .A2(n_331), .B1(n_589), .B2(n_591), .Y(n_1259) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_302), .Y(n_909) );
INVx1_ASAP7_75t_L g665 ( .A(n_303), .Y(n_665) );
INVx1_ASAP7_75t_L g1301 ( .A(n_304), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_304), .A2(n_338), .B1(n_732), .B2(n_1070), .Y(n_1317) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_305), .Y(n_906) );
INVxp67_ASAP7_75t_SL g1013 ( .A(n_306), .Y(n_1013) );
INVx1_ASAP7_75t_L g1293 ( .A(n_308), .Y(n_1293) );
INVx1_ASAP7_75t_L g1136 ( .A(n_310), .Y(n_1136) );
INVxp33_ASAP7_75t_L g955 ( .A(n_312), .Y(n_955) );
INVx1_ASAP7_75t_L g1381 ( .A(n_313), .Y(n_1381) );
INVx1_ASAP7_75t_L g577 ( .A(n_314), .Y(n_577) );
INVx1_ASAP7_75t_L g961 ( .A(n_315), .Y(n_961) );
INVxp67_ASAP7_75t_SL g1152 ( .A(n_316), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_316), .A2(n_337), .B1(n_684), .B2(n_1167), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
AND3x2_ASAP7_75t_L g1530 ( .A(n_317), .B(n_366), .C(n_1531), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_317), .B(n_366), .Y(n_1540) );
INVxp33_ASAP7_75t_SL g1092 ( .A(n_318), .Y(n_1092) );
INVx2_ASAP7_75t_L g379 ( .A(n_319), .Y(n_379) );
INVx1_ASAP7_75t_L g967 ( .A(n_321), .Y(n_967) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_322), .A2(n_478), .B(n_481), .Y(n_477) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_322), .Y(n_532) );
INVx1_ASAP7_75t_L g513 ( .A(n_325), .Y(n_513) );
INVx1_ASAP7_75t_L g1056 ( .A(n_326), .Y(n_1056) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_327), .Y(n_917) );
INVxp67_ASAP7_75t_SL g1333 ( .A(n_328), .Y(n_1333) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_329), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g1769 ( .A(n_330), .Y(n_1769) );
INVx1_ASAP7_75t_L g1328 ( .A(n_332), .Y(n_1328) );
INVx1_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
INVx2_ASAP7_75t_L g451 ( .A(n_334), .Y(n_451) );
XNOR2xp5_ASAP7_75t_L g1283 ( .A(n_335), .B(n_1284), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_337), .Y(n_1154) );
INVx1_ASAP7_75t_L g1298 ( .A(n_338), .Y(n_1298) );
INVx1_ASAP7_75t_L g510 ( .A(n_340), .Y(n_510) );
INVxp33_ASAP7_75t_L g729 ( .A(n_341), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_342), .Y(n_1430) );
CKINVDCx5p33_ASAP7_75t_R g1770 ( .A(n_344), .Y(n_1770) );
AO22x2_ASAP7_75t_L g1478 ( .A1(n_346), .A2(n_1479), .B1(n_1480), .B2(n_1516), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_346), .Y(n_1479) );
XOR2x2_ASAP7_75t_L g563 ( .A(n_348), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g1291 ( .A(n_351), .Y(n_1291) );
INVx1_ASAP7_75t_L g1085 ( .A(n_353), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_354), .A2(n_357), .B1(n_703), .B2(n_705), .Y(n_702) );
INVxp33_ASAP7_75t_L g713 ( .A(n_354), .Y(n_713) );
INVx1_ASAP7_75t_L g1345 ( .A(n_356), .Y(n_1345) );
INVxp67_ASAP7_75t_SL g715 ( .A(n_357), .Y(n_715) );
INVx1_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
AO22x1_ASAP7_75t_L g720 ( .A1(n_359), .A2(n_721), .B1(n_722), .B2(n_777), .Y(n_720) );
INVxp67_ASAP7_75t_L g721 ( .A(n_359), .Y(n_721) );
AOI21xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_382), .B(n_1518), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_369), .Y(n_363) );
AND2x4_ASAP7_75t_L g1799 ( .A(n_364), .B(n_370), .Y(n_1799) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_SL g1804 ( .A(n_365), .Y(n_1804) );
NAND2xp5_ASAP7_75t_L g1811 ( .A(n_365), .B(n_367), .Y(n_1811) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_367), .B(n_1804), .Y(n_1803) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x6_ASAP7_75t_L g608 ( .A(n_372), .B(n_558), .Y(n_608) );
OR2x2_ASAP7_75t_L g924 ( .A(n_372), .B(n_558), .Y(n_924) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g483 ( .A(n_373), .B(n_381), .Y(n_483) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_374), .B(n_596), .Y(n_1325) );
INVx8_ASAP7_75t_L g604 ( .A(n_375), .Y(n_604) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_376), .A2(n_482), .B(n_483), .Y(n_481) );
OR2x6_ASAP7_75t_L g606 ( .A(n_376), .B(n_595), .Y(n_606) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_376), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_376), .Y(n_1214) );
BUFx6f_ASAP7_75t_L g1327 ( .A(n_376), .Y(n_1327) );
INVx2_ASAP7_75t_SL g1397 ( .A(n_376), .Y(n_1397) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g453 ( .A(n_378), .Y(n_453) );
AND2x4_ASAP7_75t_L g462 ( .A(n_378), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g480 ( .A(n_378), .Y(n_480) );
INVx1_ASAP7_75t_L g496 ( .A(n_378), .Y(n_496) );
AND2x2_ASAP7_75t_L g500 ( .A(n_378), .B(n_379), .Y(n_500) );
INVx1_ASAP7_75t_L g455 ( .A(n_379), .Y(n_455) );
INVx2_ASAP7_75t_L g463 ( .A(n_379), .Y(n_463) );
INVx1_ASAP7_75t_L g469 ( .A(n_379), .Y(n_469) );
INVx1_ASAP7_75t_L g495 ( .A(n_379), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_379), .B(n_453), .Y(n_1238) );
AND2x4_ASAP7_75t_L g590 ( .A(n_380), .B(n_469), .Y(n_590) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g591 ( .A(n_381), .B(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g711 ( .A(n_381), .B(n_592), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_1131), .B2(n_1132), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_995), .B2(n_996), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
XNOR2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_779), .Y(n_386) );
XNOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_647), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_561), .B2(n_646), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221x1_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_440), .B1(n_446), .B2(n_519), .C(n_523), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_394), .B(n_413), .C(n_423), .D(n_436), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_407), .B2(n_408), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_396), .A2(n_408), .B1(n_725), .B2(n_726), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_396), .A2(n_408), .B1(n_856), .B2(n_857), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g970 ( .A1(n_396), .A2(n_408), .B1(n_971), .B2(n_972), .Y(n_970) );
AOI22xp5_ASAP7_75t_SL g1286 ( .A1(n_396), .A2(n_415), .B1(n_1287), .B2(n_1288), .Y(n_1286) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
AND2x6_ASAP7_75t_L g419 ( .A(n_397), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g568 ( .A(n_397), .B(n_400), .Y(n_568) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g849 ( .A(n_398), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g410 ( .A(n_399), .Y(n_410) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
AND2x2_ASAP7_75t_L g544 ( .A(n_399), .B(n_443), .Y(n_544) );
INVx2_ASAP7_75t_L g560 ( .A(n_399), .Y(n_560) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_401), .Y(n_634) );
INVx2_ASAP7_75t_L g701 ( .A(n_401), .Y(n_701) );
INVx2_ASAP7_75t_SL g767 ( .A(n_401), .Y(n_767) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_401), .Y(n_837) );
INVx2_ASAP7_75t_L g878 ( .A(n_401), .Y(n_878) );
INVx1_ASAP7_75t_L g1276 ( .A(n_401), .Y(n_1276) );
INVx6_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g415 ( .A(n_402), .B(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g773 ( .A(n_402), .Y(n_773) );
INVx2_ASAP7_75t_L g989 ( .A(n_402), .Y(n_989) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g411 ( .A(n_404), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g427 ( .A(n_404), .B(n_406), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g421 ( .A(n_406), .B(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_408), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_408), .A2(n_568), .B1(n_653), .B2(n_654), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_408), .A2(n_568), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_408), .A2(n_568), .B1(n_911), .B2(n_912), .Y(n_910) );
CKINVDCx6p67_ASAP7_75t_R g1017 ( .A(n_408), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_408), .A2(n_568), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_408), .A2(n_437), .B1(n_568), .B2(n_1091), .C(n_1092), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_408), .A2(n_568), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_408), .A2(n_419), .B1(n_1254), .B2(n_1255), .Y(n_1253) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_408), .A2(n_419), .B1(n_1290), .B2(n_1291), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_408), .A2(n_1498), .B1(n_1499), .B2(n_1500), .Y(n_1497) );
AND2x6_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g438 ( .A(n_409), .Y(n_438) );
INVx1_ASAP7_75t_L g1016 ( .A(n_409), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_409), .B(n_661), .Y(n_1197) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x6_ASAP7_75t_L g434 ( .A(n_410), .B(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_411), .Y(n_535) );
BUFx2_ASAP7_75t_L g637 ( .A(n_411), .Y(n_637) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_411), .Y(n_694) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_411), .Y(n_704) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_411), .Y(n_775) );
BUFx6f_ASAP7_75t_L g830 ( .A(n_411), .Y(n_830) );
INVx2_ASAP7_75t_SL g946 ( .A(n_411), .Y(n_946) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_411), .Y(n_1042) );
BUFx6f_ASAP7_75t_L g1176 ( .A(n_411), .Y(n_1176) );
BUFx3_ASAP7_75t_L g1184 ( .A(n_411), .Y(n_1184) );
INVx1_ASAP7_75t_L g529 ( .A(n_412), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_418), .B2(n_419), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g509 ( .A1(n_414), .A2(n_510), .B1(n_511), .B2(n_513), .C1(n_514), .C2(n_516), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_415), .A2(n_419), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_415), .A2(n_419), .B1(n_656), .B2(n_657), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_415), .A2(n_419), .B1(n_728), .B2(n_729), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_415), .A2(n_419), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_415), .A2(n_419), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_415), .A2(n_419), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_415), .A2(n_419), .B1(n_437), .B2(n_964), .C(n_969), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_415), .A2(n_419), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_415), .A2(n_419), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_415), .A2(n_419), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_415), .A2(n_419), .B1(n_1140), .B2(n_1154), .Y(n_1153) );
INVx4_ASAP7_75t_L g1194 ( .A(n_415), .Y(n_1194) );
AOI22xp5_ASAP7_75t_SL g1247 ( .A1(n_415), .A2(n_568), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_415), .A2(n_419), .B1(n_1491), .B2(n_1494), .Y(n_1493) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_416), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g664 ( .A(n_416), .B(n_430), .Y(n_664) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx4_ASAP7_75t_L g1202 ( .A(n_419), .Y(n_1202) );
INVx1_ASAP7_75t_L g554 ( .A(n_420), .Y(n_554) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_420), .Y(n_638) );
INVx2_ASAP7_75t_L g832 ( .A(n_420), .Y(n_832) );
INVx1_ASAP7_75t_L g939 ( .A(n_420), .Y(n_939) );
INVx1_ASAP7_75t_L g1076 ( .A(n_420), .Y(n_1076) );
BUFx6f_ASAP7_75t_L g1185 ( .A(n_420), .Y(n_1185) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g539 ( .A(n_421), .Y(n_539) );
INVx1_ASAP7_75t_L g696 ( .A(n_421), .Y(n_696) );
BUFx6f_ASAP7_75t_L g1226 ( .A(n_421), .Y(n_1226) );
INVx1_ASAP7_75t_L g528 ( .A(n_422), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_428), .B2(n_429), .C1(n_433), .C2(n_434), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g492 ( .A1(n_424), .A2(n_493), .B(n_497), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g1054 ( .A1(n_425), .A2(n_429), .B1(n_434), .B2(n_1055), .C1(n_1056), .C2(n_1057), .Y(n_1054) );
BUFx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx4f_ASAP7_75t_L g635 ( .A(n_426), .Y(n_635) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_426), .Y(n_732) );
INVx2_ASAP7_75t_SL g880 ( .A(n_426), .Y(n_880) );
INVx1_ASAP7_75t_L g943 ( .A(n_426), .Y(n_943) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_427), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_429), .A2(n_434), .B1(n_574), .B2(n_575), .C1(n_577), .C2(n_578), .Y(n_573) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_429), .A2(n_434), .B1(n_731), .B2(n_732), .C1(n_733), .C2(n_734), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g966 ( .A1(n_429), .A2(n_434), .B1(n_575), .B2(n_958), .C1(n_961), .C2(n_967), .Y(n_966) );
AOI222xp33_ASAP7_75t_L g1093 ( .A1(n_429), .A2(n_434), .B1(n_1094), .B2(n_1095), .C1(n_1096), .C2(n_1097), .Y(n_1093) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g850 ( .A(n_431), .Y(n_850) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI222xp33_ASAP7_75t_L g658 ( .A1(n_434), .A2(n_659), .B1(n_660), .B2(n_662), .C1(n_663), .C2(n_665), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g790 ( .A1(n_434), .A2(n_663), .B1(n_791), .B2(n_792), .C1(n_795), .C2(n_796), .Y(n_790) );
INVx3_ASAP7_75t_L g854 ( .A(n_434), .Y(n_854) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_434), .A2(n_664), .B1(n_902), .B2(n_903), .C1(n_905), .C2(n_906), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_434), .A2(n_849), .B1(n_1009), .B2(n_1010), .Y(n_1008) );
AOI222xp33_ASAP7_75t_L g1155 ( .A1(n_434), .A2(n_663), .B1(n_1143), .B2(n_1145), .C1(n_1156), .C2(n_1157), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_434), .A2(n_664), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
AOI222xp33_ASAP7_75t_L g1359 ( .A1(n_434), .A2(n_849), .B1(n_1345), .B2(n_1360), .C1(n_1361), .C2(n_1362), .Y(n_1359) );
AOI222xp33_ASAP7_75t_L g1410 ( .A1(n_434), .A2(n_768), .B1(n_849), .B2(n_1405), .C1(n_1411), .C2(n_1412), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_434), .A2(n_663), .B1(n_1428), .B2(n_1430), .Y(n_1439) );
AOI222xp33_ASAP7_75t_L g1495 ( .A1(n_434), .A2(n_663), .B1(n_1157), .B2(n_1487), .C1(n_1488), .C2(n_1496), .Y(n_1495) );
AOI22xp33_ASAP7_75t_L g1768 ( .A1(n_434), .A2(n_664), .B1(n_1769), .B2(n_1770), .Y(n_1768) );
NAND4xp25_ASAP7_75t_SL g651 ( .A(n_436), .B(n_652), .C(n_655), .D(n_658), .Y(n_651) );
NAND4xp25_ASAP7_75t_SL g723 ( .A(n_436), .B(n_724), .C(n_727), .D(n_730), .Y(n_723) );
BUFx2_ASAP7_75t_L g797 ( .A(n_436), .Y(n_797) );
NAND4xp25_ASAP7_75t_L g1047 ( .A(n_436), .B(n_1048), .C(n_1051), .D(n_1054), .Y(n_1047) );
NAND4xp25_ASAP7_75t_L g1149 ( .A(n_436), .B(n_1150), .C(n_1153), .D(n_1155), .Y(n_1149) );
NAND4xp25_ASAP7_75t_L g1246 ( .A(n_436), .B(n_1247), .C(n_1250), .D(n_1253), .Y(n_1246) );
NAND4xp25_ASAP7_75t_L g1285 ( .A(n_436), .B(n_1286), .C(n_1289), .D(n_1292), .Y(n_1285) );
INVx5_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx8_ASAP7_75t_R g579 ( .A(n_437), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_437), .B(n_847), .Y(n_846) );
NOR2xp33_ASAP7_75t_SL g1003 ( .A(n_437), .B(n_1004), .Y(n_1003) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_439), .Y(n_576) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_439), .Y(n_661) );
INVx2_ASAP7_75t_L g769 ( .A(n_439), .Y(n_769) );
INVx1_ASAP7_75t_L g904 ( .A(n_439), .Y(n_904) );
AOI211x1_ASAP7_75t_SL g650 ( .A1(n_440), .A2(n_651), .B(n_666), .C(n_707), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g722 ( .A1(n_440), .A2(n_723), .B(n_735), .C(n_746), .Y(n_722) );
AOI221x1_ASAP7_75t_L g782 ( .A1(n_440), .A2(n_607), .B1(n_783), .B2(n_798), .C(n_811), .Y(n_782) );
AOI221x1_ASAP7_75t_L g844 ( .A1(n_440), .A2(n_607), .B1(n_845), .B2(n_861), .C(n_874), .Y(n_844) );
INVx1_ASAP7_75t_L g1443 ( .A(n_440), .Y(n_1443) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_441), .A2(n_565), .B1(n_580), .B2(n_607), .C(n_609), .Y(n_564) );
AOI211x1_ASAP7_75t_SL g899 ( .A1(n_441), .A2(n_900), .B(n_913), .C(n_925), .Y(n_899) );
AOI221x1_ASAP7_75t_L g951 ( .A1(n_441), .A2(n_607), .B1(n_952), .B2(n_965), .C(n_973), .Y(n_951) );
OAI21xp5_ASAP7_75t_L g1001 ( .A1(n_441), .A2(n_1002), .B(n_1014), .Y(n_1001) );
INVx1_ASAP7_75t_L g1101 ( .A(n_441), .Y(n_1101) );
AOI221x1_ASAP7_75t_L g1480 ( .A1(n_441), .A2(n_607), .B1(n_1481), .B2(n_1492), .C(n_1501), .Y(n_1480) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
AND2x4_ASAP7_75t_L g1046 ( .A(n_442), .B(n_444), .Y(n_1046) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g559 ( .A(n_443), .B(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g522 ( .A(n_445), .Y(n_522) );
OR2x6_ASAP7_75t_L g1324 ( .A(n_445), .B(n_1325), .Y(n_1324) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_464), .C(n_509), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_456), .B2(n_457), .Y(n_447) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx2_ASAP7_75t_L g459 ( .A(n_450), .Y(n_459) );
AND2x4_ASAP7_75t_L g514 ( .A(n_450), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g504 ( .A(n_451), .Y(n_504) );
INVx1_ASAP7_75t_L g596 ( .A(n_451), .Y(n_596) );
INVx1_ASAP7_75t_L g491 ( .A(n_452), .Y(n_491) );
AND2x4_ASAP7_75t_L g594 ( .A(n_452), .B(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_452), .Y(n_612) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_452), .Y(n_679) );
BUFx2_ASAP7_75t_L g684 ( .A(n_452), .Y(n_684) );
BUFx2_ASAP7_75t_L g749 ( .A(n_452), .Y(n_749) );
INVx1_ASAP7_75t_L g758 ( .A(n_452), .Y(n_758) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_452), .Y(n_1061) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g475 ( .A(n_453), .Y(n_475) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
AND2x4_ASAP7_75t_L g511 ( .A(n_458), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g623 ( .A(n_460), .Y(n_623) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g891 ( .A(n_461), .Y(n_891) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g486 ( .A(n_462), .Y(n_486) );
INVx1_ASAP7_75t_L g600 ( .A(n_462), .Y(n_600) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_462), .Y(n_682) );
AND2x4_ASAP7_75t_L g479 ( .A(n_463), .B(n_480), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_487), .C(n_506), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g474 ( .A(n_471), .B(n_475), .Y(n_474) );
OR2x6_ASAP7_75t_L g507 ( .A(n_471), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_484), .Y(n_476) );
INVx2_ASAP7_75t_SL g629 ( .A(n_478), .Y(n_629) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_478), .Y(n_754) );
BUFx2_ASAP7_75t_L g1032 ( .A(n_478), .Y(n_1032) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g512 ( .A(n_479), .Y(n_512) );
AND2x4_ASAP7_75t_L g585 ( .A(n_479), .B(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_479), .Y(n_675) );
BUFx2_ASAP7_75t_L g689 ( .A(n_479), .Y(n_689) );
INVx1_ASAP7_75t_L g919 ( .A(n_479), .Y(n_919) );
BUFx3_ASAP7_75t_L g1231 ( .A(n_479), .Y(n_1231) );
OAI221xp5_ASAP7_75t_SL g524 ( .A1(n_482), .A2(n_525), .B1(n_530), .B2(n_532), .C(n_533), .Y(n_524) );
AND2x4_ASAP7_75t_L g630 ( .A(n_483), .B(n_522), .Y(n_630) );
AND2x4_ASAP7_75t_L g928 ( .A(n_483), .B(n_522), .Y(n_928) );
INVx2_ASAP7_75t_L g751 ( .A(n_485), .Y(n_751) );
INVx2_ASAP7_75t_L g760 ( .A(n_485), .Y(n_760) );
INVx1_ASAP7_75t_L g1337 ( .A(n_485), .Y(n_1337) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_486), .Y(n_489) );
INVx3_ASAP7_75t_L g1114 ( .A(n_486), .Y(n_1114) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g1065 ( .A(n_489), .Y(n_1065) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g934 ( .A(n_491), .Y(n_934) );
INVx1_ASAP7_75t_L g1030 ( .A(n_491), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g1205 ( .A1(n_493), .A2(n_1206), .B1(n_1207), .B2(n_1208), .Y(n_1205) );
OAI22xp33_ASAP7_75t_SL g1211 ( .A1(n_493), .A2(n_1212), .B1(n_1213), .B2(n_1215), .Y(n_1211) );
OAI22xp33_ASAP7_75t_L g1403 ( .A1(n_493), .A2(n_1396), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g1786 ( .A1(n_493), .A2(n_1327), .B1(n_1787), .B2(n_1788), .Y(n_1786) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g508 ( .A(n_494), .Y(n_508) );
INVx2_ASAP7_75t_L g1344 ( .A(n_494), .Y(n_1344) );
BUFx2_ASAP7_75t_L g1368 ( .A(n_494), .Y(n_1368) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_495), .B(n_496), .Y(n_1330) );
INVx1_ASAP7_75t_L g592 ( .A(n_496), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_498), .B(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g753 ( .A(n_498), .Y(n_753) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g627 ( .A(n_499), .Y(n_627) );
INVx2_ASAP7_75t_L g672 ( .A(n_499), .Y(n_672) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_500), .Y(n_515) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g981 ( .A(n_502), .B(n_522), .Y(n_981) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x6_ASAP7_75t_L g617 ( .A(n_503), .B(n_618), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g587 ( .A(n_504), .Y(n_587) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI221xp5_ASAP7_75t_SL g545 ( .A1(n_510), .A2(n_513), .B1(n_546), .B2(n_549), .C(n_552), .Y(n_545) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_512), .Y(n_583) );
INVx1_ASAP7_75t_L g894 ( .A(n_512), .Y(n_894) );
INVx3_ASAP7_75t_L g615 ( .A(n_515), .Y(n_615) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_515), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g1455 ( .A(n_515), .Y(n_1455) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
CKINVDCx8_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x6_ASAP7_75t_L g542 ( .A(n_522), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g640 ( .A(n_522), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_522), .B(n_543), .Y(n_1217) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_540), .B1(n_545), .B2(n_555), .Y(n_523) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g548 ( .A(n_527), .Y(n_548) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_527), .B(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1383 ( .A(n_527), .Y(n_1383) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g531 ( .A(n_528), .B(n_529), .Y(n_531) );
BUFx3_ASAP7_75t_L g1220 ( .A(n_530), .Y(n_1220) );
INVx1_ASAP7_75t_L g1438 ( .A(n_530), .Y(n_1438) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g551 ( .A(n_531), .Y(n_551) );
INVx1_ASAP7_75t_L g853 ( .A(n_531), .Y(n_853) );
INVx1_ASAP7_75t_L g1007 ( .A(n_531), .Y(n_1007) );
BUFx4f_ASAP7_75t_L g1386 ( .A(n_531), .Y(n_1386) );
BUFx4f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g1377 ( .A(n_535), .Y(n_1377) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g776 ( .A(n_537), .Y(n_776) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g705 ( .A(n_539), .Y(n_705) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI33xp33_ASAP7_75t_L g936 ( .A1(n_541), .A2(n_645), .A3(n_937), .B1(n_940), .B2(n_941), .B3(n_944), .Y(n_936) );
AOI33xp33_ASAP7_75t_L g1033 ( .A1(n_541), .A2(n_556), .A3(n_1034), .B1(n_1038), .B2(n_1040), .B3(n_1041), .Y(n_1033) );
AOI33xp33_ASAP7_75t_L g1502 ( .A1(n_541), .A2(n_1179), .A3(n_1503), .B1(n_1505), .B2(n_1508), .B3(n_1509), .Y(n_1502) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_542), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_542), .Y(n_833) );
OAI22xp5_ASAP7_75t_SL g1464 ( .A1(n_542), .A2(n_1180), .B1(n_1465), .B2(n_1469), .Y(n_1464) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g641 ( .A(n_544), .Y(n_641) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g1219 ( .A(n_548), .Y(n_1219) );
INVx2_ASAP7_75t_L g1349 ( .A(n_548), .Y(n_1349) );
INVx2_ASAP7_75t_L g1352 ( .A(n_548), .Y(n_1352) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_550), .A2(n_1352), .B1(n_1353), .B2(n_1354), .C(n_1355), .Y(n_1351) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
AOI33xp33_ASAP7_75t_L g875 ( .A1(n_556), .A2(n_639), .A3(n_876), .B1(n_881), .B2(n_882), .B3(n_883), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_556), .B(n_1104), .C(n_1105), .Y(n_1103) );
BUFx4f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx4f_ASAP7_75t_L g706 ( .A(n_557), .Y(n_706) );
INVx4_ASAP7_75t_L g1180 ( .A(n_557), .Y(n_1180) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x4_ASAP7_75t_L g645 ( .A(n_558), .B(n_559), .Y(n_645) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g646 ( .A(n_563), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .C(n_573), .D(n_579), .Y(n_565) );
HB1xp67_ASAP7_75t_L g1499 ( .A(n_568), .Y(n_1499) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_571), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND4xp25_ASAP7_75t_SL g900 ( .A(n_579), .B(n_901), .C(n_907), .D(n_910), .Y(n_900) );
NAND2xp5_ASAP7_75t_SL g1358 ( .A(n_579), .B(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_SL g1409 ( .A(n_579), .B(n_1410), .Y(n_1409) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_593), .C(n_602), .Y(n_580) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B(n_585), .C(n_588), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI211xp5_ASAP7_75t_L g708 ( .A1(n_583), .A2(n_585), .B(n_709), .C(n_710), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g1122 ( .A1(n_583), .A2(n_585), .B(n_1123), .C(n_1124), .Y(n_1122) );
AOI211xp5_ASAP7_75t_L g736 ( .A1(n_585), .A2(n_737), .B(n_738), .C(n_739), .Y(n_736) );
CKINVDCx11_ASAP7_75t_R g810 ( .A(n_585), .Y(n_810) );
AOI211xp5_ASAP7_75t_L g916 ( .A1(n_585), .A2(n_917), .B(n_918), .C(n_920), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g1019 ( .A(n_585), .B(n_1020), .C(n_1021), .Y(n_1019) );
AOI211xp5_ASAP7_75t_L g1078 ( .A1(n_585), .A2(n_737), .B(n_1079), .C(n_1080), .Y(n_1078) );
AOI211xp5_ASAP7_75t_L g1257 ( .A1(n_585), .A2(n_1230), .B(n_1258), .C(n_1259), .Y(n_1257) );
AOI211xp5_ASAP7_75t_L g1297 ( .A1(n_585), .A2(n_930), .B(n_1298), .C(n_1299), .Y(n_1297) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_L g806 ( .A(n_587), .Y(n_806) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g740 ( .A(n_590), .Y(n_740) );
INVx2_ASAP7_75t_L g960 ( .A(n_590), .Y(n_960) );
AOI222xp33_ASAP7_75t_L g1229 ( .A1(n_590), .A2(n_804), .B1(n_1199), .B2(n_1200), .C1(n_1224), .C2(n_1230), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1369 ( .A1(n_590), .A2(n_804), .B1(n_1361), .B2(n_1362), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_590), .A2(n_804), .B1(n_1411), .B2(n_1412), .Y(n_1416) );
AOI222xp33_ASAP7_75t_L g1427 ( .A1(n_590), .A2(n_675), .B1(n_804), .B2(n_1428), .C1(n_1429), .C2(n_1430), .Y(n_1427) );
AOI222xp33_ASAP7_75t_L g1485 ( .A1(n_590), .A2(n_804), .B1(n_867), .B2(n_1486), .C1(n_1487), .C2(n_1488), .Y(n_1485) );
AOI222xp33_ASAP7_75t_SL g1773 ( .A1(n_590), .A2(n_817), .B1(n_870), .B2(n_1769), .C1(n_1770), .C2(n_1774), .Y(n_1773) );
INVx1_ASAP7_75t_L g805 ( .A(n_592), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B1(n_598), .B2(n_601), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_594), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_594), .A2(n_598), .B1(n_742), .B2(n_743), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_594), .A2(n_598), .B1(n_800), .B2(n_801), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_594), .A2(n_714), .B1(n_863), .B2(n_864), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_594), .A2(n_714), .B1(n_922), .B2(n_923), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_594), .A2(n_598), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_594), .A2(n_598), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g1081 ( .A1(n_594), .A2(n_598), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
AOI22xp5_ASAP7_75t_SL g1127 ( .A1(n_594), .A2(n_598), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AOI22xp33_ASAP7_75t_SL g1139 ( .A1(n_594), .A2(n_873), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g1260 ( .A1(n_594), .A2(n_604), .B1(n_1261), .B2(n_1262), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_594), .A2(n_604), .B1(n_1301), .B2(n_1302), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_594), .A2(n_714), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
AND2x4_ASAP7_75t_L g598 ( .A(n_595), .B(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g714 ( .A(n_595), .B(n_599), .Y(n_714) );
INVx1_ASAP7_75t_L g1236 ( .A(n_595), .Y(n_1236) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_598), .A2(n_604), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_600), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_604), .A2(n_605), .B1(n_656), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_604), .A2(n_605), .B1(n_728), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_604), .A2(n_605), .B1(n_788), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_604), .A2(n_859), .B1(n_872), .B2(n_873), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_604), .A2(n_605), .B1(n_908), .B2(n_915), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_604), .A2(n_605), .B1(n_963), .B2(n_964), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_604), .A2(n_873), .B1(n_1049), .B2(n_1085), .Y(n_1084) );
AOI22xp5_ASAP7_75t_L g1125 ( .A1(n_604), .A2(n_873), .B1(n_1099), .B2(n_1126), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_604), .A2(n_873), .B1(n_1223), .B2(n_1233), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_604), .A2(n_605), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_604), .A2(n_873), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
AOI22xp33_ASAP7_75t_L g1775 ( .A1(n_604), .A2(n_873), .B1(n_1776), .B2(n_1777), .Y(n_1775) );
AOI22xp33_ASAP7_75t_SL g1263 ( .A1(n_605), .A2(n_714), .B1(n_1249), .B2(n_1264), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_605), .A2(n_714), .B1(n_1288), .B2(n_1304), .Y(n_1303) );
INVx5_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx4_ASAP7_75t_L g873 ( .A(n_606), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_607), .A2(n_1138), .B1(n_1149), .B2(n_1158), .C(n_1159), .Y(n_1137) );
OAI21xp5_ASAP7_75t_L g1227 ( .A1(n_607), .A2(n_1228), .B(n_1234), .Y(n_1227) );
OAI31xp33_ASAP7_75t_SL g1364 ( .A1(n_607), .A2(n_1365), .A3(n_1366), .B(n_1370), .Y(n_1364) );
OAI31xp33_ASAP7_75t_SL g1413 ( .A1(n_607), .A2(n_1414), .A3(n_1415), .B(n_1417), .Y(n_1413) );
O2A1O1Ixp33_ASAP7_75t_L g1424 ( .A1(n_607), .A2(n_1425), .B(n_1426), .C(n_1434), .Y(n_1424) );
OAI21xp5_ASAP7_75t_L g1771 ( .A1(n_607), .A2(n_1772), .B(n_1778), .Y(n_1771) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
AOI31xp33_ASAP7_75t_L g707 ( .A1(n_608), .A2(n_708), .A3(n_712), .B(n_716), .Y(n_707) );
AOI31xp33_ASAP7_75t_L g735 ( .A1(n_608), .A2(n_736), .A3(n_741), .B(n_744), .Y(n_735) );
AOI31xp33_ASAP7_75t_L g1077 ( .A1(n_608), .A2(n_1078), .A3(n_1081), .B(n_1084), .Y(n_1077) );
AOI31xp33_ASAP7_75t_SL g1121 ( .A1(n_608), .A2(n_1122), .A3(n_1125), .B(n_1127), .Y(n_1121) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_610), .B(n_620), .C(n_631), .D(n_642), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .C(n_616), .Y(n_610) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_SL g980 ( .A(n_615), .Y(n_980) );
INVx2_ASAP7_75t_L g1309 ( .A(n_615), .Y(n_1309) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_616), .B(n_756), .C(n_761), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_616), .B(n_819), .C(n_822), .Y(n_818) );
AOI33xp33_ASAP7_75t_L g884 ( .A1(n_616), .A2(n_630), .A3(n_885), .B1(n_887), .B2(n_888), .B3(n_892), .Y(n_884) );
AOI33xp33_ASAP7_75t_L g926 ( .A1(n_616), .A2(n_927), .A3(n_929), .B1(n_931), .B2(n_932), .B3(n_933), .Y(n_926) );
NAND3xp33_ASAP7_75t_L g1111 ( .A(n_616), .B(n_1112), .C(n_1115), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_616), .B(n_1166), .C(n_1169), .Y(n_1165) );
CKINVDCx8_ASAP7_75t_R g1463 ( .A(n_616), .Y(n_1463) );
INVx5_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx6_ASAP7_75t_L g690 ( .A(n_617), .Y(n_690) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .C(n_630), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g886 ( .A(n_623), .Y(n_886) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g762 ( .A(n_627), .Y(n_762) );
INVx1_ASAP7_75t_L g824 ( .A(n_627), .Y(n_824) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g930 ( .A(n_629), .Y(n_930) );
INVx2_ASAP7_75t_L g669 ( .A(n_630), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_630), .B(n_748), .C(n_752), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g974 ( .A(n_630), .B(n_975), .C(n_976), .Y(n_974) );
NAND3xp33_ASAP7_75t_L g1059 ( .A(n_630), .B(n_1060), .C(n_1062), .Y(n_1059) );
BUFx3_ASAP7_75t_L g1209 ( .A(n_630), .Y(n_1209) );
NAND3xp33_ASAP7_75t_L g1266 ( .A(n_630), .B(n_1267), .C(n_1268), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g1306 ( .A(n_630), .B(n_1307), .C(n_1308), .Y(n_1306) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .C(n_639), .Y(n_631) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx4_ASAP7_75t_L g698 ( .A(n_634), .Y(n_698) );
INVx1_ASAP7_75t_L g984 ( .A(n_634), .Y(n_984) );
INVx1_ASAP7_75t_L g1039 ( .A(n_634), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1157 ( .A(n_635), .Y(n_1157) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_639), .B(n_764), .C(n_770), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g982 ( .A(n_639), .B(n_983), .C(n_985), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g1068 ( .A(n_639), .B(n_1069), .C(n_1071), .Y(n_1068) );
NAND3xp33_ASAP7_75t_L g1274 ( .A(n_639), .B(n_1275), .C(n_1277), .Y(n_1274) );
NAND3xp33_ASAP7_75t_L g1313 ( .A(n_639), .B(n_1314), .C(n_1315), .Y(n_1313) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_SL g1347 ( .A1(n_640), .A2(n_1180), .B1(n_1348), .B2(n_1351), .Y(n_1347) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .C(n_645), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_645), .B(n_772), .C(n_774), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g986 ( .A(n_645), .B(n_987), .C(n_990), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g1072 ( .A(n_645), .B(n_1073), .C(n_1074), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1279 ( .A(n_645), .B(n_1280), .C(n_1281), .Y(n_1279) );
NAND3xp33_ASAP7_75t_L g1316 ( .A(n_645), .B(n_1317), .C(n_1318), .Y(n_1316) );
INVx1_ASAP7_75t_L g1393 ( .A(n_645), .Y(n_1393) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_719), .B1(n_720), .B2(n_778), .Y(n_647) );
INVx1_ASAP7_75t_L g778 ( .A(n_648), .Y(n_778) );
INVx1_ASAP7_75t_L g718 ( .A(n_650), .Y(n_718) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx4f_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_691), .Y(n_666) );
AOI33xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .A3(n_676), .B1(n_683), .B2(n_686), .B3(n_690), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_668), .B(n_813), .C(n_816), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g1160 ( .A(n_668), .B(n_1161), .C(n_1164), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_668), .A2(n_1445), .B1(n_1452), .B2(n_1462), .C(n_1464), .Y(n_1444) );
AOI33xp33_ASAP7_75t_L g1511 ( .A1(n_668), .A2(n_1462), .A3(n_1512), .B1(n_1513), .B2(n_1514), .B3(n_1515), .Y(n_1511) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g1170 ( .A(n_674), .Y(n_1170) );
INVx2_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_675), .Y(n_737) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
BUFx3_ASAP7_75t_L g685 ( .A(n_682), .Y(n_685) );
INVx2_ASAP7_75t_SL g815 ( .A(n_682), .Y(n_815) );
INVx4_ASAP7_75t_L g821 ( .A(n_682), .Y(n_821) );
INVx2_ASAP7_75t_SL g1168 ( .A(n_682), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1446 ( .A(n_684), .Y(n_1446) );
INVx1_ASAP7_75t_L g1458 ( .A(n_685), .Y(n_1458) );
AOI222xp33_ASAP7_75t_L g802 ( .A1(n_687), .A2(n_795), .B1(n_796), .B2(n_803), .C1(n_804), .C2(n_807), .Y(n_802) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g817 ( .A(n_688), .Y(n_817) );
INVx1_ASAP7_75t_L g867 ( .A(n_688), .Y(n_867) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g956 ( .A1(n_689), .A2(n_870), .B1(n_957), .B2(n_958), .C1(n_959), .C2(n_961), .Y(n_956) );
AOI33xp33_ASAP7_75t_L g1025 ( .A1(n_690), .A2(n_928), .A3(n_1026), .B1(n_1028), .B2(n_1029), .B3(n_1031), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1203 ( .A1(n_690), .A2(n_1204), .B1(n_1209), .B2(n_1210), .C(n_1216), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1779 ( .A1(n_690), .A2(n_1209), .B1(n_1780), .B2(n_1784), .C(n_1789), .Y(n_1779) );
AOI33xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .A3(n_697), .B1(n_699), .B2(n_702), .B3(n_706), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g1107 ( .A(n_692), .B(n_1108), .C(n_1109), .Y(n_1107) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g1177 ( .A(n_696), .Y(n_1177) );
BUFx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g1473 ( .A(n_701), .Y(n_1473) );
INVx1_ASAP7_75t_L g1470 ( .A(n_703), .Y(n_1470) );
BUFx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g1036 ( .A(n_704), .Y(n_1036) );
BUFx2_ASAP7_75t_L g1504 ( .A(n_704), .Y(n_1504) );
NAND3xp33_ASAP7_75t_L g834 ( .A(n_706), .B(n_835), .C(n_838), .Y(n_834) );
INVx5_ASAP7_75t_SL g1239 ( .A(n_714), .Y(n_1239) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g777 ( .A(n_722), .Y(n_777) );
BUFx2_ASAP7_75t_SL g1095 ( .A(n_732), .Y(n_1095) );
INVx1_ASAP7_75t_L g1188 ( .A(n_732), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1507 ( .A(n_732), .Y(n_1507) );
AOI222xp33_ASAP7_75t_L g1142 ( .A1(n_737), .A2(n_803), .B1(n_804), .B2(n_1143), .C1(n_1144), .C2(n_1145), .Y(n_1142) );
INVx1_ASAP7_75t_L g803 ( .A(n_740), .Y(n_803) );
NAND4xp25_ASAP7_75t_L g746 ( .A(n_747), .B(n_755), .C(n_763), .D(n_771), .Y(n_746) );
INVx2_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g935 ( .A(n_751), .Y(n_935) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx3_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g794 ( .A(n_769), .Y(n_794) );
AO22x2_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_896), .B1(n_897), .B2(n_994), .Y(n_779) );
INVx1_ASAP7_75t_L g994 ( .A(n_780), .Y(n_994) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_842), .Y(n_780) );
INVx1_ASAP7_75t_L g841 ( .A(n_782), .Y(n_841) );
NAND4xp25_ASAP7_75t_L g783 ( .A(n_784), .B(n_787), .C(n_790), .D(n_797), .Y(n_783) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND4xp25_ASAP7_75t_SL g1492 ( .A(n_797), .B(n_1493), .C(n_1495), .D(n_1497), .Y(n_1492) );
NAND4xp25_ASAP7_75t_SL g798 ( .A(n_799), .B(n_802), .C(n_808), .D(n_810), .Y(n_798) );
AOI222xp33_ASAP7_75t_L g865 ( .A1(n_803), .A2(n_866), .B1(n_867), .B2(n_868), .C1(n_869), .C2(n_870), .Y(n_865) );
AND2x4_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
AND2x4_ASAP7_75t_L g870 ( .A(n_805), .B(n_806), .Y(n_870) );
NAND4xp25_ASAP7_75t_SL g861 ( .A(n_810), .B(n_862), .C(n_865), .D(n_871), .Y(n_861) );
NAND4xp25_ASAP7_75t_L g952 ( .A(n_810), .B(n_953), .C(n_956), .D(n_962), .Y(n_952) );
NAND4xp25_ASAP7_75t_L g1138 ( .A(n_810), .B(n_1139), .C(n_1142), .D(n_1146), .Y(n_1138) );
NAND3xp33_ASAP7_75t_L g1228 ( .A(n_810), .B(n_1229), .C(n_1232), .Y(n_1228) );
NAND3xp33_ASAP7_75t_L g1426 ( .A(n_810), .B(n_1427), .C(n_1431), .Y(n_1426) );
NAND4xp25_ASAP7_75t_L g1481 ( .A(n_810), .B(n_1482), .C(n_1485), .D(n_1489), .Y(n_1481) );
NAND3xp33_ASAP7_75t_SL g1772 ( .A(n_810), .B(n_1773), .C(n_1775), .Y(n_1772) );
NAND4xp25_ASAP7_75t_L g811 ( .A(n_812), .B(n_818), .C(n_825), .D(n_834), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .C(n_833), .Y(n_825) );
INVx2_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
BUFx3_ASAP7_75t_L g1106 ( .A(n_830), .Y(n_1106) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g839 ( .A(n_832), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_832), .A2(n_1175), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1171 ( .A(n_833), .B(n_1172), .C(n_1173), .Y(n_1171) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g1535 ( .A1(n_840), .A2(n_1536), .B1(n_1537), .B2(n_1543), .Y(n_1535) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_855), .C(n_858), .Y(n_845) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1295 ( .A(n_849), .Y(n_1295) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_884), .Y(n_874) );
HB1xp67_ASAP7_75t_L g1506 ( .A(n_877), .Y(n_1506) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g1037 ( .A(n_880), .Y(n_1037) );
INVx1_ASAP7_75t_L g1360 ( .A(n_880), .Y(n_1360) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g1119 ( .A(n_891), .Y(n_1119) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1027 ( .A(n_894), .Y(n_1027) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_949), .B1(n_950), .B2(n_993), .Y(n_897) );
INVx1_ASAP7_75t_L g993 ( .A(n_898), .Y(n_993) );
INVx1_ASAP7_75t_L g948 ( .A(n_899), .Y(n_948) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AOI31xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_916), .A3(n_921), .B(n_924), .Y(n_913) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
AO21x1_ASAP7_75t_SL g1018 ( .A1(n_924), .A2(n_1019), .B(n_1022), .Y(n_1018) );
AOI31xp33_ASAP7_75t_L g1256 ( .A1(n_924), .A2(n_1257), .A3(n_1260), .B(n_1263), .Y(n_1256) );
AOI31xp33_ASAP7_75t_L g1296 ( .A1(n_924), .A2(n_1297), .A3(n_1300), .B(n_1303), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_936), .Y(n_925) );
BUFx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
NAND3xp33_ASAP7_75t_L g1116 ( .A(n_928), .B(n_1117), .C(n_1120), .Y(n_1116) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g1110 ( .A(n_939), .Y(n_1110) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx2_ASAP7_75t_SL g1278 ( .A(n_946), .Y(n_1278) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g992 ( .A(n_951), .Y(n_992) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_966), .B(n_968), .C(n_970), .Y(n_965) );
NAND4xp25_ASAP7_75t_L g973 ( .A(n_974), .B(n_977), .C(n_982), .D(n_986), .Y(n_973) );
NAND3xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .C(n_981), .Y(n_977) );
NAND3xp33_ASAP7_75t_L g1063 ( .A(n_981), .B(n_1064), .C(n_1066), .Y(n_1063) );
NAND3xp33_ASAP7_75t_L g1269 ( .A(n_981), .B(n_1270), .C(n_1273), .Y(n_1269) );
NAND3xp33_ASAP7_75t_L g1310 ( .A(n_981), .B(n_1311), .C(n_1312), .Y(n_1310) );
INVx1_ASAP7_75t_L g1346 ( .A(n_981), .Y(n_1346) );
BUFx2_ASAP7_75t_L g1510 ( .A(n_988), .Y(n_1510) );
INVx2_ASAP7_75t_SL g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1070 ( .A(n_989), .Y(n_1070) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B1(n_1087), .B2(n_1130), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
AO22x2_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1043), .B1(n_1044), .B2(n_1086), .Y(n_998) );
INVx1_ASAP7_75t_L g1086 ( .A(n_999), .Y(n_1086) );
NAND4xp25_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1018), .C(n_1025), .D(n_1033), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1011), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1348 ( .A1(n_1005), .A2(n_1328), .B1(n_1331), .B2(n_1349), .C(n_1350), .Y(n_1348) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
AOI211xp5_ASAP7_75t_L g1045 ( .A1(n_1046), .A2(n_1047), .B(n_1058), .C(n_1077), .Y(n_1045) );
OAI31xp33_ASAP7_75t_L g1192 ( .A1(n_1046), .A2(n_1193), .A3(n_1195), .B(n_1201), .Y(n_1192) );
AOI211xp5_ASAP7_75t_L g1245 ( .A1(n_1046), .A2(n_1246), .B(n_1256), .C(n_1265), .Y(n_1245) );
AOI211xp5_ASAP7_75t_L g1284 ( .A1(n_1046), .A2(n_1285), .B(n_1296), .C(n_1305), .Y(n_1284) );
OAI31xp33_ASAP7_75t_SL g1356 ( .A1(n_1046), .A2(n_1357), .A3(n_1358), .B(n_1363), .Y(n_1356) );
OAI31xp33_ASAP7_75t_L g1406 ( .A1(n_1046), .A2(n_1407), .A3(n_1408), .B(n_1409), .Y(n_1406) );
OAI31xp33_ASAP7_75t_SL g1764 ( .A1(n_1046), .A2(n_1765), .A3(n_1766), .B(n_1767), .Y(n_1764) );
NAND4xp25_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1063), .C(n_1068), .D(n_1072), .Y(n_1058) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1087), .Y(n_1130) );
NOR3xp33_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1102), .C(n_1121), .Y(n_1088) );
AOI31xp33_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1093), .A3(n_1098), .B(n_1101), .Y(n_1089) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1101), .Y(n_1158) );
NAND4xp25_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1107), .C(n_1111), .D(n_1116), .Y(n_1102) );
BUFx3_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1114), .Y(n_1163) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1114), .Y(n_1340) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
XOR2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1420), .Y(n_1132) );
XNOR2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1240), .Y(n_1133) );
XNOR2x2_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1189), .Y(n_1134) );
XNOR2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1578 ( .A1(n_1136), .A2(n_1539), .B1(n_1546), .B2(n_1579), .Y(n_1578) );
NAND4xp25_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1165), .C(n_1171), .D(n_1178), .Y(n_1159) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVxp67_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
BUFx3_ASAP7_75t_L g1467 ( .A(n_1176), .Y(n_1467) );
NAND3xp33_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1181), .C(n_1186), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
OAI22xp5_ASAP7_75t_SL g1216 ( .A1(n_1180), .A2(n_1217), .B1(n_1218), .B2(n_1222), .Y(n_1216) );
OAI22xp5_ASAP7_75t_SL g1789 ( .A1(n_1180), .A2(n_1217), .B1(n_1790), .B2(n_1792), .Y(n_1789) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
XNOR2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1191), .Y(n_1189) );
NAND3x1_ASAP7_75t_SL g1191 ( .A(n_1192), .B(n_1203), .C(n_1227), .Y(n_1191) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1250 ( .A1(n_1197), .A2(n_1251), .B(n_1252), .Y(n_1250) );
AOI21xp5_ASAP7_75t_L g1292 ( .A1(n_1197), .A2(n_1293), .B(n_1294), .Y(n_1292) );
OAI221xp5_ASAP7_75t_L g1218 ( .A1(n_1206), .A2(n_1208), .B1(n_1219), .B2(n_1220), .C(n_1221), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g1342 ( .A1(n_1207), .A2(n_1343), .B1(n_1344), .B2(n_1345), .Y(n_1342) );
OAI22xp5_ASAP7_75t_SL g1447 ( .A1(n_1213), .A2(n_1448), .B1(n_1449), .B2(n_1450), .Y(n_1447) );
OAI22xp5_ASAP7_75t_L g1781 ( .A1(n_1213), .A2(n_1450), .B1(n_1782), .B2(n_1783), .Y(n_1781) );
INVx3_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
OAI33xp33_ASAP7_75t_L g1374 ( .A1(n_1217), .A2(n_1375), .A3(n_1380), .B1(n_1387), .B2(n_1390), .B3(n_1393), .Y(n_1374) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_1219), .A2(n_1220), .B1(n_1223), .B2(n_1224), .C(n_1225), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g1465 ( .A1(n_1220), .A2(n_1352), .B1(n_1448), .B2(n_1449), .C(n_1466), .Y(n_1465) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_1220), .A2(n_1429), .B1(n_1470), .B2(n_1471), .C(n_1472), .Y(n_1469) );
OAI221xp5_ASAP7_75t_L g1790 ( .A1(n_1220), .A2(n_1352), .B1(n_1787), .B2(n_1788), .C(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1226), .Y(n_1379) );
BUFx6f_ASAP7_75t_L g1468 ( .A(n_1226), .Y(n_1468) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1226), .Y(n_1475) );
BUFx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
BUFx2_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1238), .Y(n_1335) );
XOR2x2_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1319), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1243), .B1(n_1282), .B2(n_1283), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
XNOR2xp5_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1245), .Y(n_1243) );
NAND4xp25_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1269), .C(n_1274), .D(n_1279), .Y(n_1265) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
NAND4xp25_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1310), .C(n_1313), .D(n_1316), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1371), .B1(n_1418), .B2(n_1419), .Y(n_1319) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1320), .Y(n_1418) );
NAND3xp33_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1356), .C(n_1364), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1347), .Y(n_1322) );
OAI33xp33_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1326), .A3(n_1332), .B1(n_1338), .B2(n_1342), .B3(n_1346), .Y(n_1323) );
OAI33xp33_ASAP7_75t_L g1394 ( .A1(n_1324), .A2(n_1346), .A3(n_1395), .B1(n_1398), .B2(n_1399), .B3(n_1403), .Y(n_1394) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1328), .B1(n_1329), .B2(n_1331), .Y(n_1326) );
OAI22xp33_ASAP7_75t_L g1395 ( .A1(n_1329), .A2(n_1381), .B1(n_1384), .B2(n_1396), .Y(n_1395) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1329), .Y(n_1451) );
BUFx3_ASAP7_75t_L g1461 ( .A(n_1329), .Y(n_1461) );
BUFx6f_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
OAI22xp33_ASAP7_75t_SL g1332 ( .A1(n_1333), .A2(n_1334), .B1(n_1336), .B2(n_1337), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_1334), .A2(n_1339), .B1(n_1340), .B2(n_1341), .Y(n_1338) );
OAI22xp33_ASAP7_75t_L g1398 ( .A1(n_1334), .A2(n_1340), .B1(n_1376), .B2(n_1378), .Y(n_1398) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1335), .Y(n_1400) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1337), .Y(n_1785) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_1340), .A2(n_1400), .B1(n_1401), .B2(n_1402), .Y(n_1399) );
OAI221xp5_ASAP7_75t_L g1792 ( .A1(n_1352), .A2(n_1774), .B1(n_1776), .B2(n_1793), .C(n_1794), .Y(n_1792) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1371), .Y(n_1419) );
NAND3xp33_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1406), .C(n_1413), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1394), .Y(n_1373) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_1376), .A2(n_1377), .B1(n_1378), .B2(n_1379), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1382), .B1(n_1384), .B2(n_1385), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_1382), .A2(n_1385), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1386), .Y(n_1793) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1477), .B1(n_1478), .B2(n_1517), .Y(n_1420) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1421), .Y(n_1517) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1444), .Y(n_1423) );
AOI21xp5_ASAP7_75t_L g1434 ( .A1(n_1435), .A2(n_1440), .B(n_1443), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx2_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1442), .Y(n_1440) );
INVx2_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
OAI22xp33_ASAP7_75t_SL g1456 ( .A1(n_1457), .A2(n_1458), .B1(n_1459), .B2(n_1460), .Y(n_1456) );
BUFx3_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx2_ASAP7_75t_SL g1477 ( .A(n_1478), .Y(n_1477) );
OAI22xp33_ASAP7_75t_L g1583 ( .A1(n_1479), .A2(n_1538), .B1(n_1544), .B2(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1480), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1511), .Y(n_1501) );
OAI221xp5_ASAP7_75t_R g1518 ( .A1(n_1519), .A2(n_1760), .B1(n_1761), .B2(n_1795), .C(n_1800), .Y(n_1518) );
AND4x1_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1687), .C(n_1701), .D(n_1733), .Y(n_1519) );
AOI211xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1548), .B(n_1649), .C(n_1663), .Y(n_1520) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1521), .B(n_1665), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1521), .B(n_1622), .Y(n_1710) );
AOI221xp5_ASAP7_75t_L g1728 ( .A1(n_1521), .A2(n_1598), .B1(n_1626), .B2(n_1729), .C(n_1730), .Y(n_1728) );
OAI333xp33_ASAP7_75t_L g1752 ( .A1(n_1521), .A2(n_1596), .A3(n_1654), .B1(n_1689), .B2(n_1753), .B3(n_1755), .C1(n_1756), .C2(n_1758), .C3(n_1759), .Y(n_1752) );
CKINVDCx5p33_ASAP7_75t_R g1521 ( .A(n_1522), .Y(n_1521) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1522), .B(n_1656), .Y(n_1689) );
OAI32xp33_ASAP7_75t_L g1709 ( .A1(n_1522), .A2(n_1562), .A3(n_1622), .B1(n_1681), .B2(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1522), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1522), .B(n_1581), .Y(n_1758) );
OR2x6_ASAP7_75t_SL g1522 ( .A(n_1523), .B(n_1535), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_1524), .A2(n_1525), .B1(n_1532), .B2(n_1533), .Y(n_1523) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1526), .Y(n_1587) );
AND2x4_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1530), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1527), .B(n_1530), .Y(n_1555) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
AND2x4_ASAP7_75t_L g1534 ( .A(n_1528), .B(n_1530), .Y(n_1534) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1529), .B(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1531), .Y(n_1542) );
INVx2_ASAP7_75t_L g1572 ( .A(n_1533), .Y(n_1572) );
INVx2_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_SL g1557 ( .A(n_1534), .Y(n_1557) );
BUFx3_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
OAI22xp5_ASAP7_75t_L g1559 ( .A1(n_1538), .A2(n_1546), .B1(n_1560), .B2(n_1561), .Y(n_1559) );
OAI22xp33_ASAP7_75t_L g1600 ( .A1(n_1538), .A2(n_1546), .B1(n_1601), .B2(n_1602), .Y(n_1600) );
BUFx6f_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
OR2x2_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1541), .Y(n_1539) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1540), .B(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1540), .Y(n_1568) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1541), .Y(n_1567) );
BUFx2_ASAP7_75t_SL g1760 ( .A(n_1543), .Y(n_1760) );
HB1xp67_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1547), .Y(n_1570) );
NAND5xp2_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1617), .C(n_1630), .D(n_1638), .E(n_1642), .Y(n_1548) );
AOI211xp5_ASAP7_75t_SL g1549 ( .A1(n_1550), .A2(n_1580), .B(n_1592), .C(n_1613), .Y(n_1549) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1550), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1562), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1551), .B(n_1595), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1551), .B(n_1596), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1551), .B(n_1564), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1641 ( .A(n_1551), .B(n_1564), .Y(n_1641) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1551), .B(n_1673), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1551), .B(n_1607), .Y(n_1684) );
OR2x2_ASAP7_75t_L g1686 ( .A(n_1551), .B(n_1607), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1551), .B(n_1606), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1551), .B(n_1573), .Y(n_1713) );
NOR2xp33_ASAP7_75t_L g1724 ( .A(n_1551), .B(n_1624), .Y(n_1724) );
NOR2xp33_ASAP7_75t_L g1754 ( .A(n_1551), .B(n_1577), .Y(n_1754) );
CKINVDCx6p67_ASAP7_75t_R g1551 ( .A(n_1552), .Y(n_1551) );
OR2x2_ASAP7_75t_L g1644 ( .A(n_1552), .B(n_1596), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1552), .B(n_1631), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1552), .B(n_1596), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1552), .B(n_1573), .Y(n_1681) );
NAND2xp5_ASAP7_75t_L g1693 ( .A(n_1552), .B(n_1694), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1552), .B(n_1595), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1552), .B(n_1606), .Y(n_1727) );
OR2x2_ASAP7_75t_L g1736 ( .A(n_1552), .B(n_1632), .Y(n_1736) );
OR2x6_ASAP7_75t_SL g1552 ( .A(n_1553), .B(n_1559), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_1554), .A2(n_1556), .B1(n_1557), .B2(n_1558), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g1585 ( .A1(n_1557), .A2(n_1586), .B1(n_1587), .B2(n_1588), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1573), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1593 ( .A(n_1563), .B(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1563), .Y(n_1605) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1563), .B(n_1658), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1694 ( .A(n_1563), .B(n_1632), .Y(n_1694) );
INVx4_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1564), .B(n_1612), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1564), .B(n_1573), .Y(n_1624) );
INVx2_ASAP7_75t_L g1636 ( .A(n_1564), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1564), .B(n_1582), .Y(n_1673) );
OR2x2_ASAP7_75t_L g1720 ( .A(n_1564), .B(n_1647), .Y(n_1720) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1564), .B(n_1727), .Y(n_1726) );
OR2x2_ASAP7_75t_L g1731 ( .A(n_1564), .B(n_1632), .Y(n_1731) );
OR2x2_ASAP7_75t_L g1735 ( .A(n_1564), .B(n_1736), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1564), .B(n_1648), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1564), .B(n_1626), .Y(n_1757) );
AND2x6_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1571), .Y(n_1564) );
AND2x4_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1568), .Y(n_1566) );
AND2x4_ASAP7_75t_L g1569 ( .A(n_1568), .B(n_1570), .Y(n_1569) );
HB1xp67_ASAP7_75t_L g1810 ( .A(n_1570), .Y(n_1810) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1577), .Y(n_1573) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1574), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1574), .B(n_1607), .Y(n_1606) );
OR2x2_ASAP7_75t_L g1632 ( .A(n_1574), .B(n_1577), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1576), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1577), .B(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1577), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_1580), .B(n_1662), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1580), .B(n_1729), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1589), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1581), .B(n_1598), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1581), .B(n_1610), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1581), .B(n_1622), .Y(n_1621) );
OR2x2_ASAP7_75t_L g1654 ( .A(n_1581), .B(n_1589), .Y(n_1654) );
INVx3_ASAP7_75t_L g1656 ( .A(n_1581), .Y(n_1656) );
AOI21xp5_ASAP7_75t_L g1748 ( .A1(n_1581), .A2(n_1749), .B(n_1752), .Y(n_1748) );
INVx3_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1615 ( .A(n_1582), .B(n_1616), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1582), .B(n_1589), .Y(n_1747) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1585), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1589), .B(n_1599), .Y(n_1598) );
OR2x2_ASAP7_75t_L g1616 ( .A(n_1589), .B(n_1599), .Y(n_1616) );
INVx2_ASAP7_75t_L g1622 ( .A(n_1589), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1589), .B(n_1610), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1589), .B(n_1610), .Y(n_1637) );
AOI22xp5_ASAP7_75t_L g1690 ( .A1(n_1589), .A2(n_1658), .B1(n_1691), .B2(n_1695), .Y(n_1690) );
OAI221xp5_ASAP7_75t_L g1717 ( .A1(n_1589), .A2(n_1716), .B1(n_1718), .B2(n_1726), .C(n_1728), .Y(n_1717) );
AND2x4_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1591), .Y(n_1589) );
OAI21xp5_ASAP7_75t_SL g1592 ( .A1(n_1593), .A2(n_1597), .B(n_1603), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1655 ( .A(n_1594), .B(n_1656), .Y(n_1655) );
A2O1A1Ixp33_ASAP7_75t_SL g1687 ( .A1(n_1594), .A2(n_1688), .B(n_1690), .C(n_1698), .Y(n_1687) );
AOI211xp5_ASAP7_75t_L g1718 ( .A1(n_1594), .A2(n_1719), .B(n_1721), .C(n_1725), .Y(n_1718) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1595), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1595), .B(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
AOI322xp5_ASAP7_75t_L g1668 ( .A1(n_1598), .A2(n_1621), .A3(n_1669), .B1(n_1671), .B2(n_1674), .C1(n_1677), .C2(n_1682), .Y(n_1668) );
INVx2_ASAP7_75t_SL g1610 ( .A(n_1599), .Y(n_1610) );
HB1xp67_ASAP7_75t_L g1620 ( .A(n_1599), .Y(n_1620) );
AOI22xp5_ASAP7_75t_L g1603 ( .A1(n_1604), .A2(n_1608), .B1(n_1609), .B2(n_1611), .Y(n_1603) );
INVxp67_ASAP7_75t_L g1759 ( .A(n_1604), .Y(n_1759) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1606), .Y(n_1670) );
NOR2xp33_ASAP7_75t_L g1753 ( .A(n_1606), .B(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1609), .Y(n_1737) );
INVx2_ASAP7_75t_SL g1648 ( .A(n_1610), .Y(n_1648) );
NOR2xp33_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1615), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1614), .B(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1615), .Y(n_1682) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1616), .Y(n_1700) );
OAI21xp33_ASAP7_75t_SL g1711 ( .A1(n_1616), .A2(n_1712), .B(n_1714), .Y(n_1711) );
AOI21xp5_ASAP7_75t_L g1617 ( .A1(n_1618), .A2(n_1623), .B(n_1625), .Y(n_1617) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1620), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1666 ( .A(n_1620), .B(n_1667), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1620), .B(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1620), .Y(n_1716) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1620), .Y(n_1723) );
AOI211xp5_ASAP7_75t_SL g1738 ( .A1(n_1621), .A2(n_1739), .B(n_1740), .C(n_1741), .Y(n_1738) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
A2O1A1Ixp33_ASAP7_75t_L g1734 ( .A1(n_1624), .A2(n_1735), .B(n_1737), .C(n_1738), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1627), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1638 ( .A(n_1626), .B(n_1639), .Y(n_1638) );
AOI21xp5_ASAP7_75t_L g1698 ( .A1(n_1626), .A2(n_1699), .B(n_1700), .Y(n_1698) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1626), .Y(n_1704) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
NOR2xp33_ASAP7_75t_L g1660 ( .A(n_1628), .B(n_1661), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1629), .B(n_1631), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1633), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1631), .B(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
OAI211xp5_ASAP7_75t_L g1683 ( .A1(n_1633), .A2(n_1656), .B(n_1684), .C(n_1685), .Y(n_1683) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
OR2x2_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1637), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1635), .B(n_1679), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1635), .B(n_1697), .Y(n_1696) );
NOR2x1_ASAP7_75t_L g1729 ( .A(n_1635), .B(n_1686), .Y(n_1729) );
INVx2_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1646 ( .A(n_1636), .B(n_1647), .Y(n_1646) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1636), .B(n_1643), .Y(n_1739) );
INVx2_ASAP7_75t_L g1658 ( .A(n_1637), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1639), .B(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
NOR2xp33_ASAP7_75t_L g1751 ( .A(n_1640), .B(n_1716), .Y(n_1751) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1641), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1645), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1648), .Y(n_1662) );
OAI21xp33_ASAP7_75t_L g1749 ( .A1(n_1648), .A2(n_1675), .B(n_1750), .Y(n_1749) );
OAI221xp5_ASAP7_75t_L g1649 ( .A1(n_1650), .A2(n_1654), .B1(n_1655), .B2(n_1657), .C(n_1659), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1652), .Y(n_1650) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_SL g1665 ( .A(n_1656), .Y(n_1665) );
NOR3xp33_ASAP7_75t_L g1741 ( .A(n_1656), .B(n_1670), .C(n_1720), .Y(n_1741) );
INVxp67_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
NOR2xp33_ASAP7_75t_L g1692 ( .A(n_1662), .B(n_1693), .Y(n_1692) );
OAI211xp5_ASAP7_75t_SL g1663 ( .A1(n_1664), .A2(n_1666), .B(n_1668), .C(n_1683), .Y(n_1663) );
OAI311xp33_ASAP7_75t_L g1701 ( .A1(n_1664), .A2(n_1702), .A3(n_1703), .B1(n_1711), .C1(n_1717), .Y(n_1701) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1667), .Y(n_1706) );
OR2x2_ASAP7_75t_L g1675 ( .A(n_1670), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
NAND2xp33_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1680), .Y(n_1677) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1693), .Y(n_1725) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1695), .Y(n_1702) );
INVxp67_ASAP7_75t_L g1745 ( .A(n_1696), .Y(n_1745) );
OAI21xp33_ASAP7_75t_L g1703 ( .A1(n_1704), .A2(n_1705), .B(n_1709), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1707), .Y(n_1705) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
A2O1A1Ixp33_ASAP7_75t_L g1744 ( .A1(n_1714), .A2(n_1745), .B(n_1746), .C(n_1748), .Y(n_1744) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1724), .Y(n_1722) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1727), .Y(n_1732) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1731), .B(n_1732), .Y(n_1730) );
AOI21xp5_ASAP7_75t_L g1733 ( .A1(n_1734), .A2(n_1742), .B(n_1744), .Y(n_1733) );
CKINVDCx14_ASAP7_75t_R g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
INVxp33_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1763), .Y(n_1808) );
NAND3x1_ASAP7_75t_L g1763 ( .A(n_1764), .B(n_1771), .C(n_1779), .Y(n_1763) );
CKINVDCx5p33_ASAP7_75t_R g1795 ( .A(n_1796), .Y(n_1795) );
BUFx2_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1799), .Y(n_1798) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
CKINVDCx5p33_ASAP7_75t_R g1802 ( .A(n_1803), .Y(n_1802) );
OAI21xp5_ASAP7_75t_L g1809 ( .A1(n_1804), .A2(n_1810), .B(n_1811), .Y(n_1809) );
INVxp33_ASAP7_75t_SL g1805 ( .A(n_1806), .Y(n_1805) );
endmodule