module fake_jpeg_21153_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_29),
.C(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_42),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_31),
.B1(n_20),
.B2(n_28),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_55),
.B1(n_24),
.B2(n_21),
.Y(n_74)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_52),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_60),
.Y(n_89)
);

BUFx2_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_39),
.B1(n_37),
.B2(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_23),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_35),
.B(n_21),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_76),
.B(n_77),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_39),
.B1(n_41),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_18),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_83),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_24),
.B1(n_29),
.B2(n_25),
.Y(n_75)
);

AND2x4_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_41),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_41),
.B1(n_19),
.B2(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_41),
.C(n_22),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_23),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_59),
.B1(n_57),
.B2(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_23),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_56),
.B1(n_24),
.B2(n_60),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_66),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_23),
.B(n_19),
.C(n_26),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_115),
.B1(n_117),
.B2(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_22),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_91),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_110),
.B1(n_106),
.B2(n_103),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_137),
.B1(n_140),
.B2(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_125),
.B1(n_136),
.B2(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_132),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_84),
.B1(n_67),
.B2(n_69),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_130),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_89),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_133),
.B(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_82),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_84),
.C(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_86),
.B1(n_68),
.B2(n_63),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_19),
.Y(n_167)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_63),
.B1(n_71),
.B2(n_88),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_22),
.C(n_19),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_143),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_93),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_95),
.B1(n_98),
.B2(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_156),
.B1(n_162),
.B2(n_169),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_123),
.Y(n_173)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_168),
.B1(n_170),
.B2(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_116),
.B1(n_87),
.B2(n_85),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_168)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_30),
.B1(n_18),
.B2(n_26),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_30),
.B1(n_18),
.B2(n_3),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_129),
.B(n_133),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_169),
.B1(n_8),
.B2(n_9),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_179),
.CI(n_158),
.CON(n_192),
.SN(n_192)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_142),
.B(n_30),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_0),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_181),
.C(n_159),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_185),
.Y(n_194)
);

XOR2x2_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_3),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_152),
.C(n_154),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_5),
.B(n_7),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_5),
.B(n_7),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_13),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_204),
.C(n_176),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_161),
.C(n_152),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_210)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_147),
.C(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_191),
.C(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_157),
.C(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_171),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_169),
.B1(n_8),
.B2(n_10),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_169),
.B1(n_15),
.B2(n_14),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_187),
.B(n_182),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_194),
.B(n_192),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_203),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_216),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_190),
.B(n_179),
.C(n_178),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_219),
.B(n_205),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_189),
.B(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_220),
.C(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_208),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_171),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_201),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_14),
.CI(n_8),
.CON(n_231),
.SN(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_222),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_193),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_228),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_230),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_192),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_224),
.B(n_229),
.C(n_230),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_215),
.B1(n_212),
.B2(n_11),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_215),
.C(n_10),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_215),
.C(n_11),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_231),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_242),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_7),
.B(n_12),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_12),
.B(n_239),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_235),
.B(n_232),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_245),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_248),
.B(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_234),
.C(n_12),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_250),
.C(n_253),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_255),
.Y(n_256)
);


endmodule