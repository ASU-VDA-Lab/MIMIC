module real_aes_1830_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g226 ( .A(n_0), .B(n_141), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_1), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g132 ( .A(n_2), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_3), .B(n_125), .Y(n_124) );
NAND2xp33_ASAP7_75t_SL g211 ( .A(n_4), .B(n_131), .Y(n_211) );
INVx1_ASAP7_75t_L g202 ( .A(n_5), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_6), .B(n_145), .Y(n_476) );
INVx1_ASAP7_75t_L g519 ( .A(n_7), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g806 ( .A(n_8), .Y(n_806) );
AND2x2_ASAP7_75t_L g119 ( .A(n_9), .B(n_120), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_10), .Y(n_533) );
INVx2_ASAP7_75t_L g121 ( .A(n_11), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_12), .Y(n_426) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_12), .B(n_805), .C(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g484 ( .A(n_13), .Y(n_484) );
AOI221x1_ASAP7_75t_L g205 ( .A1(n_14), .A2(n_134), .B1(n_206), .B2(n_208), .C(n_210), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_15), .B(n_125), .Y(n_192) );
INVx1_ASAP7_75t_L g430 ( .A(n_16), .Y(n_430) );
NOR2xp33_ASAP7_75t_SL g802 ( .A(n_16), .B(n_431), .Y(n_802) );
INVx1_ASAP7_75t_L g482 ( .A(n_17), .Y(n_482) );
INVx1_ASAP7_75t_SL g469 ( .A(n_18), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_19), .B(n_126), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_20), .A2(n_134), .B(n_139), .Y(n_133) );
AOI221xp5_ASAP7_75t_SL g216 ( .A1(n_21), .A2(n_38), .B1(n_125), .B2(n_134), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_22), .B(n_141), .Y(n_140) );
AOI33xp33_ASAP7_75t_L g499 ( .A1(n_23), .A2(n_52), .A3(n_178), .B1(n_185), .B2(n_500), .B3(n_501), .Y(n_499) );
AOI22x1_ASAP7_75t_R g757 ( .A1(n_24), .A2(n_36), .B1(n_758), .B2(n_759), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_24), .Y(n_759) );
INVx1_ASAP7_75t_L g527 ( .A(n_25), .Y(n_527) );
OR2x2_ASAP7_75t_L g122 ( .A(n_26), .B(n_93), .Y(n_122) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_26), .A2(n_93), .B(n_121), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_27), .B(n_143), .Y(n_196) );
INVxp67_ASAP7_75t_L g204 ( .A(n_28), .Y(n_204) );
AND2x2_ASAP7_75t_L g165 ( .A(n_29), .B(n_155), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g780 ( .A1(n_29), .A2(n_90), .B1(n_781), .B2(n_782), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_29), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_30), .B(n_176), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_31), .A2(n_134), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_32), .B(n_143), .Y(n_218) );
AND2x2_ASAP7_75t_L g131 ( .A(n_33), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g135 ( .A(n_33), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g184 ( .A(n_33), .Y(n_184) );
OR2x6_ASAP7_75t_L g428 ( .A(n_34), .B(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g807 ( .A(n_34), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_35), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_36), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_37), .B(n_176), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_39), .A2(n_145), .B1(n_209), .B2(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_40), .B(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_41), .A2(n_83), .B1(n_134), .B2(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_42), .B(n_126), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_43), .B(n_141), .Y(n_163) );
XOR2xp5_ASAP7_75t_L g433 ( .A(n_44), .B(n_434), .Y(n_433) );
AOI22x1_ASAP7_75t_SL g788 ( .A1(n_44), .A2(n_68), .B1(n_789), .B2(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_44), .Y(n_789) );
XNOR2x2_ASAP7_75t_SL g756 ( .A(n_45), .B(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_46), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_47), .B(n_172), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_48), .B(n_126), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_49), .Y(n_446) );
AND2x2_ASAP7_75t_L g229 ( .A(n_50), .B(n_155), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_51), .B(n_155), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_53), .B(n_126), .Y(n_511) );
INVxp33_ASAP7_75t_L g809 ( .A(n_54), .Y(n_809) );
INVx1_ASAP7_75t_L g128 ( .A(n_55), .Y(n_128) );
INVx1_ASAP7_75t_L g138 ( .A(n_55), .Y(n_138) );
AND2x2_ASAP7_75t_L g512 ( .A(n_56), .B(n_155), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_57), .A2(n_75), .B1(n_176), .B2(n_182), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_58), .B(n_176), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_59), .B(n_125), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_60), .B(n_209), .Y(n_535) );
AOI21xp5_ASAP7_75t_SL g456 ( .A1(n_61), .A2(n_182), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g156 ( .A(n_62), .B(n_155), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_63), .B(n_143), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_64), .B(n_141), .Y(n_152) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_65), .B(n_120), .Y(n_197) );
INVx1_ASAP7_75t_L g479 ( .A(n_66), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_67), .A2(n_134), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_68), .Y(n_790) );
INVx1_ASAP7_75t_L g510 ( .A(n_69), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_70), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_71), .B(n_172), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_72), .A2(n_182), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g130 ( .A(n_73), .Y(n_130) );
INVx1_ASAP7_75t_L g136 ( .A(n_73), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_74), .B(n_176), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_76), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g471 ( .A(n_77), .B(n_208), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_78), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_79), .A2(n_182), .B(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_80), .A2(n_171), .B(n_182), .C(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_81), .B(n_125), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_82), .A2(n_86), .B1(n_125), .B2(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g431 ( .A(n_84), .Y(n_431) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_85), .B(n_208), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_87), .A2(n_182), .B1(n_497), .B2(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_88), .B(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_89), .B(n_141), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_90), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g755 ( .A(n_91), .B(n_756), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_92), .A2(n_134), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g458 ( .A(n_94), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_95), .B(n_143), .Y(n_151) );
AND2x2_ASAP7_75t_L g503 ( .A(n_96), .B(n_208), .Y(n_503) );
OAI22xp33_ASAP7_75t_SL g786 ( .A1(n_97), .A2(n_787), .B1(n_788), .B2(n_791), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_97), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_98), .A2(n_525), .B(n_526), .C(n_528), .Y(n_524) );
INVxp67_ASAP7_75t_L g207 ( .A(n_99), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_100), .B(n_125), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_101), .B(n_143), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_102), .A2(n_134), .B(n_194), .Y(n_193) );
BUFx2_ASAP7_75t_L g771 ( .A(n_103), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_104), .B(n_126), .Y(n_459) );
AOI21xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_796), .B(n_808), .Y(n_105) );
OA22x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_767), .B1(n_776), .B2(n_794), .Y(n_106) );
OAI21xp5_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_755), .B(n_760), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OAI22x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_423), .B1(n_432), .B2(n_753), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g762 ( .A(n_111), .Y(n_762) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_345), .Y(n_111) );
NOR3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_269), .C(n_319), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_249), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_188), .B(n_230), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_166), .Y(n_116) );
INVx1_ASAP7_75t_SL g355 ( .A(n_117), .Y(n_355) );
AOI32xp33_ASAP7_75t_L g386 ( .A1(n_117), .A2(n_368), .A3(n_387), .B1(n_388), .B2(n_389), .Y(n_386) );
AND2x2_ASAP7_75t_L g388 ( .A(n_117), .B(n_245), .Y(n_388) );
AND2x4_ASAP7_75t_SL g117 ( .A(n_118), .B(n_146), .Y(n_117) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
INVx5_ASAP7_75t_L g248 ( .A(n_118), .Y(n_248) );
OR2x2_ASAP7_75t_L g255 ( .A(n_118), .B(n_247), .Y(n_255) );
INVx2_ASAP7_75t_L g260 ( .A(n_118), .Y(n_260) );
AND2x2_ASAP7_75t_L g272 ( .A(n_118), .B(n_147), .Y(n_272) );
AND2x2_ASAP7_75t_L g277 ( .A(n_118), .B(n_157), .Y(n_277) );
OR2x2_ASAP7_75t_L g284 ( .A(n_118), .B(n_169), .Y(n_284) );
AND2x4_ASAP7_75t_L g293 ( .A(n_118), .B(n_158), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_SL g335 ( .A1(n_118), .A2(n_251), .B(n_286), .C(n_324), .Y(n_335) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
AND2x2_ASAP7_75t_SL g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x4_ASAP7_75t_L g145 ( .A(n_121), .B(n_122), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_133), .B(n_145), .Y(n_123) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
INVx1_ASAP7_75t_L g212 ( .A(n_126), .Y(n_212) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
AND2x6_ASAP7_75t_L g141 ( .A(n_127), .B(n_136), .Y(n_141) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g143 ( .A(n_129), .B(n_138), .Y(n_143) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx5_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_131), .Y(n_528) );
AND2x2_ASAP7_75t_L g137 ( .A(n_132), .B(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
BUFx3_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
INVx2_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
AND2x4_ASAP7_75t_L g182 ( .A(n_137), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_142), .B(n_144), .Y(n_139) );
INVxp67_ASAP7_75t_L g483 ( .A(n_141), .Y(n_483) );
INVxp67_ASAP7_75t_L g485 ( .A(n_143), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_144), .A2(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_144), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_144), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_144), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_144), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_144), .A2(n_449), .B(n_450), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_144), .A2(n_452), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g468 ( .A1(n_144), .A2(n_452), .B(n_469), .C(n_470), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_144), .B(n_145), .Y(n_486) );
INVx1_ASAP7_75t_L g497 ( .A(n_144), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_144), .A2(n_452), .B(n_510), .C(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_144), .A2(n_452), .B(n_519), .C(n_520), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_145), .B(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_145), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_145), .B(n_207), .Y(n_206) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_145), .B(n_211), .C(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_145), .A2(n_456), .B(n_460), .Y(n_455) );
INVx3_ASAP7_75t_SL g285 ( .A(n_146), .Y(n_285) );
AND2x2_ASAP7_75t_L g331 ( .A(n_146), .B(n_248), .Y(n_331) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_157), .Y(n_146) );
AND2x2_ASAP7_75t_L g168 ( .A(n_147), .B(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_L g262 ( .A(n_147), .B(n_158), .Y(n_262) );
AND2x2_ASAP7_75t_L g266 ( .A(n_147), .B(n_245), .Y(n_266) );
INVx1_ASAP7_75t_L g292 ( .A(n_147), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_147), .B(n_158), .Y(n_314) );
INVx2_ASAP7_75t_L g318 ( .A(n_147), .Y(n_318) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_147), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_147), .B(n_248), .Y(n_395) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_154), .B(n_156), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_154), .A2(n_159), .B(n_165), .Y(n_158) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_154), .A2(n_159), .B(n_165), .Y(n_247) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_154), .A2(n_465), .B(n_471), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_155), .Y(n_154) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_155), .A2(n_216), .B(n_220), .Y(n_215) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g329 ( .A(n_158), .B(n_169), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g339 ( .A(n_167), .Y(n_339) );
NAND2xp33_ASAP7_75t_SL g364 ( .A(n_167), .B(n_256), .Y(n_364) );
AND2x2_ASAP7_75t_L g406 ( .A(n_168), .B(n_248), .Y(n_406) );
AND2x2_ASAP7_75t_L g317 ( .A(n_169), .B(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g380 ( .A(n_169), .Y(n_380) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
AOI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_187), .Y(n_170) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_171), .A2(n_495), .B(n_503), .Y(n_494) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_171), .A2(n_495), .B(n_503), .Y(n_543) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_192), .B(n_193), .Y(n_191) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_172), .A2(n_517), .B(n_521), .Y(n_516) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g209 ( .A(n_173), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_181), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_176), .A2(n_182), .B1(n_201), .B2(n_203), .Y(n_200) );
INVx1_ASAP7_75t_L g536 ( .A(n_176), .Y(n_536) );
AND2x4_ASAP7_75t_L g176 ( .A(n_177), .B(n_180), .Y(n_176) );
INVx1_ASAP7_75t_L g444 ( .A(n_177), .Y(n_444) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
OR2x6_ASAP7_75t_L g452 ( .A(n_178), .B(n_186), .Y(n_452) );
INVxp33_ASAP7_75t_L g500 ( .A(n_178), .Y(n_500) );
INVx1_ASAP7_75t_L g445 ( .A(n_180), .Y(n_445) );
INVxp67_ASAP7_75t_L g534 ( .A(n_182), .Y(n_534) );
NOR2x1p5_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
INVx1_ASAP7_75t_L g501 ( .A(n_185), .Y(n_501) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_188), .A2(n_271), .B1(n_373), .B2(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_213), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_189), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_189), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_198), .Y(n_189) );
INVx2_ASAP7_75t_L g236 ( .A(n_190), .Y(n_236) );
OR2x2_ASAP7_75t_L g240 ( .A(n_190), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_190), .B(n_253), .Y(n_258) );
AND2x4_ASAP7_75t_SL g268 ( .A(n_190), .B(n_199), .Y(n_268) );
OR2x2_ASAP7_75t_L g275 ( .A(n_190), .B(n_215), .Y(n_275) );
OR2x2_ASAP7_75t_L g287 ( .A(n_190), .B(n_199), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_190), .B(n_215), .Y(n_301) );
INVx1_ASAP7_75t_L g306 ( .A(n_190), .Y(n_306) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_190), .Y(n_324) );
AND2x2_ASAP7_75t_L g387 ( .A(n_190), .B(n_307), .Y(n_387) );
INVx2_ASAP7_75t_L g391 ( .A(n_190), .Y(n_391) );
OR2x2_ASAP7_75t_L g398 ( .A(n_190), .B(n_288), .Y(n_398) );
OR2x2_ASAP7_75t_L g420 ( .A(n_190), .B(n_421), .Y(n_420) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_197), .Y(n_190) );
AND2x2_ASAP7_75t_L g237 ( .A(n_198), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_198), .B(n_221), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_198), .B(n_297), .Y(n_359) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
AND2x4_ASAP7_75t_L g307 ( .A(n_199), .B(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_199), .B(n_252), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_199), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_199), .B(n_241), .Y(n_400) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_205), .Y(n_199) );
INVx3_ASAP7_75t_L g505 ( .A(n_208), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_208), .A2(n_505), .B1(n_524), .B2(n_529), .Y(n_523) );
INVx4_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AOI21x1_ASAP7_75t_L g222 ( .A1(n_209), .A2(n_223), .B(n_229), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_209), .B(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_212), .A2(n_452), .B1(n_479), .B2(n_480), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_212), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g267 ( .A(n_213), .B(n_268), .Y(n_267) );
AO221x1_ASAP7_75t_L g341 ( .A1(n_213), .A2(n_256), .B1(n_287), .B2(n_342), .C(n_343), .Y(n_341) );
OAI322xp33_ASAP7_75t_L g393 ( .A1(n_213), .A2(n_313), .A3(n_394), .B1(n_396), .B2(n_397), .C1(n_398), .C2(n_399), .Y(n_393) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_221), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx3_ASAP7_75t_L g235 ( .A(n_215), .Y(n_235) );
INVx2_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
AND2x2_ASAP7_75t_L g253 ( .A(n_215), .B(n_221), .Y(n_253) );
INVx1_ASAP7_75t_L g298 ( .A(n_215), .Y(n_298) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_215), .Y(n_354) );
INVx1_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
OR2x2_ASAP7_75t_L g288 ( .A(n_221), .B(n_241), .Y(n_288) );
INVx2_ASAP7_75t_L g308 ( .A(n_221), .Y(n_308) );
INVx1_ASAP7_75t_L g361 ( .A(n_221), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_221), .B(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OAI21xp33_ASAP7_75t_SL g231 ( .A1(n_232), .A2(n_239), .B(n_242), .Y(n_231) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_232), .A2(n_271), .B1(n_273), .B2(n_277), .C(n_278), .Y(n_270) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
NOR2x1p5_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g357 ( .A(n_236), .Y(n_357) );
INVx1_ASAP7_75t_SL g276 ( .A(n_237), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_237), .A2(n_382), .B(n_384), .Y(n_381) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_238), .Y(n_281) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_241), .Y(n_344) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_244), .A2(n_320), .B(n_325), .C(n_336), .Y(n_319) );
OR2x2_ASAP7_75t_L g409 ( .A(n_244), .B(n_314), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_244), .B(n_277), .Y(n_411) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g251 ( .A(n_245), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g313 ( .A(n_245), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g351 ( .A(n_245), .B(n_318), .Y(n_351) );
OA33x2_ASAP7_75t_L g358 ( .A1(n_245), .A2(n_275), .A3(n_359), .B1(n_360), .B2(n_362), .B3(n_364), .Y(n_358) );
OR2x2_ASAP7_75t_L g369 ( .A(n_245), .B(n_354), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_245), .B(n_293), .Y(n_383) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g271 ( .A(n_247), .B(n_272), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g320 ( .A1(n_247), .A2(n_277), .B1(n_321), .B2(n_322), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_248), .B(n_328), .C(n_361), .Y(n_360) );
AOI322xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .A3(n_256), .B1(n_257), .B2(n_259), .C1(n_263), .C2(n_267), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g356 ( .A(n_252), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_253), .A2(n_268), .B(n_312), .C(n_315), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_254), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
NAND4xp25_ASAP7_75t_SL g375 ( .A(n_255), .B(n_284), .C(n_376), .D(n_378), .Y(n_375) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g265 ( .A(n_260), .Y(n_265) );
OR2x2_ASAP7_75t_L g310 ( .A(n_260), .B(n_262), .Y(n_310) );
AND2x2_ASAP7_75t_L g379 ( .A(n_261), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g384 ( .A(n_265), .B(n_379), .Y(n_384) );
BUFx2_ASAP7_75t_L g377 ( .A(n_266), .Y(n_377) );
INVx1_ASAP7_75t_SL g407 ( .A(n_267), .Y(n_407) );
AND2x4_ASAP7_75t_L g343 ( .A(n_268), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g396 ( .A(n_268), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_289), .C(n_311), .Y(n_269) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_SL g333 ( .A(n_275), .Y(n_333) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_275), .A2(n_402), .B(n_403), .C(n_412), .Y(n_401) );
OR2x2_ASAP7_75t_L g323 ( .A(n_276), .B(n_324), .Y(n_323) );
OAI22xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B1(n_285), .B2(n_286), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_280), .B(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_283), .B(n_340), .Y(n_422) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g397 ( .A(n_284), .B(n_285), .Y(n_397) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B1(n_299), .B2(n_303), .C1(n_304), .C2(n_309), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_292), .Y(n_303) );
AND2x2_ASAP7_75t_L g350 ( .A(n_293), .B(n_351), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_293), .A2(n_366), .B1(n_371), .B2(n_375), .Y(n_365) );
INVx2_ASAP7_75t_SL g418 ( .A(n_293), .Y(n_418) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g374 ( .A(n_298), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_298), .B(n_361), .Y(n_421) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g334 ( .A(n_302), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_304), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g372 ( .A(n_306), .Y(n_372) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_307), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g415 ( .A(n_307), .B(n_344), .Y(n_415) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g419 ( .A(n_317), .Y(n_419) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_330), .B(n_332), .C(n_335), .Y(n_325) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g370 ( .A(n_332), .Y(n_370) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_341), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_385), .C(n_401), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_365), .C(n_381), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B1(n_355), .B2(n_356), .C(n_358), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g394 ( .A(n_380), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g402 ( .A(n_384), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_392), .Y(n_385) );
INVx2_ASAP7_75t_L g408 ( .A(n_387), .Y(n_408) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g399 ( .A(n_390), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_408), .B2(n_409), .C(n_410), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_420), .B2(n_422), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
CKINVDCx11_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_425), .A2(n_433), .B1(n_753), .B2(n_762), .Y(n_761) );
OR2x6_ASAP7_75t_SL g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AND2x6_ASAP7_75t_SL g754 ( .A(n_426), .B(n_428), .Y(n_754) );
OR2x2_ASAP7_75t_L g766 ( .A(n_426), .B(n_428), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_426), .B(n_427), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AO22x1_ASAP7_75t_L g784 ( .A1(n_434), .A2(n_785), .B1(n_786), .B2(n_792), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_434), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g434 ( .A(n_435), .B(n_604), .C(n_670), .D(n_733), .Y(n_434) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_567), .Y(n_435) );
OR3x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_537), .C(n_564), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_472), .B(n_492), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_461), .Y(n_439) );
AND2x2_ASAP7_75t_L g667 ( .A(n_440), .B(n_637), .Y(n_667) );
INVx1_ASAP7_75t_L g740 ( .A(n_440), .Y(n_740) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_453), .Y(n_440) );
INVx2_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_441), .Y(n_555) );
AND2x2_ASAP7_75t_L g559 ( .A(n_441), .B(n_475), .Y(n_559) );
AND2x4_ASAP7_75t_L g575 ( .A(n_441), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_441), .Y(n_579) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_447), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .C(n_446), .Y(n_443) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g525 ( .A(n_452), .Y(n_525) );
AND2x2_ASAP7_75t_L g473 ( .A(n_453), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g556 ( .A(n_453), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_453), .B(n_546), .Y(n_560) );
INVx2_ASAP7_75t_L g574 ( .A(n_453), .Y(n_574) );
AND2x4_ASAP7_75t_L g578 ( .A(n_453), .B(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_453), .Y(n_613) );
OR2x2_ASAP7_75t_L g619 ( .A(n_453), .B(n_464), .Y(n_619) );
NOR2x1_ASAP7_75t_SL g648 ( .A(n_453), .B(n_475), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_453), .B(n_722), .Y(n_750) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x2_ASAP7_75t_L g647 ( .A(n_461), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2x1_ASAP7_75t_L g681 ( .A(n_462), .B(n_474), .Y(n_681) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g488 ( .A(n_464), .Y(n_488) );
INVx2_ASAP7_75t_L g547 ( .A(n_464), .Y(n_547) );
AND2x2_ASAP7_75t_L g570 ( .A(n_464), .B(n_475), .Y(n_570) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_464), .Y(n_597) );
INVx1_ASAP7_75t_L g638 ( .A(n_464), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_487), .Y(n_472) );
AND2x2_ASAP7_75t_L g650 ( .A(n_473), .B(n_545), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_474), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g717 ( .A(n_474), .Y(n_717) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g576 ( .A(n_475), .Y(n_576) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_481), .B(n_486), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_481) );
OAI211xp5_ASAP7_75t_SL g653 ( .A1(n_487), .A2(n_654), .B(n_658), .C(n_664), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x2_ASAP7_75t_SL g569 ( .A(n_489), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g700 ( .A(n_489), .Y(n_700) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g622 ( .A(n_491), .B(n_576), .Y(n_622) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_513), .Y(n_492) );
AOI32xp33_ASAP7_75t_L g658 ( .A1(n_493), .A2(n_642), .A3(n_659), .B1(n_660), .B2(n_662), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
INVx2_ASAP7_75t_L g584 ( .A(n_494), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_494), .B(n_516), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g596 ( .A(n_504), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_504), .B(n_522), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_504), .B(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_504), .Y(n_714) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_504) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OR2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_616), .Y(n_615) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g566 ( .A(n_514), .B(n_540), .Y(n_566) );
AND2x2_ASAP7_75t_L g715 ( .A(n_514), .B(n_713), .Y(n_715) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g552 ( .A(n_516), .Y(n_552) );
AND2x4_ASAP7_75t_L g591 ( .A(n_516), .B(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_L g625 ( .A(n_516), .Y(n_625) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_516), .Y(n_633) );
AND2x2_ASAP7_75t_L g642 ( .A(n_516), .B(n_522), .Y(n_642) );
INVx1_ASAP7_75t_L g726 ( .A(n_516), .Y(n_726) );
INVx2_ASAP7_75t_L g563 ( .A(n_522), .Y(n_563) );
INVx1_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
INVx1_ASAP7_75t_L g657 ( .A(n_522), .Y(n_657) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_530), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI32xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_548), .A3(n_553), .B1(n_557), .B2(n_561), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_539), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_540), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g641 ( .A(n_540), .B(n_642), .Y(n_641) );
INVxp67_ASAP7_75t_L g666 ( .A(n_540), .Y(n_666) );
AND2x2_ASAP7_75t_L g747 ( .A(n_540), .B(n_589), .Y(n_747) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g562 ( .A(n_542), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g661 ( .A(n_542), .B(n_584), .Y(n_661) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_542), .B(n_563), .Y(n_683) );
NOR2x1_ASAP7_75t_L g725 ( .A(n_542), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g592 ( .A(n_543), .Y(n_592) );
INVx1_ASAP7_75t_L g616 ( .A(n_543), .Y(n_616) );
AND2x2_ASAP7_75t_L g631 ( .A(n_543), .B(n_563), .Y(n_631) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g659 ( .A(n_545), .B(n_648), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_545), .B(n_578), .Y(n_729) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_546), .Y(n_698) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_547), .Y(n_680) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g581 ( .A(n_550), .B(n_582), .Y(n_581) );
NOR2xp67_ASAP7_75t_L g665 ( .A(n_550), .B(n_666), .Y(n_665) );
NOR2xp67_ASAP7_75t_SL g752 ( .A(n_550), .B(n_690), .Y(n_752) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g609 ( .A(n_552), .B(n_563), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_553), .B(n_619), .Y(n_677) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_554), .B(n_570), .Y(n_643) );
AND2x4_ASAP7_75t_SL g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_556), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g708 ( .A(n_556), .B(n_579), .Y(n_708) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_556), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_557), .B(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
OR2x2_ASAP7_75t_L g679 ( .A(n_558), .B(n_680), .Y(n_679) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_558), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g668 ( .A(n_559), .B(n_613), .Y(n_668) );
INVxp33_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g582 ( .A(n_562), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g742 ( .A(n_562), .B(n_624), .Y(n_742) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_585), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .B(n_580), .Y(n_568) );
AND2x2_ASAP7_75t_L g703 ( .A(n_570), .B(n_578), .Y(n_703) );
NAND2xp33_ASAP7_75t_R g571 ( .A(n_572), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g745 ( .A(n_574), .Y(n_745) );
INVx4_ASAP7_75t_L g603 ( .A(n_575), .Y(n_603) );
INVx1_ASAP7_75t_L g722 ( .A(n_576), .Y(n_722) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g716 ( .A(n_578), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_578), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_581), .A2(n_646), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g610 ( .A(n_584), .B(n_596), .Y(n_610) );
AND2x2_ASAP7_75t_L g624 ( .A(n_584), .B(n_625), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_593), .B(n_598), .C(n_601), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g672 ( .A(n_588), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g600 ( .A(n_589), .Y(n_600) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g660 ( .A(n_590), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g669 ( .A(n_590), .B(n_591), .Y(n_669) );
INVx1_ASAP7_75t_L g701 ( .A(n_590), .Y(n_701) );
AND2x4_ASAP7_75t_L g682 ( .A(n_591), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g704 ( .A(n_591), .B(n_595), .Y(n_704) );
AND2x2_ASAP7_75t_L g712 ( .A(n_591), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g687 ( .A(n_595), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_595), .B(n_609), .Y(n_689) );
AND2x2_ASAP7_75t_L g692 ( .A(n_595), .B(n_642), .Y(n_692) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_596), .B(n_657), .Y(n_706) );
AND2x2_ASAP7_75t_L g634 ( .A(n_597), .B(n_622), .Y(n_634) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g730 ( .A(n_600), .B(n_610), .Y(n_730) );
BUFx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_602), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g614 ( .A(n_603), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_603), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_644), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_628), .Y(n_605) );
OAI222xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_611), .B1(n_615), .B2(n_617), .C1(n_620), .C2(n_623), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_613), .B(n_622), .Y(n_621) );
OR2x6_ASAP7_75t_L g693 ( .A(n_613), .B(n_663), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g696 ( .A(n_613), .B(n_616), .C(n_632), .D(n_697), .E(n_699), .Y(n_696) );
NAND2x1_ASAP7_75t_L g732 ( .A(n_614), .B(n_618), .Y(n_732) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_619), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_621), .A2(n_712), .B1(n_715), .B2(n_716), .Y(n_711) );
INVx2_ASAP7_75t_L g663 ( .A(n_622), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_622), .B(n_638), .Y(n_675) );
INVx3_ASAP7_75t_L g710 ( .A(n_623), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
AND2x2_ASAP7_75t_L g655 ( .A(n_624), .B(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g688 ( .A(n_624), .Y(n_688) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g651 ( .A(n_627), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_629), .B(n_640), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .B(n_635), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g639 ( .A(n_631), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_634), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_639), .Y(n_635) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_SL g721 ( .A(n_638), .B(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_653), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .B(n_651), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g690 ( .A(n_661), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_664) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_694), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .C(n_684), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OA21x2_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B(n_682), .Y(n_676) );
NAND2xp33_ASAP7_75t_SL g678 ( .A(n_679), .B(n_681), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_691), .B(n_693), .Y(n_684) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_689), .C(n_690), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_688), .A2(n_728), .B1(n_730), .B2(n_731), .Y(n_727) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_718), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_696), .B(n_702), .C(n_709), .D(n_711), .Y(n_695) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g707 ( .A(n_698), .B(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g738 ( .A(n_701), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_707), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_707), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g718 ( .A1(n_719), .A2(n_723), .B(n_727), .Y(n_718) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_748), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_738), .B(n_739), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_743), .B2(n_746), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx11_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_755), .A2(n_761), .B(n_763), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
BUFx3_ASAP7_75t_L g795 ( .A(n_769), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI21x1_ASAP7_75t_SL g776 ( .A1(n_772), .A2(n_777), .B(n_779), .Y(n_776) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx3_ASAP7_75t_L g778 ( .A(n_775), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .B1(n_784), .B2(n_793), .Y(n_779) );
INVx1_ASAP7_75t_L g793 ( .A(n_780), .Y(n_793) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g792 ( .A(n_786), .Y(n_792) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx3_ASAP7_75t_SL g810 ( .A(n_800), .Y(n_810) );
OR2x2_ASAP7_75t_SL g800 ( .A(n_801), .B(n_803), .Y(n_800) );
CKINVDCx16_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
endmodule