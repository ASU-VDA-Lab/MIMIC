module fake_ariane_1795_n_1111 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1111);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1111;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_1029;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_926;
wire n_813;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_1099;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_455;
wire n_429;
wire n_238;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_931;
wire n_827;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_26),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_78),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_52),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_55),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_133),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_71),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_50),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_138),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_113),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_151),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_99),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_131),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_80),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_93),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_33),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_36),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_121),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_105),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_162),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_115),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_23),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_28),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_92),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_200),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_110),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_12),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_41),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_146),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_191),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_97),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_81),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_79),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_61),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_111),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_207),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_182),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_118),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_65),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_129),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_56),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_147),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_169),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_47),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_87),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_101),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_34),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_4),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_89),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_252),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_283),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_283),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_257),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_225),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_220),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_244),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_239),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_251),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_263),
.Y(n_316)
);

BUFx6f_ASAP7_75t_SL g317 ( 
.A(n_278),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_260),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_256),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_235),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_277),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_261),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_219),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_235),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_0),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_310),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_332),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_333),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_334),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_232),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_313),
.B(n_265),
.Y(n_350)
);

CKINVDCx6p67_ASAP7_75t_R g351 ( 
.A(n_302),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_336),
.A2(n_284),
.B(n_224),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_313),
.B(n_230),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_262),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_337),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_297),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_284),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_317),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_304),
.B(n_268),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

CKINVDCx6p67_ASAP7_75t_R g368 ( 
.A(n_325),
.Y(n_368)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_232),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_323),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_328),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_319),
.B(n_222),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_301),
.B(n_223),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_300),
.B(n_232),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_232),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_301),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_295),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_296),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_290),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_290),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_226),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_371),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_339),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_339),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_315),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_228),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_R g405 ( 
.A(n_352),
.B(n_342),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_368),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_348),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_380),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_380),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_382),
.B(n_380),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_380),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_379),
.B(n_315),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_364),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_380),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_382),
.A2(n_255),
.B1(n_288),
.B2(n_286),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_390),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_390),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_R g429 ( 
.A(n_352),
.B(n_318),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_385),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_231),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_390),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_390),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_390),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_373),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_387),
.B(n_373),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_387),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_392),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_365),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_361),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_365),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_386),
.Y(n_448)
);

AOI21x1_ASAP7_75t_L g449 ( 
.A1(n_352),
.A2(n_369),
.B(n_338),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_359),
.B(n_234),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_338),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_345),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_392),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_389),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_389),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_384),
.B(n_236),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_360),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_391),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_391),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_354),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_364),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_354),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NOR2x1p5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_366),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_462),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_353),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_L g471 ( 
.A(n_416),
.B(n_364),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_464),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_395),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_403),
.B(n_383),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_400),
.B(n_381),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_417),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_418),
.A2(n_414),
.B1(n_446),
.B2(n_404),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_383),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_455),
.B(n_362),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_411),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_412),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_405),
.A2(n_457),
.B1(n_425),
.B2(n_448),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_424),
.B(n_379),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_444),
.B(n_379),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_394),
.B(n_381),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_405),
.B(n_372),
.C(n_363),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_362),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_420),
.B(n_350),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_430),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_434),
.A2(n_352),
.B1(n_377),
.B2(n_367),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_435),
.A2(n_441),
.B1(n_445),
.B2(n_456),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_378),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_456),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_437),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_401),
.B(n_375),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_429),
.A2(n_378),
.B1(n_363),
.B2(n_372),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_406),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_451),
.B(n_378),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_432),
.B(n_363),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_410),
.B(n_362),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_428),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_396),
.B(n_454),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_413),
.B(n_363),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_421),
.B(n_318),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_422),
.B(n_367),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_427),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_377),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_463),
.B(n_343),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_421),
.B(n_341),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_402),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_440),
.B(n_364),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_438),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_408),
.B(n_343),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_402),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_449),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_463),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

INVx4_ASAP7_75t_SL g539 ( 
.A(n_429),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_409),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_461),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_341),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_460),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_452),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_452),
.B(n_372),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_393),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_341),
.Y(n_548)
);

AOI22x1_ASAP7_75t_L g549 ( 
.A1(n_531),
.A2(n_372),
.B1(n_358),
.B2(n_357),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_358),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_545),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_544),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_465),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_468),
.B(n_372),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_470),
.Y(n_555)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_L g557 ( 
.A1(n_490),
.A2(n_357),
.B1(n_346),
.B2(n_282),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_498),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_542),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_484),
.B(n_346),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_544),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_539),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_477),
.B(n_237),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_490),
.B(n_238),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_477),
.B(n_240),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_532),
.B(n_242),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_500),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_546),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_344),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_532),
.B(n_344),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_467),
.B(n_281),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_478),
.Y(n_575)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_539),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_504),
.B(n_243),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_504),
.B(n_513),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_513),
.B(n_246),
.Y(n_579)
);

OAI221xp5_ASAP7_75t_L g580 ( 
.A1(n_467),
.A2(n_280),
.B1(n_275),
.B2(n_273),
.C(n_272),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_495),
.Y(n_581)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_476),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_501),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_510),
.Y(n_586)
);

NAND2x1p5_ASAP7_75t_L g587 ( 
.A(n_511),
.B(n_5),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

AOI22x1_ASAP7_75t_L g589 ( 
.A1(n_506),
.A2(n_271),
.B1(n_259),
.B2(n_254),
.Y(n_589)
);

NAND2x1p5_ASAP7_75t_L g590 ( 
.A(n_511),
.B(n_5),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_507),
.B(n_6),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_519),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_473),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_483),
.B(n_250),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_475),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_515),
.B(n_6),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_518),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_499),
.B(n_253),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_495),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_516),
.B(n_469),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_485),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_537),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_520),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_479),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_505),
.B(n_10),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

AO22x2_ASAP7_75t_L g612 ( 
.A1(n_539),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_609),
.B(n_474),
.C(n_480),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_603),
.B(n_487),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_578),
.A2(n_471),
.B(n_508),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_601),
.B(n_543),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_533),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_558),
.A2(n_480),
.B1(n_503),
.B2(n_547),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_561),
.B(n_533),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_577),
.A2(n_514),
.B(n_535),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_581),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_556),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_580),
.B(n_523),
.C(n_522),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_559),
.A2(n_547),
.B1(n_469),
.B2(n_523),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_563),
.B(n_543),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_560),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_569),
.B(n_528),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_573),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_579),
.A2(n_491),
.B(n_492),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_574),
.A2(n_466),
.B(n_525),
.C(n_533),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_551),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_554),
.A2(n_534),
.B(n_496),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_570),
.A2(n_534),
.B(n_496),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_598),
.B(n_541),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_594),
.A2(n_534),
.B(n_496),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_608),
.B(n_541),
.C(n_493),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_594),
.B(n_493),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_599),
.A2(n_494),
.B(n_502),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_566),
.A2(n_494),
.B(n_529),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_610),
.B(n_541),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_568),
.B(n_488),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_565),
.A2(n_509),
.B1(n_502),
.B2(n_530),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_599),
.A2(n_540),
.B(n_536),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_SL g646 ( 
.A(n_587),
.B(n_509),
.C(n_11),
.Y(n_646)
);

AOI21xp33_ASAP7_75t_L g647 ( 
.A1(n_557),
.A2(n_530),
.B(n_536),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_567),
.A2(n_538),
.B1(n_497),
.B2(n_527),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_610),
.B(n_13),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_605),
.A2(n_538),
.B(n_527),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_562),
.B(n_497),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_551),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_611),
.A2(n_538),
.B(n_527),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_611),
.A2(n_497),
.B(n_521),
.Y(n_654)
);

CKINVDCx10_ASAP7_75t_R g655 ( 
.A(n_582),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_550),
.B(n_521),
.Y(n_656)
);

AO32x1_ASAP7_75t_L g657 ( 
.A1(n_583),
.A2(n_521),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_595),
.A2(n_30),
.B(n_29),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_581),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_591),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_550),
.B(n_16),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_590),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_593),
.B(n_18),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_581),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_553),
.Y(n_665)
);

NOR3xp33_ASAP7_75t_L g666 ( 
.A(n_593),
.B(n_19),
.C(n_20),
.Y(n_666)
);

NAND2x1_ASAP7_75t_L g667 ( 
.A(n_592),
.B(n_31),
.Y(n_667)
);

NAND2x1_ASAP7_75t_L g668 ( 
.A(n_592),
.B(n_32),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_548),
.B(n_21),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_602),
.B(n_21),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_556),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_615),
.A2(n_597),
.B(n_596),
.C(n_606),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_617),
.B(n_555),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_616),
.A2(n_549),
.B(n_564),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_666),
.A2(n_572),
.B(n_571),
.C(n_588),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_652),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_638),
.A2(n_612),
.B1(n_564),
.B2(n_576),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_655),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_627),
.B(n_555),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_622),
.A2(n_612),
.B(n_576),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_R g682 ( 
.A(n_624),
.B(n_582),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_613),
.A2(n_585),
.B(n_586),
.C(n_584),
.Y(n_683)
);

AO21x1_ASAP7_75t_L g684 ( 
.A1(n_644),
.A2(n_589),
.B(n_604),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_648),
.A2(n_604),
.B(n_589),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_631),
.A2(n_22),
.B(n_23),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_632),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_671),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_634),
.A2(n_24),
.B(n_25),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_621),
.B(n_27),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_643),
.B(n_35),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_628),
.B(n_217),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_633),
.B(n_642),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_665),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_614),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_645),
.A2(n_37),
.B(n_38),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_630),
.Y(n_697)
);

CKINVDCx6p67_ASAP7_75t_R g698 ( 
.A(n_618),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_661),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_629),
.B(n_39),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_626),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_635),
.A2(n_44),
.B(n_46),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_620),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_659),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_646),
.A2(n_662),
.B(n_647),
.C(n_639),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_641),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_620),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_636),
.B(n_649),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_625),
.B(n_651),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_663),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_660),
.A2(n_54),
.B(n_57),
.C(n_58),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_654),
.A2(n_59),
.B(n_60),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_670),
.B(n_62),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_659),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_670),
.B(n_216),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_619),
.B(n_63),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_SL g717 ( 
.A(n_669),
.B(n_64),
.C(n_66),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_659),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_650),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_623),
.B(n_72),
.Y(n_720)
);

AO21x1_ASAP7_75t_L g721 ( 
.A1(n_640),
.A2(n_73),
.B(n_74),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_623),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_664),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_656),
.Y(n_725)
);

NOR2x1_ASAP7_75t_SL g726 ( 
.A(n_653),
.B(n_75),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_637),
.B(n_76),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_710),
.B(n_668),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_707),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

BUFx2_ASAP7_75t_SL g731 ( 
.A(n_688),
.Y(n_731)
);

NAND2x1p5_ASAP7_75t_L g732 ( 
.A(n_704),
.B(n_667),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_714),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_693),
.B(n_77),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_672),
.Y(n_735)
);

CKINVDCx14_ASAP7_75t_R g736 ( 
.A(n_682),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_698),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_718),
.Y(n_738)
);

BUFx2_ASAP7_75t_R g739 ( 
.A(n_679),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_708),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_694),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_677),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_706),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_695),
.Y(n_744)
);

INVx3_ASAP7_75t_SL g745 ( 
.A(n_722),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_722),
.Y(n_746)
);

BUFx12f_ASAP7_75t_L g747 ( 
.A(n_703),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_704),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_724),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_690),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_691),
.B(n_658),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_697),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_723),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_725),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_674),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_684),
.Y(n_756)
);

BUFx8_ASAP7_75t_SL g757 ( 
.A(n_713),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

INVx5_ASAP7_75t_SL g759 ( 
.A(n_676),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_699),
.B(n_82),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_678),
.B(n_83),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_715),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_709),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_683),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_681),
.A2(n_657),
.B1(n_85),
.B2(n_86),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_687),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_720),
.Y(n_767)
);

INVx6_ASAP7_75t_SL g768 ( 
.A(n_726),
.Y(n_768)
);

CKINVDCx11_ASAP7_75t_R g769 ( 
.A(n_705),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_692),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_716),
.A2(n_657),
.B1(n_88),
.B2(n_90),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_721),
.Y(n_772)
);

BUFx6f_ASAP7_75t_SL g773 ( 
.A(n_717),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_719),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_673),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_700),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_727),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_689),
.Y(n_778)
);

BUFx4f_ASAP7_75t_L g779 ( 
.A(n_711),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_685),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_689),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_686),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_686),
.Y(n_783)
);

BUFx12f_ASAP7_75t_L g784 ( 
.A(n_681),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_701),
.Y(n_785)
);

BUFx12f_ASAP7_75t_L g786 ( 
.A(n_702),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_675),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_675),
.Y(n_788)
);

OAI21x1_ASAP7_75t_SL g789 ( 
.A1(n_776),
.A2(n_696),
.B(n_712),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_733),
.B(n_696),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_741),
.Y(n_791)
);

OAI22xp33_ASAP7_75t_L g792 ( 
.A1(n_747),
.A2(n_657),
.B1(n_91),
.B2(n_94),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_782),
.A2(n_84),
.B(n_95),
.Y(n_793)
);

AO21x2_ASAP7_75t_L g794 ( 
.A1(n_756),
.A2(n_96),
.B(n_98),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_731),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_751),
.A2(n_100),
.B(n_102),
.C(n_103),
.Y(n_796)
);

CKINVDCx11_ASAP7_75t_R g797 ( 
.A(n_729),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_742),
.Y(n_798)
);

INVx4_ASAP7_75t_SL g799 ( 
.A(n_745),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_733),
.B(n_104),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_769),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_787),
.A2(n_215),
.B(n_112),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_745),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_777),
.A2(n_109),
.B(n_114),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_763),
.B(n_116),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_767),
.A2(n_119),
.B(n_120),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_787),
.A2(n_122),
.B(n_124),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_746),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_779),
.A2(n_125),
.B(n_126),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_732),
.A2(n_756),
.B(n_764),
.Y(n_810)
);

AOI22x1_ASAP7_75t_L g811 ( 
.A1(n_766),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

OAI21x1_ASAP7_75t_SL g813 ( 
.A1(n_771),
.A2(n_132),
.B(n_134),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_737),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_769),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_788),
.A2(n_139),
.B(n_140),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_SL g817 ( 
.A1(n_784),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_817)
);

AOI221xp5_ASAP7_75t_L g818 ( 
.A1(n_779),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.C(n_150),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_758),
.B(n_214),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_737),
.Y(n_820)
);

AO21x2_ASAP7_75t_L g821 ( 
.A1(n_788),
.A2(n_152),
.B(n_153),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_735),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_732),
.A2(n_154),
.B(n_155),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_740),
.B(n_156),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_744),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_757),
.B(n_739),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_767),
.B(n_157),
.Y(n_827)
);

CKINVDCx14_ASAP7_75t_R g828 ( 
.A(n_736),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_735),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_770),
.A2(n_158),
.B(n_159),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_767),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_751),
.A2(n_165),
.B(n_166),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_740),
.B(n_167),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_750),
.A2(n_168),
.B(n_170),
.C(n_171),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_755),
.B(n_213),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_761),
.A2(n_775),
.B1(n_773),
.B2(n_765),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_748),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_775),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_757),
.B(n_175),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_728),
.A2(n_176),
.B(n_177),
.C(n_178),
.Y(n_841)
);

NAND2x1_ASAP7_75t_L g842 ( 
.A(n_763),
.B(n_180),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_767),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_738),
.B(n_181),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_730),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_837),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_SL g847 ( 
.A(n_836),
.B(n_765),
.C(n_728),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_791),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_790),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_790),
.B(n_753),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_825),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_839),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_799),
.B(n_753),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_814),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_798),
.B(n_783),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_810),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_819),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_812),
.B(n_783),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_816),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_803),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_819),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_835),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_827),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_835),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_795),
.B(n_781),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_832),
.B(n_781),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_845),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_832),
.A2(n_773),
.B1(n_759),
.B2(n_786),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_816),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_802),
.Y(n_870)
);

OAI321xp33_ASAP7_75t_L g871 ( 
.A1(n_809),
.A2(n_763),
.A3(n_760),
.B1(n_762),
.B2(n_734),
.C(n_780),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_843),
.B(n_778),
.Y(n_872)
);

CKINVDCx11_ASAP7_75t_R g873 ( 
.A(n_797),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_803),
.B(n_763),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_843),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_821),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_802),
.B(n_743),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_806),
.B(n_778),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_799),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_821),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_794),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_818),
.A2(n_759),
.B1(n_762),
.B2(n_774),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_827),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_822),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_820),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_800),
.B(n_762),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_794),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_800),
.B(n_754),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_844),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_848),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_822),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_846),
.B(n_822),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_882),
.A2(n_809),
.B(n_806),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_846),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_850),
.B(n_829),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_851),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_884),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_873),
.B(n_828),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_866),
.A2(n_759),
.B1(n_772),
.B2(n_774),
.Y(n_899)
);

INVx6_ASAP7_75t_SL g900 ( 
.A(n_888),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_847),
.A2(n_774),
.B(n_831),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_SL g902 ( 
.A(n_879),
.B(n_829),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_888),
.B(n_829),
.Y(n_903)
);

BUFx5_ASAP7_75t_L g904 ( 
.A(n_876),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_850),
.B(n_808),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_866),
.A2(n_818),
.B(n_815),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_851),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_868),
.A2(n_815),
.B1(n_792),
.B2(n_774),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_873),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_848),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_854),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_858),
.B(n_762),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_858),
.B(n_826),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_852),
.Y(n_914)
);

AO21x1_ASAP7_75t_L g915 ( 
.A1(n_889),
.A2(n_831),
.B(n_840),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_885),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_860),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_890),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_894),
.B(n_849),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_913),
.B(n_849),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_891),
.B(n_849),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_904),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_909),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_892),
.B(n_865),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_905),
.B(n_865),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_890),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_904),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_891),
.B(n_850),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_904),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_910),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_904),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_905),
.B(n_855),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_898),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_912),
.B(n_857),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_914),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_917),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_896),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_915),
.B(n_857),
.Y(n_938)
);

AO21x2_ASAP7_75t_L g939 ( 
.A1(n_906),
.A2(n_887),
.B(n_876),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_907),
.B(n_855),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_938),
.A2(n_859),
.B(n_869),
.Y(n_941)
);

AO21x2_ASAP7_75t_L g942 ( 
.A1(n_939),
.A2(n_893),
.B(n_901),
.Y(n_942)
);

AO21x2_ASAP7_75t_L g943 ( 
.A1(n_939),
.A2(n_887),
.B(n_880),
.Y(n_943)
);

AO21x2_ASAP7_75t_L g944 ( 
.A1(n_939),
.A2(n_880),
.B(n_929),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_936),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_928),
.A2(n_902),
.B(n_908),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_918),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_933),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_918),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_922),
.A2(n_859),
.B(n_869),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_926),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_933),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_926),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_928),
.A2(n_871),
.B(n_903),
.Y(n_954)
);

OAI22xp33_ASAP7_75t_L g955 ( 
.A1(n_940),
.A2(n_886),
.B1(n_863),
.B2(n_883),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_924),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_935),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_944),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_949),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_948),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_948),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_948),
.Y(n_962)
);

NAND4xp25_ASAP7_75t_SL g963 ( 
.A(n_946),
.B(n_923),
.C(n_925),
.D(n_932),
.Y(n_963)
);

INVx5_ASAP7_75t_SL g964 ( 
.A(n_942),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_956),
.B(n_925),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_947),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_944),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_949),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_947),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_956),
.B(n_934),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_952),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_959),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_970),
.B(n_961),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_968),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_960),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_971),
.B(n_952),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_962),
.B(n_952),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_966),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_962),
.B(n_952),
.Y(n_979)
);

OAI22xp33_ASAP7_75t_L g980 ( 
.A1(n_973),
.A2(n_954),
.B1(n_964),
.B2(n_969),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_972),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_974),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_977),
.B(n_963),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_978),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_975),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_979),
.B(n_969),
.C(n_966),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_985),
.B(n_977),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_980),
.A2(n_964),
.B1(n_942),
.B2(n_967),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_984),
.B(n_976),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_981),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_986),
.B(n_945),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_965),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_982),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_981),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_985),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_985),
.B(n_957),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_986),
.B(n_964),
.C(n_967),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_995),
.B(n_911),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_990),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_987),
.B(n_739),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_992),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_990),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_991),
.Y(n_1003)
);

NOR2x1_ASAP7_75t_L g1004 ( 
.A(n_997),
.B(n_942),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_994),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_996),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1006),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_998),
.B(n_989),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_999),
.Y(n_1009)
);

XOR2x2_ASAP7_75t_L g1010 ( 
.A(n_1000),
.B(n_988),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_998),
.B(n_993),
.Y(n_1011)
);

AOI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_1001),
.A2(n_958),
.B(n_944),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_1005),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_1003),
.B(n_947),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_1004),
.A2(n_951),
.B1(n_953),
.B2(n_957),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1013),
.B(n_1002),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1007),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1014),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1009),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_1011),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1008),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_SL g1022 ( 
.A(n_1010),
.B(n_736),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_951),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1020),
.B(n_1012),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_1022),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1021),
.B(n_916),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_SL g1027 ( 
.A1(n_1017),
.A2(n_860),
.B(n_958),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_1016),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1018),
.B(n_951),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1019),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1023),
.B(n_953),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_1026),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_1030),
.B(n_796),
.C(n_955),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_811),
.C(n_824),
.Y(n_1034)
);

NAND4xp75_ASAP7_75t_L g1035 ( 
.A(n_1028),
.B(n_833),
.C(n_805),
.D(n_867),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1029),
.Y(n_1036)
);

AOI221x1_ASAP7_75t_L g1037 ( 
.A1(n_1024),
.A2(n_957),
.B1(n_930),
.B2(n_922),
.C(n_931),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_1027),
.B(n_941),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_1036),
.Y(n_1039)
);

AOI211xp5_ASAP7_75t_L g1040 ( 
.A1(n_1032),
.A2(n_1031),
.B(n_841),
.C(n_834),
.Y(n_1040)
);

AOI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_1038),
.A2(n_813),
.B1(n_943),
.B2(n_930),
.C(n_935),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1037),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1039),
.A2(n_1035),
.B1(n_927),
.B2(n_929),
.Y(n_1044)
);

AOI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_1042),
.A2(n_1043),
.B1(n_1040),
.B2(n_1041),
.C(n_943),
.Y(n_1045)
);

AOI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_1042),
.A2(n_943),
.B1(n_927),
.B2(n_931),
.C(n_862),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1039),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_1042),
.A2(n_861),
.B1(n_864),
.B2(n_870),
.C(n_801),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1039),
.Y(n_1049)
);

INVx8_ASAP7_75t_L g1050 ( 
.A(n_1039),
.Y(n_1050)
);

XOR2xp5_ASAP7_75t_L g1051 ( 
.A(n_1039),
.B(n_817),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_1039),
.A2(n_842),
.B(n_838),
.C(n_874),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1047),
.A2(n_884),
.B1(n_768),
.B2(n_924),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_1049),
.B(n_884),
.Y(n_1054)
);

NAND3x1_ASAP7_75t_SL g1055 ( 
.A(n_1045),
.B(n_920),
.C(n_932),
.Y(n_1055)
);

OAI321xp33_ASAP7_75t_L g1056 ( 
.A1(n_1046),
.A2(n_863),
.A3(n_856),
.B1(n_903),
.B2(n_934),
.C(n_878),
.Y(n_1056)
);

OAI211xp5_ASAP7_75t_SL g1057 ( 
.A1(n_1050),
.A2(n_899),
.B(n_883),
.C(n_940),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1048),
.B(n_920),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1051),
.A2(n_768),
.B1(n_919),
.B2(n_897),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1044),
.A2(n_919),
.B1(n_897),
.B2(n_785),
.Y(n_1060)
);

OAI32xp33_ASAP7_75t_L g1061 ( 
.A1(n_1052),
.A2(n_878),
.A3(n_875),
.B1(n_883),
.B2(n_870),
.Y(n_1061)
);

OAI32xp33_ASAP7_75t_L g1062 ( 
.A1(n_1047),
.A2(n_878),
.A3(n_875),
.B1(n_856),
.B2(n_941),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1054),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1055),
.Y(n_1064)
);

INVx3_ASAP7_75t_SL g1065 ( 
.A(n_1058),
.Y(n_1065)
);

AND4x1_ASAP7_75t_L g1066 ( 
.A(n_1061),
.B(n_900),
.C(n_186),
.D(n_188),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1060),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_1053),
.B(n_184),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_1056),
.B(n_189),
.C(n_190),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1057),
.B(n_950),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1059),
.A2(n_853),
.B1(n_950),
.B2(n_895),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_1062),
.B(n_875),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_1058),
.B(n_928),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_1058),
.B(n_853),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1054),
.B(n_921),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1063),
.B(n_853),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1064),
.B(n_823),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1065),
.B(n_895),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_1067),
.B(n_192),
.Y(n_1079)
);

AOI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1068),
.A2(n_807),
.B(n_793),
.C(n_804),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1069),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1073),
.B(n_772),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_772),
.Y(n_1083)
);

XNOR2xp5_ASAP7_75t_L g1084 ( 
.A(n_1066),
.B(n_830),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1079),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1081),
.B(n_1075),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1078),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1076),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1076),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1077),
.A2(n_1072),
.B1(n_1070),
.B2(n_1071),
.Y(n_1090)
);

XNOR2x1_ASAP7_75t_L g1091 ( 
.A(n_1084),
.B(n_194),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1088),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1089),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1086),
.A2(n_1083),
.B(n_1082),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1095),
.A2(n_1087),
.B(n_1093),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_1096),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1097),
.A2(n_1090),
.B1(n_1091),
.B2(n_1085),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_1094),
.B(n_1080),
.C(n_199),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_900),
.B1(n_928),
.B2(n_921),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1098),
.B(n_196),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_863),
.B1(n_921),
.B2(n_785),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_921),
.B(n_863),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_863),
.B1(n_780),
.B2(n_772),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_1102),
.B1(n_872),
.B2(n_785),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1101),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1106),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1105),
.A2(n_204),
.B(n_205),
.Y(n_1108)
);

AO221x1_ASAP7_75t_L g1109 ( 
.A1(n_1104),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.C(n_785),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_1107),
.A2(n_881),
.B1(n_937),
.B2(n_877),
.C(n_789),
.Y(n_1110)
);

AOI211xp5_ASAP7_75t_L g1111 ( 
.A1(n_1110),
.A2(n_1109),
.B(n_1108),
.C(n_881),
.Y(n_1111)
);


endmodule