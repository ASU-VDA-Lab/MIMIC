module real_jpeg_29014_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_344, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_344;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_0),
.Y(n_107)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_1),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_23),
.B1(n_26),
.B2(n_117),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_117),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_1),
.A2(n_60),
.B1(n_62),
.B2(n_117),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_32),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_32),
.B(n_164),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_122),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_57),
.B(n_60),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_79),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_2),
.A2(n_99),
.B1(n_102),
.B2(n_215),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_49),
.B1(n_60),
.B2(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_4),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_4),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_23),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_38),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_7),
.A2(n_38),
.B1(n_60),
.B2(n_62),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_8),
.A2(n_28),
.B1(n_32),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_8),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_119),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_8),
.A2(n_60),
.B1(n_62),
.B2(n_119),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_119),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_25),
.B1(n_60),
.B2(n_62),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_10),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_10),
.A2(n_47),
.B1(n_60),
.B2(n_62),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_47),
.Y(n_272)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_23),
.B1(n_26),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_12),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_12),
.A2(n_28),
.B1(n_32),
.B2(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_124),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_12),
.A2(n_60),
.B1(n_62),
.B2(n_124),
.Y(n_215)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_15),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_342),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_84),
.B(n_340),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_20),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_21),
.A2(n_45),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_22),
.A2(n_34),
.B(n_83),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_22),
.A2(n_27),
.B(n_34),
.Y(n_342)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_27),
.B(n_30),
.C(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_30),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_23),
.B(n_122),
.CON(n_121),
.SN(n_121)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_27),
.A2(n_34),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_28),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_28),
.A2(n_35),
.B1(n_121),
.B2(n_136),
.Y(n_135)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_28),
.A2(n_54),
.A3(n_68),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_30),
.B(n_32),
.Y(n_136)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_33),
.A2(n_46),
.B(n_50),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_34),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_40),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_76),
.C(n_81),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_41),
.A2(n_42),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.C(n_65),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_43),
.A2(n_44),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_45),
.A2(n_50),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_45),
.A2(n_50),
.B1(n_130),
.B2(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_51),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_51),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_51),
.A2(n_65),
.B1(n_308),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_59),
.B(n_63),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_63),
.B(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_52),
.A2(n_59),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_52),
.A2(n_172),
.B(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_52),
.A2(n_59),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_52),
.A2(n_59),
.B1(n_171),
.B2(n_190),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_52),
.A2(n_59),
.B1(n_94),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_52),
.A2(n_112),
.B(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_55),
.B(n_69),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_55),
.A2(n_58),
.B(n_122),
.C(n_192),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_59),
.B(n_122),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_62),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_64),
.B(n_113),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_65),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_66),
.A2(n_78),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_74),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_74),
.B1(n_116),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_67),
.A2(n_74),
.B1(n_147),
.B2(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_67),
.B(n_73),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_67),
.A2(n_74),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_72),
.A2(n_79),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_78),
.A2(n_80),
.B(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_78),
.A2(n_258),
.B(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_81),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_333),
.B(n_339),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_303),
.A3(n_325),
.B1(n_331),
.B2(n_332),
.C(n_344),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_284),
.B(n_302),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_262),
.B(n_283),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_154),
.B(n_239),
.C(n_261),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_139),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_90),
.B(n_139),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_125),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_109),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_92),
.B(n_109),
.C(n_125),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_93),
.B(n_98),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_95),
.B(n_182),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B(n_104),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_99),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_99),
.A2(n_207),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_99),
.A2(n_151),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_100),
.A2(n_105),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_100),
.A2(n_202),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_120),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_122),
.B(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_134),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_127),
.B(n_132),
.C(n_134),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_137),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_140),
.A2(n_141),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_152),
.B(n_201),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_238),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_231),
.B(n_237),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_183),
.B(n_230),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_173),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_158),
.B(n_173),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.C(n_169),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_159),
.A2(n_160),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_162),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_180),
.C(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_224),
.B(n_229),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_203),
.B(n_223),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_186),
.B(n_193),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_211),
.B(n_222),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_209),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_217),
.B(n_221),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_259),
.B2(n_260),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_249),
.B2(n_250),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_250),
.C(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_253),
.C(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_264),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_282),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_276),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_276),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_271),
.C(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_278),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_280),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_296),
.B(n_299),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_286),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_300),
.B2(n_301),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_295),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_295),
.C(n_301),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B(n_294),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_305),
.C(n_315),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_305),
.B1(n_306),
.B2(n_330),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_294),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_317),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_317),
.Y(n_332)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_310),
.C(n_312),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_314),
.B1(n_319),
.B2(n_323),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_323),
.C(n_324),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_316),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_324),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);


endmodule