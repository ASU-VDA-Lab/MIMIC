module fake_jpeg_17117_n_289 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_27),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_16),
.C(n_28),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_37),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_35),
.B1(n_14),
.B2(n_33),
.Y(n_58)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_25),
.Y(n_64)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_33),
.B1(n_17),
.B2(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_58),
.B1(n_67),
.B2(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_62),
.B(n_64),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_43),
.B(n_41),
.C(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_36),
.B1(n_35),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_18),
.B1(n_21),
.B2(n_51),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_40),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_35),
.B1(n_21),
.B2(n_23),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_78),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_42),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_103),
.B(n_71),
.Y(n_107)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_63),
.B1(n_39),
.B2(n_45),
.Y(n_129)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_43),
.B1(n_54),
.B2(n_45),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_101),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_0),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_97),
.Y(n_139)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_111),
.Y(n_156)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_67),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_73),
.B1(n_69),
.B2(n_54),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_60),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_61),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_73),
.B1(n_95),
.B2(n_81),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_57),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_63),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_100),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_90),
.B(n_104),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_105),
.B(n_20),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_87),
.B1(n_79),
.B2(n_92),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_157),
.B1(n_29),
.B2(n_23),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_109),
.B1(n_110),
.B2(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_143),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_145),
.C(n_148),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_94),
.B(n_81),
.C(n_102),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_53),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_30),
.C(n_40),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_122),
.C(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_20),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_18),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_115),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_89),
.B1(n_29),
.B2(n_23),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_120),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_161),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_151),
.B(n_140),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_183),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_172),
.B(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_109),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_77),
.B(n_89),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_111),
.B1(n_22),
.B2(n_29),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_175),
.B1(n_187),
.B2(n_142),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_139),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_20),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_22),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_134),
.B(n_22),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_189),
.A2(n_197),
.B1(n_203),
.B2(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_204),
.C(n_206),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_133),
.C(n_148),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_181),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_144),
.B1(n_131),
.B2(n_150),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_207),
.Y(n_219)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_145),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_142),
.C(n_132),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_157),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_212),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_159),
.B1(n_164),
.B2(n_171),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_210),
.B1(n_165),
.B2(n_28),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_169),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_192),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_168),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_160),
.B1(n_183),
.B2(n_174),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_208),
.B1(n_189),
.B2(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_225),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_164),
.B1(n_175),
.B2(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_224),
.A2(n_228),
.B1(n_201),
.B2(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_1),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_191),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_176),
.C(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_236),
.B1(n_230),
.B2(n_237),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_233),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_237),
.C(n_242),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_165),
.B1(n_210),
.B2(n_134),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_214),
.B(n_9),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_77),
.C(n_28),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_217),
.C(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_246),
.C(n_248),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_211),
.C(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_218),
.C(n_226),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_222),
.C(n_77),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_222),
.C(n_20),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_3),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_8),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_231),
.B1(n_232),
.B2(n_3),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_244),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_9),
.B1(n_4),
.B2(n_6),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_9),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_252),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_3),
.C(n_4),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_270),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_6),
.B(n_7),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_271),
.B1(n_265),
.B2(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_278),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_264),
.B(n_257),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_274),
.B(n_275),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_263),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_281),
.A2(n_276),
.B(n_268),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_282),
.B(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_284),
.B(n_11),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_283),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_13),
.C(n_11),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_12),
.Y(n_289)
);


endmodule