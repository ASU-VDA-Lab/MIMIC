module real_jpeg_30306_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_1),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_1),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_1),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_1),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_2),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_6),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_9),
.B(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_11),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_30),
.Y(n_139)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_14),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_33),
.Y(n_32)
);

AND2x4_ASAP7_75t_SL g92 ( 
.A(n_15),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_15),
.B(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_15),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_142),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_19),
.B(n_122),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_64),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_32),
.C(n_36),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_23),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_129)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_31),
.Y(n_183)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_31),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_32),
.B(n_36),
.Y(n_127)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_49),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_48),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_57),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_106),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_82),
.C(n_95),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_71),
.C(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_95),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.C(n_92),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_84),
.B1(n_92),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_88),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_92),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_101),
.Y(n_109)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_124),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_128),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.C(n_133),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2x2_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_138),
.Y(n_222)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_170),
.B(n_238),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_167),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_145),
.B(n_167),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_163),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.C(n_159),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_150),
.B1(n_159),
.B2(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_188),
.B(n_237),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_172),
.B(n_186),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_184),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_176),
.B1(n_184),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_203),
.B(n_236),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_196),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_192),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_196),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_229),
.B(n_235),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_224),
.B(n_228),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_214),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_223),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);


endmodule