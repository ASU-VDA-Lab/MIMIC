module fake_jpeg_24322_n_284 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_17),
.B1(n_27),
.B2(n_23),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_23),
.B1(n_14),
.B2(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_14),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_7),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_73),
.B1(n_30),
.B2(n_43),
.Y(n_104)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_34),
.B(n_37),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_37),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_38),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_81),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_36),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_90),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_30),
.B1(n_43),
.B2(n_41),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_97),
.B1(n_43),
.B2(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_30),
.A3(n_59),
.B1(n_38),
.B2(n_36),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_74),
.B(n_49),
.Y(n_107)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_71),
.B1(n_59),
.B2(n_56),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_67),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_81),
.B1(n_77),
.B2(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_49),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_65),
.B(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_48),
.B1(n_44),
.B2(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_35),
.B(n_37),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_112),
.B1(n_92),
.B2(n_101),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_127),
.B(n_129),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_81),
.B1(n_77),
.B2(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_114),
.B1(n_122),
.B2(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_36),
.B1(n_38),
.B2(n_48),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_119),
.B1(n_126),
.B2(n_83),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_82),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_98),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_36),
.B1(n_59),
.B2(n_71),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_29),
.B1(n_25),
.B2(n_19),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_57),
.B1(n_37),
.B2(n_35),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_26),
.B(n_35),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_26),
.B(n_35),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_89),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_136),
.B(n_137),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_102),
.B(n_103),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_102),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_138),
.A2(n_144),
.B1(n_133),
.B2(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_102),
.B1(n_96),
.B2(n_86),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_143),
.B1(n_148),
.B2(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_145),
.C(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_130),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_83),
.B1(n_91),
.B2(n_90),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_35),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_105),
.B1(n_78),
.B2(n_68),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_153),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_37),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_105),
.B1(n_94),
.B2(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_29),
.B1(n_25),
.B2(n_19),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_118),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_129),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_152),
.B(n_26),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_117),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_16),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_140),
.B1(n_138),
.B2(n_132),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_186),
.B1(n_191),
.B2(n_196),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_132),
.B1(n_153),
.B2(n_106),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_167),
.B1(n_168),
.B2(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_16),
.C(n_1),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_155),
.C(n_158),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_7),
.C(n_12),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

OAI22x1_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_7),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_175),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_159),
.B1(n_161),
.B2(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_184),
.C(n_182),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_174),
.C(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_212),
.C(n_214),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_208),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_163),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_218),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_165),
.C(n_160),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_179),
.C(n_193),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_162),
.C(n_176),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_0),
.C(n_3),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_164),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_183),
.B1(n_186),
.B2(n_156),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_232),
.B1(n_212),
.B2(n_206),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_229),
.C(n_234),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_197),
.C(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_156),
.B1(n_191),
.B2(n_4),
.Y(n_232)
);

BUFx12f_ASAP7_75t_SL g233 ( 
.A(n_213),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_213),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_8),
.C(n_12),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_240),
.B1(n_231),
.B2(n_228),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_202),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_242),
.Y(n_256)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_248),
.Y(n_249)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_246),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_0),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_235),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_240),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_220),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_9),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_3),
.C(n_4),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_238),
.C(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_266),
.C(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_268),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_239),
.CI(n_10),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_6),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_3),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_4),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_272),
.B(n_274),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_11),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_13),
.B(n_5),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_265),
.C(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_266),
.B(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_271),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_279),
.C(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_278),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_5),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_5),
.Y(n_284)
);


endmodule