module fake_aes_9060_n_35 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_13;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx16_ASAP7_75t_R g9 ( .A(n_5), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_7), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_0), .B(n_5), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_10), .B(n_15), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_9), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx1_ASAP7_75t_SL g19 ( .A(n_9), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_14), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
CKINVDCx16_ASAP7_75t_R g24 ( .A(n_19), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_21), .B(n_16), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_21), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx2_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
AOI211xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_26), .B(n_23), .C(n_22), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_23), .B1(n_25), .B2(n_24), .C(n_16), .Y(n_31) );
NAND2x1p5_ASAP7_75t_L g32 ( .A(n_30), .B(n_29), .Y(n_32) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
OAI22xp5_ASAP7_75t_SL g34 ( .A1(n_32), .A2(n_13), .B1(n_12), .B2(n_29), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_33), .B1(n_4), .B2(n_6), .Y(n_35) );
endmodule