module real_aes_8903_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g478 ( .A1(n_0), .A2(n_157), .B(n_479), .C(n_482), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_1), .B(n_473), .Y(n_483) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g155 ( .A(n_3), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_4), .B(n_158), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_5), .A2(n_468), .B(n_541), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_6), .A2(n_105), .B1(n_430), .B2(n_438), .C1(n_441), .C2(n_745), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_6), .A2(n_78), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_6), .Y(n_116) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_6), .A2(n_180), .B(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_7), .A2(n_40), .B1(n_145), .B2(n_203), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_8), .A2(n_9), .B1(n_736), .B2(n_737), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_8), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_9), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_10), .B(n_180), .Y(n_188) );
AND2x6_ASAP7_75t_L g160 ( .A(n_11), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_12), .A2(n_160), .B(n_459), .C(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_13), .B(n_41), .Y(n_113) );
INVx1_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
INVx1_ASAP7_75t_L g136 ( .A(n_15), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_16), .B(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_17), .B(n_158), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_18), .B(n_132), .Y(n_190) );
AO32x2_ASAP7_75t_L g241 ( .A1(n_19), .A2(n_131), .A3(n_174), .B1(n_180), .B2(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_20), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_20), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_21), .A2(n_32), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_21), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_22), .B(n_145), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_23), .B(n_132), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_24), .A2(n_57), .B1(n_145), .B2(n_203), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_25), .A2(n_83), .B1(n_141), .B2(n_145), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_26), .B(n_145), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_27), .A2(n_174), .B(n_459), .C(n_490), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_28), .A2(n_174), .B(n_459), .C(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_29), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_30), .A2(n_734), .B1(n_735), .B2(n_738), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_30), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_31), .B(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_32), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_32), .A2(n_122), .B1(n_123), .B2(n_124), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_33), .A2(n_468), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_34), .B(n_176), .Y(n_218) );
INVx2_ASAP7_75t_L g143 ( .A(n_35), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_36), .A2(n_465), .B(n_508), .C(n_509), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_37), .B(n_145), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_38), .B(n_176), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_39), .B(n_225), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_42), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_43), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_44), .B(n_158), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_45), .B(n_468), .Y(n_550) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_46), .A2(n_443), .B1(n_729), .B2(n_730), .C1(n_739), .C2(n_742), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_47), .A2(n_465), .B(n_508), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_48), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_49), .B(n_145), .Y(n_183) );
INVx1_ASAP7_75t_L g480 ( .A(n_50), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_51), .A2(n_92), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g533 ( .A(n_52), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_53), .B(n_145), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_54), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_55), .B(n_468), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_56), .B(n_153), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g194 ( .A1(n_58), .A2(n_62), .B1(n_141), .B2(n_145), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_59), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_60), .B(n_145), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_61), .B(n_145), .Y(n_222) );
INVx1_ASAP7_75t_L g161 ( .A(n_63), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_64), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_65), .B(n_473), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_66), .A2(n_147), .B(n_153), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_67), .B(n_145), .Y(n_156) );
INVx1_ASAP7_75t_L g135 ( .A(n_68), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_69), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_70), .B(n_158), .Y(n_511) );
AO32x2_ASAP7_75t_L g200 ( .A1(n_71), .A2(n_174), .A3(n_180), .B1(n_201), .B2(n_206), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_72), .B(n_159), .Y(n_524) );
INVx1_ASAP7_75t_L g170 ( .A(n_73), .Y(n_170) );
INVx1_ASAP7_75t_L g213 ( .A(n_74), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_75), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_76), .B(n_492), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_77), .A2(n_459), .B(n_461), .C(n_465), .Y(n_458) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_79), .B(n_141), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_80), .Y(n_542) );
INVx1_ASAP7_75t_L g437 ( .A(n_81), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_82), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_84), .B(n_203), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_85), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_86), .B(n_141), .Y(n_217) );
INVx2_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_88), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_89), .B(n_173), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_90), .B(n_141), .Y(n_184) );
OR2x2_ASAP7_75t_L g109 ( .A(n_91), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g446 ( .A(n_91), .B(n_111), .Y(n_446) );
INVx2_ASAP7_75t_L g450 ( .A(n_91), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_93), .A2(n_103), .B1(n_141), .B2(n_142), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_94), .B(n_468), .Y(n_506) );
INVx1_ASAP7_75t_L g510 ( .A(n_95), .Y(n_510) );
INVxp67_ASAP7_75t_L g545 ( .A(n_96), .Y(n_545) );
XNOR2xp5_ASAP7_75t_L g118 ( .A(n_97), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_98), .B(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_99), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g462 ( .A(n_100), .Y(n_462) );
INVx1_ASAP7_75t_L g520 ( .A(n_101), .Y(n_520) );
AND2x2_ASAP7_75t_L g535 ( .A(n_102), .B(n_176), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_114), .B(n_428), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g429 ( .A(n_109), .Y(n_429) );
BUFx2_ASAP7_75t_L g440 ( .A(n_109), .Y(n_440) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_110), .B(n_450), .Y(n_744) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g449 ( .A(n_111), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
XNOR2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B1(n_124), .B2(n_427), .Y(n_119) );
INVx1_ASAP7_75t_L g427 ( .A(n_120), .Y(n_427) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR5x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_318), .C(n_376), .D(n_412), .E(n_419), .Y(n_124) );
NAND3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_264), .C(n_288), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_196), .B1(n_230), .B2(n_235), .C(n_245), .Y(n_126) );
OAI21xp5_ASAP7_75t_SL g398 ( .A1(n_127), .A2(n_399), .B(n_401), .Y(n_398) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_177), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_128), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
INVx2_ASAP7_75t_L g234 ( .A(n_129), .Y(n_234) );
AND2x2_ASAP7_75t_L g247 ( .A(n_129), .B(n_179), .Y(n_247) );
AND2x2_ASAP7_75t_L g301 ( .A(n_129), .B(n_178), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_129), .B(n_164), .Y(n_316) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_162), .Y(n_129) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_130), .A2(n_165), .B(n_175), .Y(n_164) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_131), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_133), .B(n_134), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_151), .B(n_160), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_144), .C(n_147), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_140), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_140), .A2(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
INVx3_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_145), .Y(n_464) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
AND2x6_ASAP7_75t_L g459 ( .A(n_146), .B(n_460), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_147), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_148), .A2(n_216), .B(n_217), .Y(n_215) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g492 ( .A(n_149), .Y(n_492) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
INVx1_ASAP7_75t_L g225 ( .A(n_150), .Y(n_225) );
INVx1_ASAP7_75t_L g460 ( .A(n_150), .Y(n_460) );
AND2x2_ASAP7_75t_L g469 ( .A(n_150), .B(n_154), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_156), .C(n_157), .Y(n_151) );
O2A1O1Ixp5_ASAP7_75t_L g169 ( .A1(n_152), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_152), .A2(n_491), .B(n_493), .Y(n_490) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_157), .A2(n_186), .B(n_187), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_157), .A2(n_173), .B1(n_193), .B2(n_194), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_157), .A2(n_173), .B1(n_243), .B2(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_158), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_158), .A2(n_183), .B(n_184), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_SL g211 ( .A1(n_158), .A2(n_212), .B(n_213), .C(n_214), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_158), .B(n_545), .Y(n_544) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g201 ( .A1(n_159), .A2(n_173), .B1(n_202), .B2(n_205), .Y(n_201) );
BUFx3_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_160), .A2(n_182), .B(n_185), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_211), .B(n_215), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_221), .B(n_226), .Y(n_220) );
INVx4_ASAP7_75t_SL g466 ( .A(n_160), .Y(n_466) );
AND2x4_ASAP7_75t_L g468 ( .A(n_160), .B(n_469), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_160), .B(n_469), .Y(n_521) );
AND2x2_ASAP7_75t_L g334 ( .A(n_163), .B(n_275), .Y(n_334) );
AND2x2_ASAP7_75t_L g367 ( .A(n_163), .B(n_179), .Y(n_367) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OR2x2_ASAP7_75t_L g274 ( .A(n_164), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g287 ( .A(n_164), .B(n_179), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_164), .B(n_275), .Y(n_294) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_164), .Y(n_303) );
AND2x2_ASAP7_75t_L g310 ( .A(n_164), .B(n_178), .Y(n_310) );
INVx1_ASAP7_75t_L g341 ( .A(n_164), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_174), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_172), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g481 ( .A(n_173), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_174), .B(n_192), .C(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_210), .B(n_218), .Y(n_209) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_176), .A2(n_220), .B(n_229), .Y(n_219) );
INVx1_ASAP7_75t_L g498 ( .A(n_176), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_176), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_176), .A2(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g317 ( .A(n_177), .Y(n_317) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_189), .Y(n_177) );
INVx2_ASAP7_75t_L g273 ( .A(n_178), .Y(n_273) );
AND2x2_ASAP7_75t_L g295 ( .A(n_178), .B(n_234), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_178), .B(n_341), .Y(n_346) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_179), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g418 ( .A(n_179), .B(n_382), .Y(n_418) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_188), .Y(n_179) );
INVx4_ASAP7_75t_L g195 ( .A(n_180), .Y(n_195) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_180), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_180), .A2(n_550), .B(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
INVx3_ASAP7_75t_L g333 ( .A(n_189), .Y(n_333) );
OR2x2_ASAP7_75t_L g363 ( .A(n_189), .B(n_364), .Y(n_363) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_189), .B(n_273), .Y(n_389) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx1_ASAP7_75t_L g276 ( .A(n_190), .Y(n_276) );
AO21x1_ASAP7_75t_L g275 ( .A1(n_192), .A2(n_195), .B(n_276), .Y(n_275) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_195), .A2(n_457), .B(n_470), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_195), .B(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g473 ( .A(n_195), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_195), .B(n_514), .Y(n_513) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_195), .A2(n_519), .B(n_526), .Y(n_518) );
AOI33xp33_ASAP7_75t_L g409 ( .A1(n_196), .A2(n_247), .A3(n_261), .B1(n_333), .B2(n_410), .B3(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
OR2x2_ASAP7_75t_L g262 ( .A(n_198), .B(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_198), .B(n_259), .Y(n_321) );
OR2x2_ASAP7_75t_L g374 ( .A(n_198), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g300 ( .A(n_199), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g325 ( .A(n_199), .B(n_207), .Y(n_325) );
AND2x2_ASAP7_75t_L g392 ( .A(n_199), .B(n_237), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_199), .A2(n_292), .B(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
INVx1_ASAP7_75t_L g252 ( .A(n_200), .Y(n_252) );
AND2x2_ASAP7_75t_L g271 ( .A(n_200), .B(n_241), .Y(n_271) );
AND2x2_ASAP7_75t_L g320 ( .A(n_200), .B(n_240), .Y(n_320) );
INVx2_ASAP7_75t_L g482 ( .A(n_204), .Y(n_482) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_204), .Y(n_512) );
INVx1_ASAP7_75t_L g495 ( .A(n_206), .Y(n_495) );
INVx2_ASAP7_75t_SL g362 ( .A(n_207), .Y(n_362) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
INVx2_ASAP7_75t_L g282 ( .A(n_208), .Y(n_282) );
INVx1_ASAP7_75t_L g413 ( .A(n_208), .Y(n_413) );
AND2x2_ASAP7_75t_L g426 ( .A(n_208), .B(n_307), .Y(n_426) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g253 ( .A(n_209), .Y(n_253) );
OR2x2_ASAP7_75t_L g259 ( .A(n_209), .B(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_219), .Y(n_237) );
AND2x2_ASAP7_75t_L g254 ( .A(n_219), .B(n_240), .Y(n_254) );
INVx1_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
INVx1_ASAP7_75t_L g267 ( .A(n_219), .Y(n_267) );
AND2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_241), .Y(n_292) );
INVx2_ASAP7_75t_L g308 ( .A(n_219), .Y(n_308) );
AND2x2_ASAP7_75t_L g401 ( .A(n_219), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_219), .B(n_282), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
INVx1_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_232), .B(n_316), .Y(n_382) );
INVx1_ASAP7_75t_SL g342 ( .A(n_233), .Y(n_342) );
INVx2_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
AND2x2_ASAP7_75t_L g332 ( .A(n_234), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g348 ( .A(n_234), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
INVx1_ASAP7_75t_L g410 ( .A(n_236), .Y(n_410) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g368 ( .A(n_238), .B(n_358), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_238), .A2(n_379), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g281 ( .A(n_239), .B(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
INVx1_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
OR2x2_ASAP7_75t_L g394 ( .A(n_240), .B(n_253), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_240), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g307 ( .A(n_241), .B(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_248), .B1(n_255), .B2(n_257), .Y(n_245) );
OR2x2_ASAP7_75t_L g324 ( .A(n_246), .B(n_274), .Y(n_324) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_247), .A2(n_366), .B1(n_368), .B2(n_369), .C1(n_370), .C2(n_373), .Y(n_365) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g312 ( .A(n_251), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_253), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_253), .Y(n_337) );
AND2x2_ASAP7_75t_L g385 ( .A(n_253), .B(n_254), .Y(n_385) );
INVx1_ASAP7_75t_L g403 ( .A(n_253), .Y(n_403) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g369 ( .A(n_256), .B(n_295), .Y(n_369) );
AND2x2_ASAP7_75t_L g411 ( .A(n_256), .B(n_287), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_258), .B(n_306), .Y(n_393) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_259), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g286 ( .A(n_263), .B(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g354 ( .A(n_263), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B(n_272), .C(n_277), .Y(n_264) );
INVxp67_ASAP7_75t_L g278 ( .A(n_265), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_266), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_266), .B(n_313), .Y(n_408) );
BUFx3_ASAP7_75t_L g372 ( .A(n_267), .Y(n_372) );
INVx1_ASAP7_75t_L g279 ( .A(n_268), .Y(n_279) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g298 ( .A(n_270), .B(n_292), .Y(n_298) );
INVx1_ASAP7_75t_SL g338 ( .A(n_271), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g328 ( .A(n_273), .Y(n_328) );
AND2x2_ASAP7_75t_L g351 ( .A(n_273), .B(n_334), .Y(n_351) );
INVx1_ASAP7_75t_SL g322 ( .A(n_274), .Y(n_322) );
INVx1_ASAP7_75t_L g349 ( .A(n_275), .Y(n_349) );
AOI31xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .A3(n_280), .B(n_283), .Y(n_277) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g370 ( .A(n_281), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g344 ( .A(n_282), .Y(n_344) );
BUFx2_ASAP7_75t_L g358 ( .A(n_282), .Y(n_358) );
AND2x2_ASAP7_75t_L g386 ( .A(n_282), .B(n_307), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g359 ( .A(n_286), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_287), .B(n_354), .Y(n_400) );
AND2x2_ASAP7_75t_L g407 ( .A(n_287), .B(n_333), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_293), .B(n_296), .C(n_311), .Y(n_288) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_293), .A2(n_320), .B1(n_321), .B2(n_322), .C(n_323), .Y(n_319) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g327 ( .A(n_294), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
OAI32xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .A3(n_302), .B1(n_304), .B2(n_309), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_298), .A2(n_351), .B(n_352), .C(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_306), .A2(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g375 ( .A(n_307), .Y(n_375) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_313), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g361 ( .A(n_313), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND4xp25_ASAP7_75t_SL g318 ( .A(n_319), .B(n_331), .C(n_350), .D(n_365), .Y(n_318) );
AND2x2_ASAP7_75t_L g357 ( .A(n_320), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g379 ( .A(n_320), .B(n_372), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_322), .B(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_326), .B2(n_329), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_324), .A2(n_375), .B1(n_406), .B2(n_408), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g412 ( .A1(n_324), .A2(n_413), .B(n_414), .C(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g383 ( .A(n_325), .Y(n_383) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_327), .A2(n_361), .B1(n_378), .B2(n_379), .C1(n_380), .C2(n_383), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_335), .C(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g397 ( .A(n_332), .Y(n_397) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_336), .A2(n_340), .B1(n_343), .B2(n_345), .Y(n_339) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g366 ( .A(n_348), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g424 ( .A(n_351), .Y(n_424) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B1(n_360), .B2(n_363), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_358), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g415 ( .A(n_363), .Y(n_415) );
INVx1_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_369), .Y(n_423) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND5xp2_ASAP7_75t_L g376 ( .A(n_377), .B(n_384), .C(n_398), .D(n_404), .E(n_409), .Y(n_376) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_387), .C(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI31xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .A3(n_394), .B(n_395), .Y(n_390) );
INVx1_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g419 ( .A1(n_406), .A2(n_408), .B1(n_420), .B2(n_423), .C1(n_424), .C2(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g748 ( .A(n_429), .Y(n_748) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_434), .A2(n_435), .B(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g747 ( .A(n_434), .B(n_436), .Y(n_747) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B1(n_448), .B2(n_451), .Y(n_444) );
INVx2_ASAP7_75t_L g740 ( .A(n_445), .Y(n_740) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_447), .A2(n_451), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g741 ( .A(n_448), .Y(n_741) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_637), .C(n_686), .Y(n_451) );
NAND5xp2_ASAP7_75t_L g452 ( .A(n_453), .B(n_571), .C(n_600), .D(n_608), .E(n_623), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_499), .B(n_515), .C(n_555), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_484), .Y(n_454) );
AND2x2_ASAP7_75t_L g566 ( .A(n_455), .B(n_563), .Y(n_566) );
AND2x2_ASAP7_75t_L g599 ( .A(n_455), .B(n_485), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_455), .B(n_503), .Y(n_692) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_472), .Y(n_455) );
INVx2_ASAP7_75t_L g502 ( .A(n_456), .Y(n_502) );
BUFx2_ASAP7_75t_L g666 ( .A(n_456), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_467), .Y(n_457) );
INVx5_ASAP7_75t_L g477 ( .A(n_459), .Y(n_477) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_466), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_466), .A2(n_477), .B(n_542), .C(n_543), .Y(n_541) );
BUFx2_ASAP7_75t_L g488 ( .A(n_468), .Y(n_488) );
AND2x2_ASAP7_75t_L g484 ( .A(n_472), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g564 ( .A(n_472), .Y(n_564) );
AND2x2_ASAP7_75t_L g650 ( .A(n_472), .B(n_563), .Y(n_650) );
AND2x2_ASAP7_75t_L g705 ( .A(n_472), .B(n_502), .Y(n_705) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_483), .Y(n_472) );
INVx2_ASAP7_75t_L g508 ( .A(n_477), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g622 ( .A(n_484), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_484), .B(n_503), .Y(n_669) );
INVx5_ASAP7_75t_L g563 ( .A(n_485), .Y(n_563) );
AND2x4_ASAP7_75t_L g584 ( .A(n_485), .B(n_564), .Y(n_584) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_485), .Y(n_606) );
AND2x2_ASAP7_75t_L g681 ( .A(n_485), .B(n_666), .Y(n_681) );
AND2x2_ASAP7_75t_L g684 ( .A(n_485), .B(n_504), .Y(n_684) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_489), .B(n_495), .Y(n_486) );
INVx2_ASAP7_75t_L g494 ( .A(n_492), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_494), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_494), .A2(n_512), .B(n_533), .C(n_534), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_499), .B(n_564), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_499), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
AND2x2_ASAP7_75t_L g589 ( .A(n_501), .B(n_564), .Y(n_589) );
AND2x2_ASAP7_75t_L g607 ( .A(n_501), .B(n_504), .Y(n_607) );
INVx1_ASAP7_75t_L g627 ( .A(n_501), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_501), .B(n_563), .Y(n_672) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_501), .Y(n_714) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_502), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_503), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_503), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_503), .A2(n_559), .B(n_620), .C(n_622), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_503), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g635 ( .A(n_503), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g639 ( .A(n_503), .B(n_563), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_503), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g654 ( .A(n_503), .B(n_564), .Y(n_654) );
AND2x2_ASAP7_75t_L g704 ( .A(n_503), .B(n_705), .Y(n_704) );
INVx5_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g568 ( .A(n_504), .Y(n_568) );
AND2x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_562), .Y(n_609) );
AND2x2_ASAP7_75t_L g621 ( .A(n_504), .B(n_596), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_504), .B(n_650), .Y(n_668) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_536), .Y(n_515) );
INVx1_ASAP7_75t_L g557 ( .A(n_516), .Y(n_557) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
OR2x2_ASAP7_75t_L g559 ( .A(n_517), .B(n_528), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_517), .B(n_566), .C(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_517), .B(n_538), .Y(n_576) );
OR2x2_ASAP7_75t_L g591 ( .A(n_517), .B(n_579), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_517), .B(n_547), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_517), .B(n_728), .Y(n_727) );
INVx5_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_518), .B(n_538), .Y(n_594) );
AND2x2_ASAP7_75t_L g633 ( .A(n_518), .B(n_548), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_518), .B(n_547), .Y(n_661) );
OR2x2_ASAP7_75t_L g664 ( .A(n_518), .B(n_547), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_522), .Y(n_519) );
INVx5_ASAP7_75t_SL g579 ( .A(n_528), .Y(n_579) );
OR2x2_ASAP7_75t_L g585 ( .A(n_528), .B(n_537), .Y(n_585) );
AND2x2_ASAP7_75t_L g601 ( .A(n_528), .B(n_602), .Y(n_601) );
AOI321xp33_ASAP7_75t_L g608 ( .A1(n_528), .A2(n_609), .A3(n_610), .B1(n_611), .B2(n_617), .C(n_619), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_528), .B(n_536), .Y(n_618) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_528), .Y(n_631) );
OR2x2_ASAP7_75t_L g678 ( .A(n_528), .B(n_576), .Y(n_678) );
AND2x2_ASAP7_75t_L g700 ( .A(n_528), .B(n_597), .Y(n_700) );
AND2x2_ASAP7_75t_L g719 ( .A(n_528), .B(n_538), .Y(n_719) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_535), .Y(n_528) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_538), .B(n_547), .Y(n_560) );
AND2x2_ASAP7_75t_L g569 ( .A(n_538), .B(n_570), .Y(n_569) );
INVx3_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_538), .B(n_597), .Y(n_602) );
INVxp67_ASAP7_75t_L g632 ( .A(n_538), .Y(n_632) );
OR2x2_ASAP7_75t_L g674 ( .A(n_538), .B(n_579), .Y(n_674) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_546), .Y(n_538) );
OR2x2_ASAP7_75t_L g556 ( .A(n_547), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g570 ( .A(n_547), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_547), .B(n_559), .Y(n_603) );
AND2x2_ASAP7_75t_L g652 ( .A(n_547), .B(n_596), .Y(n_652) );
AND2x2_ASAP7_75t_L g690 ( .A(n_547), .B(n_579), .Y(n_690) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_548), .B(n_579), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .B(n_561), .C(n_565), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_556), .A2(n_558), .B1(n_683), .B2(n_685), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_558), .A2(n_581), .B1(n_636), .B2(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_SL g710 ( .A(n_559), .Y(n_710) );
INVx1_ASAP7_75t_SL g610 ( .A(n_560), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_562), .B(n_582), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g623 ( .A1(n_562), .A2(n_603), .B1(n_610), .B2(n_624), .C1(n_628), .C2(n_634), .Y(n_623) );
AND2x2_ASAP7_75t_L g713 ( .A(n_562), .B(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g588 ( .A(n_563), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_563), .B(n_583), .Y(n_658) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_563), .Y(n_695) );
AND2x2_ASAP7_75t_L g698 ( .A(n_563), .B(n_607), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_563), .B(n_714), .Y(n_724) );
INVx1_ASAP7_75t_L g615 ( .A(n_564), .Y(n_615) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_564), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g706 ( .A1(n_566), .A2(n_707), .B(n_708), .C(n_711), .Y(n_706) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_568), .B(n_630), .C(n_633), .Y(n_629) );
OR2x2_ASAP7_75t_L g657 ( .A(n_568), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_568), .B(n_584), .Y(n_685) );
OR2x2_ASAP7_75t_L g590 ( .A(n_570), .B(n_591), .Y(n_590) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_580), .C(n_592), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_573), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g679 ( .A(n_574), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_575), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g593 ( .A(n_578), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_579), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g647 ( .A(n_579), .B(n_597), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_579), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_579), .B(n_596), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B1(n_586), .B2(n_590), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_582), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_584), .B(n_626), .Y(n_625) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_585), .A2(n_649), .B1(n_651), .B2(n_653), .C(n_655), .Y(n_648) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g703 ( .A(n_588), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g716 ( .A(n_588), .B(n_705), .Y(n_716) );
INVx1_ASAP7_75t_L g636 ( .A(n_589), .Y(n_636) );
INVx1_ASAP7_75t_L g707 ( .A(n_590), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_591), .A2(n_674), .B(n_697), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B(n_598), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_603), .B(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g640 ( .A(n_601), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_602), .A2(n_688), .B1(n_691), .B2(n_693), .C(n_696), .Y(n_687) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_610), .A2(n_700), .B1(n_701), .B2(n_703), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g676 ( .A(n_612), .Y(n_676) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2xp67_ASAP7_75t_SL g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g680 ( .A(n_616), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g645 ( .A(n_621), .Y(n_645) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_626), .B(n_650), .Y(n_702) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_632), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g718 ( .A(n_633), .B(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g725 ( .A(n_633), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI211xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_640), .B(n_641), .C(n_675), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B(n_648), .C(n_667), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g728 ( .A(n_652), .Y(n_728) );
AND2x2_ASAP7_75t_L g665 ( .A(n_654), .B(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_663), .B2(n_665), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OR2x2_ASAP7_75t_L g673 ( .A(n_661), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g726 ( .A(n_662), .Y(n_726) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI31xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .A3(n_670), .B(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_679), .C(n_682), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
NAND5xp2_ASAP7_75t_L g686 ( .A(n_687), .B(n_699), .C(n_706), .D(n_720), .E(n_723), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_698), .A2(n_724), .B1(n_725), .B2(n_727), .Y(n_723) );
INVx1_ASAP7_75t_SL g722 ( .A(n_700), .Y(n_722) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B(n_717), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
CKINVDCx14_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx3_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
NAND2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
endmodule