module fake_jpeg_13818_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_24),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_50),
.B1(n_57),
.B2(n_55),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_64),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_1),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_67),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_72),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_53),
.B1(n_45),
.B2(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_7),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_52),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_63),
.B1(n_65),
.B2(n_4),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_22),
.B1(n_40),
.B2(n_39),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_95),
.Y(n_103)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_9),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_9),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_11),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_69),
.B(n_79),
.C(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_10),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_111),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_10),
.B(n_11),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_28),
.C(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_117),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_17),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_88),
.Y(n_113)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_18),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_19),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_103),
.C(n_112),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_35),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_114),
.B(n_101),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_107),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_113),
.B(n_110),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_126),
.B1(n_105),
.B2(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_131),
.B1(n_102),
.B2(n_125),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_102),
.A3(n_119),
.B1(n_124),
.B2(n_120),
.C1(n_106),
.C2(n_41),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_119),
.C(n_36),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_37),
.Y(n_139)
);


endmodule