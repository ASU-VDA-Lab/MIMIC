module fake_jpeg_20692_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_23),
.Y(n_46)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_50),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_33),
.B1(n_27),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_41),
.B1(n_42),
.B2(n_38),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_25),
.B1(n_36),
.B2(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_20),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_30),
.B1(n_31),
.B2(n_26),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_38),
.B1(n_42),
.B2(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_61),
.B(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_67),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_38),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_71),
.B(n_74),
.Y(n_104)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_37),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NAND2x1p5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NAND2x1_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_36),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_81),
.B1(n_47),
.B2(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_12),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_12),
.Y(n_77)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_77),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_36),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_83),
.B1(n_86),
.B2(n_44),
.Y(n_113)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_73),
.B1(n_87),
.B2(n_47),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_41),
.C(n_43),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_44),
.C(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_26),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_38),
.B(n_42),
.C(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_109),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_38),
.B1(n_42),
.B2(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_98),
.B1(n_116),
.B2(n_103),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_70),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_43),
.B1(n_39),
.B2(n_35),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_43),
.B1(n_39),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_114),
.B1(n_85),
.B2(n_69),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_26),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_90),
.C(n_92),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_43),
.B1(n_39),
.B2(n_35),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_80),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_22),
.B1(n_32),
.B2(n_24),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_83),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_86),
.B1(n_65),
.B2(n_74),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_129),
.Y(n_167)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_125),
.B(n_133),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_86),
.B(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_138),
.B(n_97),
.Y(n_174)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_132),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_62),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_86),
.B(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_10),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_92),
.B1(n_69),
.B2(n_62),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_35),
.B1(n_39),
.B2(n_79),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_15),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_144),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_39),
.B1(n_35),
.B2(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_35),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_72),
.B1(n_64),
.B2(n_22),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_147),
.B1(n_106),
.B2(n_98),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_117),
.B1(n_96),
.B2(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_20),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_108),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_175),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_159),
.B1(n_161),
.B2(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_104),
.C(n_103),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_158),
.C(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_94),
.C(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_100),
.B1(n_98),
.B2(n_111),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_111),
.B1(n_107),
.B2(n_110),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_123),
.C(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_142),
.B(n_22),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_0),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_110),
.C(n_93),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_93),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_32),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_210),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_158),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_198),
.B(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_131),
.B1(n_143),
.B2(n_135),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_201),
.B1(n_203),
.B2(n_157),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_133),
.B(n_135),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_135),
.B1(n_125),
.B2(n_124),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_212),
.B1(n_156),
.B2(n_167),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_124),
.B1(n_127),
.B2(n_137),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_183),
.B1(n_184),
.B2(n_163),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_0),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_176),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_17),
.B1(n_16),
.B2(n_24),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_170),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_179),
.A2(n_0),
.B(n_1),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_1),
.B(n_2),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_152),
.C(n_155),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_189),
.C(n_209),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_172),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

XOR2x2_ASAP7_75t_SL g256 ( 
.A(n_221),
.B(n_4),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_180),
.B1(n_171),
.B2(n_165),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_229),
.B1(n_234),
.B2(n_235),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_17),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_16),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_197),
.B1(n_201),
.B2(n_208),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_240),
.B1(n_187),
.B2(n_214),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_3),
.B(n_4),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_196),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_191),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_244),
.B(n_246),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_215),
.C(n_189),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_253),
.C(n_232),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_195),
.B1(n_198),
.B2(n_185),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_229),
.B1(n_235),
.B2(n_219),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_202),
.B(n_188),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_239),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_212),
.C(n_213),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_216),
.B1(n_222),
.B2(n_234),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_10),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_226),
.Y(n_261)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_7),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_258),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_259),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_263),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_245),
.C(n_254),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_247),
.C(n_233),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_271),
.C(n_250),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_220),
.C(n_255),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_216),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_241),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_227),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_277),
.B1(n_242),
.B2(n_273),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_277),
.B1(n_242),
.B2(n_256),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

INVxp33_ASAP7_75t_SL g279 ( 
.A(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_280),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_249),
.C(n_245),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_222),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_283),
.Y(n_292)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_238),
.C(n_221),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_299),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_264),
.B(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_266),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_272),
.B1(n_238),
.B2(n_240),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_279),
.B(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_284),
.B1(n_288),
.B2(n_280),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_261),
.B1(n_10),
.B2(n_11),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_11),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_15),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_312),
.B(n_13),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_298),
.C(n_11),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_307),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_5),
.B(n_6),
.Y(n_320)
);

NOR4xp25_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_309),
.C(n_305),
.D(n_13),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_319),
.A2(n_320),
.B(n_316),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_321),
.B(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_5),
.Y(n_326)
);


endmodule