module fake_jpeg_9826_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_55),
.B(n_63),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_25),
.B1(n_42),
.B2(n_51),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_24),
.B1(n_31),
.B2(n_34),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_25),
.B1(n_30),
.B2(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_74),
.B1(n_23),
.B2(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_17),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_60),
.B(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_75),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_33),
.B1(n_21),
.B2(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_26),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_20),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_91),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_24),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_101),
.C(n_105),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_93)
);

OAI22x1_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_104),
.B1(n_23),
.B2(n_6),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_96),
.B1(n_112),
.B2(n_90),
.Y(n_140)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_32),
.C(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_17),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_112),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_33),
.B1(n_34),
.B2(n_12),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_56),
.B(n_32),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_29),
.B1(n_26),
.B2(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_75),
.B(n_22),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_118),
.Y(n_136)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_115),
.Y(n_143)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_23),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_23),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

OR2x2_ASAP7_75t_SL g126 ( 
.A(n_54),
.B(n_32),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_32),
.C(n_29),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_26),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_73),
.B1(n_80),
.B2(n_69),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_151),
.B1(n_157),
.B2(n_94),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_97),
.B1(n_106),
.B2(n_127),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_80),
.C(n_69),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_154),
.C(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_147),
.B1(n_153),
.B2(n_156),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_73),
.B1(n_54),
.B2(n_32),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_116),
.B(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_98),
.A2(n_90),
.B1(n_113),
.B2(n_120),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_29),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_123),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_108),
.A2(n_29),
.B1(n_26),
.B2(n_9),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_89),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_164),
.Y(n_195)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_89),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_183),
.B1(n_184),
.B2(n_97),
.Y(n_207)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_166),
.B(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_105),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_105),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_126),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_192),
.B(n_129),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_105),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_175),
.C(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_151),
.B1(n_132),
.B2(n_130),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_180),
.B1(n_131),
.B2(n_142),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_124),
.C(n_95),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_87),
.Y(n_179)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_88),
.B1(n_91),
.B2(n_103),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_87),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_185),
.Y(n_203)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g197 ( 
.A(n_187),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_193),
.B1(n_97),
.B2(n_92),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_146),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_12),
.B(n_11),
.C(n_9),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_12),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_123),
.B(n_107),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_199),
.C(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_134),
.B1(n_137),
.B2(n_144),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_196),
.A2(n_206),
.B1(n_208),
.B2(n_216),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_168),
.B(n_179),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_146),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_192),
.B1(n_166),
.B2(n_191),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_218),
.B1(n_220),
.B2(n_222),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_157),
.B1(n_139),
.B2(n_131),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_211),
.B1(n_172),
.B2(n_160),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_141),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_222),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_150),
.B(n_146),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_225),
.C(n_8),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_221),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_187),
.B1(n_161),
.B2(n_164),
.Y(n_216)
);

XNOR2x2_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_13),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_115),
.B1(n_114),
.B2(n_122),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_170),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_92),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_226),
.B(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_186),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_232),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_252),
.B1(n_217),
.B2(n_211),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_238),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_235),
.B(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_197),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_240),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_172),
.B1(n_183),
.B2(n_169),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_250),
.B1(n_199),
.B2(n_219),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_197),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_14),
.Y(n_243)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_230),
.C(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_0),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_195),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_250),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_251),
.B1(n_252),
.B2(n_238),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_194),
.B1(n_213),
.B2(n_204),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_271),
.B1(n_229),
.B2(n_234),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_205),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_239),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.C(n_269),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_204),
.C(n_225),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_240),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_201),
.C(n_223),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_219),
.B(n_215),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_201),
.B1(n_212),
.B2(n_203),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_277),
.B(n_282),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_253),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_265),
.C(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_237),
.C(n_251),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_249),
.C(n_233),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_241),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_289),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_288),
.B(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_261),
.B(n_227),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_290),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_257),
.CI(n_255),
.CON(n_292),
.SN(n_292)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_258),
.B(n_257),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_275),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_273),
.B1(n_268),
.B2(n_232),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_305),
.B1(n_302),
.B2(n_294),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_SL g304 ( 
.A1(n_279),
.A2(n_231),
.A3(n_256),
.B1(n_264),
.B2(n_261),
.C1(n_268),
.C2(n_273),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_284),
.Y(n_310)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_310),
.B(n_298),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_281),
.B1(n_275),
.B2(n_226),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_293),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_274),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_300),
.C(n_301),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_295),
.B(n_297),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_274),
.B1(n_1),
.B2(n_2),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_312),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_301),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_323),
.C(n_314),
.Y(n_330)
);

INVx11_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_292),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_326),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_323),
.A2(n_300),
.B(n_309),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_330),
.B(n_321),
.Y(n_333)
);

OAI321xp33_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_329),
.A3(n_318),
.B1(n_319),
.B2(n_317),
.C(n_306),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_316),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_322),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_335),
.B(n_6),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_325),
.B1(n_306),
.B2(n_313),
.Y(n_335)
);

AOI311xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.A3(n_8),
.B(n_4),
.C(n_5),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_0),
.B(n_3),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_0),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_3),
.C(n_4),
.Y(n_340)
);


endmodule