module fake_netlist_6_207_n_1909 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1909);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1909;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_474;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_44),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_23),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_79),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_122),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_110),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_50),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_72),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_43),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_24),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_40),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_101),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_90),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_78),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_38),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_62),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_16),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_152),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_28),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_44),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_111),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_61),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_82),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_63),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_126),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_62),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_116),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_74),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_86),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_28),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_63),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_37),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_89),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_39),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_53),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_77),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_76),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_150),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_129),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_45),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_102),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_124),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_43),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_38),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_34),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_105),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_19),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_145),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_112),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_23),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_31),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_147),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_155),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_133),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_16),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_115),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_47),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_56),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_20),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_26),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_32),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_0),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_3),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_48),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_108),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_100),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_113),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_60),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_120),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_18),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_50),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_12),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_80),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_64),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_93),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_29),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_168),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_162),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_39),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_123),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_159),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_104),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_69),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_169),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_26),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_91),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_65),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_20),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_118),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_84),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_10),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_109),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_56),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_3),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_33),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_73),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_144),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_42),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_36),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_51),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_59),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_103),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_134),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_96),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_153),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_11),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_61),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_8),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_57),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_95),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_87),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_167),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_35),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_30),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_27),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_19),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_22),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_136),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_161),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_57),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_21),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_259),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_266),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_179),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_173),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_260),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_177),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_231),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_231),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_178),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_231),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_182),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_261),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_261),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_182),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_261),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_269),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_172),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_179),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_174),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_240),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_240),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_197),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_240),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_180),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_239),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_246),
.B(n_0),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_185),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_242),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_171),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_171),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_257),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_181),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_181),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_183),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_187),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_266),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_308),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_179),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_183),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_189),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_260),
.B(n_2),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_336),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_196),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_196),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_205),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_190),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_205),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_192),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_246),
.B(n_2),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_222),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_222),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_198),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_202),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_308),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_225),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_246),
.B(n_4),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_225),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_203),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_211),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_220),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_175),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_226),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_175),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_322),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_228),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_228),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_229),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_234),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_201),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_346),
.B(n_246),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_346),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_340),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_329),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_201),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_363),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_389),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_356),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_344),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_344),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_389),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_417),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_375),
.B(n_338),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_348),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_R g450 ( 
.A(n_393),
.B(n_338),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_352),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_342),
.A2(n_290),
.B1(n_310),
.B2(n_224),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_366),
.B(n_329),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_362),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_402),
.A2(n_215),
.B(n_204),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_367),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_353),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_353),
.A2(n_250),
.B(n_235),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_355),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_402),
.A2(n_215),
.B(n_204),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_357),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_367),
.B(n_236),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_358),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_409),
.B(n_201),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_358),
.B(n_204),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_360),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_369),
.B(n_238),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_360),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_369),
.B(n_337),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_372),
.B(n_337),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_372),
.B(n_176),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_374),
.B(n_337),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_414),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_443),
.B(n_409),
.C(n_394),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_457),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_347),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_351),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_464),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g507 ( 
.A(n_428),
.B(n_395),
.C(n_349),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_448),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_478),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_478),
.A2(n_341),
.B1(n_370),
.B2(n_364),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_448),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_460),
.B(n_431),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_428),
.B(n_416),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_354),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_L g519 ( 
.A(n_464),
.B(n_378),
.C(n_374),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

BUFx8_ASAP7_75t_SL g522 ( 
.A(n_457),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_424),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_478),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_424),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_424),
.Y(n_529)
);

CKINVDCx6p67_ASAP7_75t_R g530 ( 
.A(n_498),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_450),
.A2(n_268),
.B1(n_319),
.B2(n_237),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_464),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_436),
.A2(n_387),
.B1(n_388),
.B2(n_342),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_471),
.B(n_371),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_424),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_450),
.A2(n_230),
.B1(n_252),
.B2(n_224),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_376),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_436),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_424),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_453),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_483),
.B(n_416),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_431),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_453),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_425),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_426),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_483),
.B(n_386),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_426),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_498),
.B(n_206),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_427),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_458),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_460),
.B(n_392),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_431),
.A2(n_494),
.B1(n_496),
.B2(n_493),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_427),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_461),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_493),
.B(n_399),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_429),
.Y(n_559)
);

BUFx12f_ASAP7_75t_L g560 ( 
.A(n_441),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_456),
.A2(n_407),
.B1(n_387),
.B2(n_388),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_425),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_425),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_495),
.B(n_215),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_493),
.B(n_295),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_460),
.B(n_407),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_430),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_494),
.A2(n_361),
.B1(n_391),
.B2(n_176),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_456),
.B(n_295),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_425),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_425),
.Y(n_576)
);

AO21x2_ASAP7_75t_L g577 ( 
.A1(n_458),
.A2(n_468),
.B(n_209),
.Y(n_577)
);

INVx6_ASAP7_75t_L g578 ( 
.A(n_447),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_494),
.B(n_401),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_437),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_439),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_425),
.Y(n_582)
);

OAI21xp33_ASAP7_75t_SL g583 ( 
.A1(n_458),
.A2(n_250),
.B(n_235),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_468),
.B(n_295),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_425),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_447),
.B(n_405),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_455),
.B(n_406),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_432),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_439),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_442),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_432),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_432),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_432),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_468),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_496),
.A2(n_264),
.B1(n_382),
.B2(n_270),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_442),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_455),
.B(n_411),
.Y(n_597)
);

AND3x2_ASAP7_75t_L g598 ( 
.A(n_496),
.B(n_209),
.C(n_188),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_432),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_495),
.B(n_207),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_432),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_438),
.B(n_378),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_444),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_432),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_444),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_497),
.B(n_451),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_432),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_447),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_447),
.B(n_412),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_449),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_449),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_489),
.B(n_413),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_L g613 ( 
.A1(n_451),
.A2(n_230),
.B1(n_252),
.B2(n_276),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_459),
.A2(n_276),
.B1(n_339),
.B2(n_335),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_433),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_459),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_447),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_497),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_447),
.B(n_415),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_433),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_433),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_497),
.Y(n_622)
);

AO21x2_ASAP7_75t_L g623 ( 
.A1(n_438),
.A2(n_210),
.B(n_188),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_438),
.B(n_210),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_489),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_462),
.B(n_465),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_447),
.B(n_420),
.Y(n_627)
);

INVxp67_ASAP7_75t_SL g628 ( 
.A(n_433),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_489),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_433),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_447),
.B(n_421),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_447),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_489),
.A2(n_265),
.B1(n_334),
.B2(n_331),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_462),
.B(n_216),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_446),
.B(n_206),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_461),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_433),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_465),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_433),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_489),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_433),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_446),
.B(n_216),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_403),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_446),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_434),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_472),
.B(n_403),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_434),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_472),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_466),
.B(n_214),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_534),
.B(n_491),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_549),
.B(n_491),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_513),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_626),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_555),
.B(n_491),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_551),
.B(n_368),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_551),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_612),
.B(n_491),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_543),
.B(n_491),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_505),
.B(n_373),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_506),
.A2(n_223),
.B(n_219),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_543),
.B(n_473),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_513),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_516),
.B(n_492),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_516),
.B(n_492),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_512),
.B(n_207),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_513),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_528),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_579),
.A2(n_377),
.B1(n_379),
.B2(n_255),
.Y(n_670)
);

BUFx6f_ASAP7_75t_SL g671 ( 
.A(n_521),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_499),
.B(n_473),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_618),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_650),
.B(n_492),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_567),
.B(n_207),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_506),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_512),
.B(n_207),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

OAI221xp5_ASAP7_75t_L g682 ( 
.A1(n_633),
.A2(n_272),
.B1(n_270),
.B2(n_331),
.C(n_265),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_650),
.B(n_492),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_618),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_539),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_539),
.B(n_475),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_566),
.B(n_492),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_566),
.B(n_492),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_541),
.B(n_475),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_510),
.A2(n_532),
.B(n_583),
.C(n_519),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_214),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_606),
.B(n_476),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_524),
.B(n_207),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_606),
.B(n_476),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_542),
.B(n_255),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_644),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_648),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_616),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_207),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_566),
.B(n_492),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_647),
.B(n_492),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_524),
.B(n_233),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_647),
.B(n_466),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_648),
.B(n_479),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_SL g706 ( 
.A(n_561),
.B(n_184),
.C(n_170),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_622),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_544),
.B(n_479),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_622),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_645),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_616),
.B(n_233),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_558),
.A2(n_517),
.B1(n_499),
.B2(n_504),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_404),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_510),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_554),
.B(n_638),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_647),
.B(n_466),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_567),
.B(n_233),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_616),
.B(n_233),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_518),
.A2(n_191),
.B1(n_251),
.B2(n_298),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_567),
.A2(n_292),
.B1(n_291),
.B2(n_289),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_532),
.B(n_466),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_568),
.B(n_186),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_600),
.B(n_466),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_600),
.B(n_470),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_548),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_548),
.Y(n_726)
);

NOR3xp33_ASAP7_75t_L g727 ( 
.A(n_587),
.B(n_597),
.C(n_533),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_550),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_568),
.B(n_193),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_SL g730 ( 
.A1(n_557),
.A2(n_244),
.B1(n_199),
.B2(n_208),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_616),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_507),
.B(n_194),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_645),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_553),
.B(n_233),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_550),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_552),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_557),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_507),
.B(n_200),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_625),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_553),
.B(n_233),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_552),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_553),
.B(n_241),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_636),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_531),
.B(n_212),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_634),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_600),
.B(n_470),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_556),
.B(n_470),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_594),
.B(n_247),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_634),
.B(n_480),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_522),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_556),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_531),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_559),
.B(n_563),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_559),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_594),
.B(n_254),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_536),
.B(n_213),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_563),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_569),
.B(n_470),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_594),
.B(n_258),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_569),
.B(n_470),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_570),
.B(n_487),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_570),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_567),
.A2(n_273),
.B1(n_262),
.B2(n_263),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_536),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_572),
.B(n_487),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_636),
.Y(n_766)
);

OR2x2_ASAP7_75t_SL g767 ( 
.A(n_613),
.B(n_272),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_572),
.B(n_487),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_580),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_634),
.B(n_480),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_514),
.B(n_217),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_634),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_580),
.B(n_487),
.Y(n_773)
);

NOR2x1p5_ASAP7_75t_L g774 ( 
.A(n_530),
.B(n_218),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_581),
.B(n_490),
.Y(n_775)
);

INVx8_ASAP7_75t_L g776 ( 
.A(n_567),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_581),
.B(n_490),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_614),
.B(n_221),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_567),
.A2(n_275),
.B1(n_277),
.B2(n_279),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_503),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_589),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_560),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_589),
.B(n_490),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_590),
.B(n_490),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_625),
.B(n_281),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_590),
.B(n_219),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_596),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_596),
.B(n_223),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_614),
.Y(n_789)
);

BUFx6f_ASAP7_75t_SL g790 ( 
.A(n_521),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_603),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_603),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_605),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_625),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_571),
.B(n_484),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_484),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_605),
.B(n_610),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_610),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_611),
.B(n_227),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_611),
.B(n_227),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_583),
.A2(n_488),
.B(n_485),
.C(n_274),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_629),
.B(n_243),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_635),
.B(n_232),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_629),
.B(n_243),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_640),
.B(n_294),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_509),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_602),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_509),
.Y(n_809)
);

NOR2x1p5_ASAP7_75t_L g810 ( 
.A(n_530),
.B(n_245),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_640),
.B(n_609),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_640),
.B(n_282),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_602),
.Y(n_813)
);

O2A1O1Ixp5_ASAP7_75t_L g814 ( 
.A1(n_651),
.A2(n_288),
.B(n_292),
.C(n_291),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_509),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_519),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_547),
.B(n_296),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_619),
.B(n_248),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_567),
.B(n_282),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_599),
.B(n_286),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_623),
.B(n_485),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_634),
.A2(n_288),
.B1(n_289),
.B2(n_286),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_624),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_662),
.A2(n_628),
.B(n_584),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_691),
.B(n_586),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_675),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_794),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_752),
.B(n_643),
.C(n_624),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_652),
.A2(n_584),
.B(n_631),
.Y(n_829)
);

BUFx12f_ASAP7_75t_L g830 ( 
.A(n_782),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_808),
.B(n_574),
.Y(n_831)
);

NAND2x1p5_ASAP7_75t_L g832 ( 
.A(n_668),
.B(n_547),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_653),
.A2(n_584),
.B(n_608),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_813),
.B(n_823),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_661),
.B(n_643),
.C(n_627),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_685),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_817),
.A2(n_584),
.B(n_525),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_690),
.A2(n_574),
.B(n_623),
.C(n_584),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_659),
.A2(n_617),
.B(n_608),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_677),
.A2(n_632),
.B(n_617),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_677),
.A2(n_632),
.B(n_547),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_782),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_700),
.A2(n_547),
.B(n_577),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_690),
.A2(n_525),
.B(n_523),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_663),
.B(n_692),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_794),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_663),
.B(n_574),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_700),
.A2(n_577),
.B(n_525),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_692),
.B(n_694),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_737),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_750),
.B(n_560),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_695),
.A2(n_738),
.B(n_732),
.C(n_771),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_655),
.B(n_598),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_715),
.B(n_560),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_717),
.A2(n_577),
.B(n_526),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_717),
.A2(n_688),
.B(n_687),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_794),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_694),
.B(n_574),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_678),
.B(n_574),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_714),
.B(n_623),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_778),
.A2(n_595),
.B(n_646),
.C(n_641),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_701),
.A2(n_577),
.B(n_526),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_803),
.B(n_540),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_675),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_776),
.A2(n_526),
.B(n_523),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_684),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_540),
.B1(n_575),
.B2(n_604),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_674),
.B(n_540),
.Y(n_868)
);

OAI321xp33_ASAP7_75t_L g869 ( 
.A1(n_744),
.A2(n_317),
.A3(n_316),
.B1(n_280),
.B2(n_274),
.C(n_334),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_713),
.B(n_488),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_801),
.A2(n_520),
.B(n_515),
.C(n_511),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_776),
.A2(n_527),
.B(n_523),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_794),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_756),
.A2(n_649),
.B(n_646),
.C(n_641),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_734),
.A2(n_284),
.B(n_280),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_680),
.A2(n_520),
.B(n_515),
.C(n_511),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_713),
.B(n_521),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_705),
.B(n_540),
.Y(n_878)
);

NOR2x1p5_ASAP7_75t_L g879 ( 
.A(n_686),
.B(n_249),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_776),
.A2(n_529),
.B(n_527),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_805),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_671),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_764),
.B(n_521),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_698),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_776),
.A2(n_529),
.B(n_527),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_707),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_722),
.A2(n_649),
.B(n_646),
.C(n_641),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_816),
.A2(n_535),
.B(n_529),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_665),
.A2(n_537),
.B(n_535),
.Y(n_889)
);

AOI21x1_ASAP7_75t_L g890 ( 
.A1(n_817),
.A2(n_537),
.B(n_535),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_666),
.A2(n_545),
.B(n_537),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_658),
.B(n_404),
.Y(n_892)
);

BUFx4f_ASAP7_75t_L g893 ( 
.A(n_749),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_699),
.B(n_297),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_709),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_656),
.A2(n_562),
.B(n_545),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_705),
.B(n_575),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_668),
.B(n_546),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_811),
.A2(n_562),
.B(n_545),
.Y(n_899)
);

CKINVDCx6p67_ASAP7_75t_R g900 ( 
.A(n_671),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_725),
.B(n_575),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_726),
.B(n_575),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_728),
.B(n_604),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_668),
.A2(n_564),
.B(n_562),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_742),
.A2(n_515),
.B(n_520),
.C(n_511),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_764),
.B(n_253),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_734),
.A2(n_565),
.B(n_564),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_604),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_740),
.A2(n_565),
.B(n_564),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_709),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_727),
.A2(n_604),
.B1(n_607),
.B2(n_615),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_740),
.A2(n_721),
.B(n_660),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_729),
.A2(n_649),
.B(n_639),
.C(n_565),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_805),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_789),
.A2(n_591),
.B(n_639),
.C(n_585),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_667),
.A2(n_582),
.B(n_576),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_710),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_796),
.A2(n_821),
.B(n_818),
.C(n_696),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_702),
.A2(n_582),
.B(n_576),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_796),
.A2(n_591),
.B(n_639),
.C(n_585),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_710),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_736),
.B(n_607),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_751),
.B(n_607),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_733),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_754),
.B(n_607),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_757),
.B(n_615),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_733),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_742),
.A2(n_500),
.B(n_501),
.C(n_502),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_704),
.A2(n_716),
.B(n_753),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_739),
.B(n_615),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_797),
.A2(n_576),
.B(n_582),
.Y(n_931)
);

NOR2xp67_ASAP7_75t_L g932 ( 
.A(n_780),
.B(n_670),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_739),
.B(n_615),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_741),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_689),
.B(n_195),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_699),
.B(n_301),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_708),
.B(n_195),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_723),
.A2(n_585),
.B(n_588),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_821),
.A2(n_697),
.B(n_681),
.C(n_664),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_762),
.B(n_637),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_769),
.B(n_637),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_805),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_724),
.A2(n_593),
.B(n_588),
.Y(n_943)
);

BUFx12f_ASAP7_75t_L g944 ( 
.A(n_774),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_814),
.A2(n_588),
.B(n_591),
.C(n_630),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_795),
.B(n_256),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_746),
.A2(n_601),
.B(n_592),
.Y(n_947)
);

AOI33xp33_ASAP7_75t_L g948 ( 
.A1(n_822),
.A2(n_325),
.A3(n_284),
.B1(n_316),
.B2(n_317),
.B3(n_419),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_748),
.A2(n_637),
.B1(n_592),
.B2(n_630),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_805),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_654),
.A2(n_592),
.B1(n_593),
.B2(n_630),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_654),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_741),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_781),
.B(n_637),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_793),
.B(n_798),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_664),
.B(n_593),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_787),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_667),
.A2(n_693),
.B(n_679),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_669),
.B(n_601),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_743),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_669),
.A2(n_601),
.B1(n_621),
.B2(n_620),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_676),
.A2(n_621),
.B(n_620),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_683),
.A2(n_621),
.B(n_620),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_672),
.B(n_267),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_672),
.A2(n_673),
.B(n_679),
.Y(n_965)
);

AO22x1_ASAP7_75t_L g966 ( 
.A1(n_749),
.A2(n_271),
.B1(n_278),
.B2(n_283),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_787),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_749),
.B(n_408),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_748),
.A2(n_502),
.B(n_500),
.C(n_508),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_766),
.B(n_408),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_673),
.A2(n_325),
.B1(n_195),
.B2(n_481),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_693),
.A2(n_642),
.B(n_573),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_791),
.B(n_792),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_703),
.A2(n_642),
.B(n_573),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_703),
.A2(n_642),
.B(n_573),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_791),
.B(n_546),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_755),
.A2(n_323),
.B1(n_302),
.B2(n_328),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_792),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_731),
.B(n_546),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_770),
.A2(n_501),
.B(n_500),
.C(n_502),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_731),
.B(n_546),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_770),
.B(n_410),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_770),
.B(n_546),
.Y(n_983)
);

AND3x1_ASAP7_75t_SL g984 ( 
.A(n_810),
.B(n_419),
.C(n_418),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_657),
.B(n_719),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_755),
.A2(n_330),
.B1(n_304),
.B2(n_321),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_747),
.A2(n_508),
.B(n_501),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_786),
.B(n_546),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_820),
.A2(n_573),
.B(n_642),
.Y(n_989)
);

OR2x2_ASAP7_75t_SL g990 ( 
.A(n_767),
.B(n_410),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_807),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_759),
.A2(n_508),
.B(n_418),
.C(n_463),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_745),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_730),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_788),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_809),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_799),
.B(n_573),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_809),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_800),
.B(n_758),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_711),
.A2(n_642),
.B(n_573),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_815),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_711),
.A2(n_642),
.B(n_440),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_706),
.Y(n_1003)
);

BUFx4f_ASAP7_75t_SL g1004 ( 
.A(n_759),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_760),
.A2(n_423),
.B(n_481),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_SL g1006 ( 
.A(n_671),
.B(n_305),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_802),
.B(n_309),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_718),
.A2(n_440),
.B(n_434),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_745),
.A2(n_320),
.B(n_313),
.C(n_306),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_772),
.B(n_785),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_772),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_804),
.B(n_452),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_812),
.B(n_452),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_826),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_834),
.B(n_718),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_SL g1016 ( 
.A1(n_985),
.A2(n_790),
.B1(n_682),
.B2(n_195),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_852),
.A2(n_720),
.B1(n_819),
.B2(n_763),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_SL g1018 ( 
.A1(n_939),
.A2(n_785),
.B(n_806),
.C(n_768),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_824),
.A2(n_856),
.B(n_843),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_838),
.A2(n_806),
.B(n_765),
.C(n_761),
.Y(n_1020)
);

OAI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_946),
.A2(n_287),
.B(n_293),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_838),
.A2(n_773),
.B(n_784),
.C(n_783),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_881),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_829),
.A2(n_833),
.B(n_918),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_912),
.A2(n_775),
.B(n_777),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_848),
.A2(n_815),
.B(n_779),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_881),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_SL g1028 ( 
.A(n_906),
.B(n_327),
.C(n_303),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_855),
.A2(n_445),
.B(n_434),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_845),
.B(n_849),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_991),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_883),
.A2(n_790),
.B1(n_578),
.B2(n_299),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_828),
.B(n_307),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_968),
.B(n_790),
.Y(n_1034)
);

O2A1O1Ixp5_ASAP7_75t_L g1035 ( 
.A1(n_825),
.A2(n_486),
.B(n_454),
.C(n_477),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_SL g1036 ( 
.A(n_883),
.B(n_311),
.C(n_315),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_893),
.A2(n_318),
.B1(n_324),
.B2(n_326),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_881),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_866),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_946),
.A2(n_332),
.B(n_333),
.C(n_454),
.Y(n_1040)
);

OAI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_1004),
.A2(n_578),
.B1(n_486),
.B2(n_454),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_836),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_893),
.B(n_452),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_828),
.B(n_454),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_877),
.B(n_452),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_995),
.B(n_463),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_906),
.A2(n_463),
.B(n_467),
.C(n_474),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_841),
.A2(n_434),
.B(n_445),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_935),
.A2(n_467),
.B(n_477),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_831),
.A2(n_578),
.B1(n_440),
.B2(n_434),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_907),
.A2(n_474),
.B(n_486),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_836),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_881),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_832),
.A2(n_999),
.B(n_863),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_835),
.A2(n_467),
.B(n_477),
.C(n_474),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_832),
.A2(n_434),
.B(n_445),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_850),
.B(n_4),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_952),
.Y(n_1058)
);

AOI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_869),
.A2(n_467),
.B1(n_477),
.B2(n_474),
.C(n_486),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_955),
.B(n_463),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_854),
.B(n_482),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_991),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_960),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_835),
.A2(n_440),
.B(n_452),
.C(n_482),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_1004),
.B(n_482),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_884),
.Y(n_1066)
);

AO32x1_ASAP7_75t_L g1067 ( 
.A1(n_951),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_950),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_888),
.A2(n_445),
.B(n_434),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_862),
.A2(n_445),
.B(n_440),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_884),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_842),
.B(n_67),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_830),
.B(n_578),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_968),
.Y(n_1074)
);

OR2x6_ASAP7_75t_SL g1075 ( 
.A(n_882),
.B(n_5),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_950),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_858),
.A2(n_452),
.B(n_482),
.C(n_445),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_864),
.Y(n_1078)
);

AOI22x1_ASAP7_75t_L g1079 ( 
.A1(n_929),
.A2(n_482),
.B1(n_452),
.B2(n_445),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_898),
.A2(n_872),
.B(n_865),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_950),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_892),
.B(n_482),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_988),
.A2(n_445),
.B(n_482),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_847),
.A2(n_578),
.B1(n_482),
.B2(n_452),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_994),
.B(n_6),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_997),
.A2(n_860),
.B(n_899),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_973),
.A2(n_423),
.B(n_481),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_982),
.B(n_164),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_SL g1089 ( 
.A1(n_983),
.A2(n_10),
.B(n_11),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_964),
.B(n_982),
.Y(n_1090)
);

NOR2x1p5_ASAP7_75t_L g1091 ( 
.A(n_900),
.B(n_163),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1003),
.A2(n_1010),
.B1(n_964),
.B2(n_1011),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1010),
.A2(n_481),
.B1(n_423),
.B2(n_17),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_965),
.A2(n_423),
.B(n_481),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_870),
.B(n_481),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_932),
.B(n_12),
.C(n_14),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_990),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_895),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_L g1099 ( 
.A1(n_887),
.A2(n_114),
.B(n_70),
.C(n_154),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_879),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_853),
.B(n_149),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_921),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_886),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_878),
.B(n_481),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_880),
.A2(n_423),
.B(n_481),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_897),
.B(n_481),
.Y(n_1106)
);

BUFx4f_ASAP7_75t_L g1107 ( 
.A(n_944),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_970),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_851),
.B(n_140),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_924),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_927),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1006),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_861),
.A2(n_14),
.B(n_17),
.C(n_21),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_898),
.A2(n_885),
.B(n_956),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_953),
.B(n_481),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_937),
.A2(n_948),
.B(n_977),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_957),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_853),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_993),
.B(n_135),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_978),
.B(n_481),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_909),
.A2(n_423),
.B(n_131),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1011),
.B(n_127),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_993),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_934),
.B(n_423),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_967),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_984),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_993),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_910),
.B(n_423),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_993),
.B(n_950),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_SL g1130 ( 
.A(n_1009),
.B(n_22),
.C(n_24),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_952),
.B(n_119),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_917),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_952),
.B(n_117),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_966),
.B(n_952),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_859),
.A2(n_986),
.B1(n_1007),
.B2(n_911),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_846),
.B(n_423),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_913),
.A2(n_107),
.B(n_99),
.C(n_98),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_839),
.A2(n_85),
.B(n_83),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_827),
.B(n_88),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_827),
.B(n_75),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_959),
.A2(n_68),
.B(n_27),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_894),
.B(n_25),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_840),
.A2(n_30),
.B(n_32),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_983),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_846),
.B(n_33),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_867),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_SL g1147 ( 
.A(n_936),
.B(n_41),
.C(n_46),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_873),
.B(n_47),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_984),
.A2(n_59),
.B1(n_49),
.B2(n_52),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_873),
.B(n_48),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_981),
.A2(n_52),
.B(n_54),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_914),
.B(n_54),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_868),
.A2(n_55),
.B(n_58),
.Y(n_1153)
);

NOR2x1_ASAP7_75t_L g1154 ( 
.A(n_857),
.B(n_55),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_914),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_976),
.A2(n_58),
.B(n_844),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_920),
.A2(n_1013),
.B(n_1012),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_857),
.B(n_942),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_942),
.B(n_996),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_998),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_989),
.A2(n_874),
.B(n_896),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_SL g1162 ( 
.A1(n_992),
.A2(n_876),
.B(n_905),
.C(n_1005),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_938),
.A2(n_947),
.B(n_943),
.Y(n_1163)
);

AND2x2_ASAP7_75t_SL g1164 ( 
.A(n_971),
.B(n_902),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_979),
.B(n_901),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_933),
.B(n_930),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_L g1167 ( 
.A(n_971),
.B(n_915),
.C(n_992),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_889),
.A2(n_891),
.B(n_931),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1001),
.B(n_940),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_933),
.B(n_875),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1142),
.A2(n_876),
.B(n_905),
.C(n_980),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1014),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1097),
.A2(n_926),
.B1(n_954),
.B2(n_941),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1026),
.A2(n_837),
.B(n_890),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1029),
.A2(n_987),
.B(n_916),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_SL g1176 ( 
.A(n_1166),
.B(n_958),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1030),
.B(n_1090),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1023),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1020),
.A2(n_949),
.B(n_919),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_904),
.B(n_962),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1063),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1092),
.B(n_903),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1019),
.A2(n_963),
.B(n_961),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_L g1184 ( 
.A(n_1108),
.B(n_908),
.Y(n_1184)
);

OAI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1085),
.A2(n_922),
.B1(n_923),
.B2(n_925),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1116),
.A2(n_871),
.B(n_928),
.C(n_969),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1039),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1015),
.B(n_871),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1019),
.A2(n_1000),
.B(n_974),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1146),
.A2(n_972),
.B1(n_975),
.B2(n_1002),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1024),
.A2(n_928),
.B(n_969),
.Y(n_1191)
);

OAI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1149),
.A2(n_945),
.B1(n_1008),
.B2(n_1134),
.Y(n_1192)
);

INVx6_ASAP7_75t_SL g1193 ( 
.A(n_1034),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1028),
.A2(n_945),
.B1(n_1126),
.B2(n_1021),
.Y(n_1194)
);

AOI221x1_ASAP7_75t_L g1195 ( 
.A1(n_1156),
.A2(n_1024),
.B1(n_1096),
.B2(n_1161),
.C(n_1163),
.Y(n_1195)
);

AOI221x1_ASAP7_75t_L g1196 ( 
.A1(n_1161),
.A2(n_1163),
.B1(n_1168),
.B2(n_1086),
.C(n_1157),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1086),
.A2(n_1026),
.B(n_1018),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1071),
.B(n_1066),
.Y(n_1198)
);

INVxp67_ASAP7_75t_SL g1199 ( 
.A(n_1052),
.Y(n_1199)
);

BUFx16f_ASAP7_75t_R g1200 ( 
.A(n_1034),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1033),
.B(n_1160),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1042),
.B(n_1074),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1118),
.B(n_1101),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1155),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1023),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1154),
.A2(n_1122),
.B1(n_1057),
.B2(n_1150),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1029),
.A2(n_1080),
.B(n_1070),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1070),
.A2(n_1114),
.B(n_1051),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1025),
.A2(n_1135),
.B(n_1157),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1023),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_SL g1212 ( 
.A1(n_1162),
.A2(n_1133),
.B(n_1131),
.C(n_1119),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1025),
.A2(n_1017),
.B(n_1022),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1165),
.A2(n_1164),
.B(n_1064),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1037),
.B(n_1112),
.Y(n_1215)
);

BUFx5_ASAP7_75t_L g1216 ( 
.A(n_1140),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1168),
.A2(n_1077),
.B(n_1069),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1027),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1101),
.B(n_1088),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1069),
.A2(n_1079),
.B(n_1099),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1100),
.B(n_1088),
.Y(n_1221)
);

INVx6_ASAP7_75t_L g1222 ( 
.A(n_1122),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_SL g1223 ( 
.A(n_1166),
.B(n_1061),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1123),
.B(n_1127),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1055),
.A2(n_1084),
.A3(n_1050),
.B(n_1040),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1095),
.A2(n_1167),
.B(n_1106),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1083),
.A2(n_1048),
.B(n_1121),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1083),
.A2(n_1056),
.B(n_1035),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1107),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1098),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1027),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1138),
.A2(n_1143),
.A3(n_1094),
.B(n_1145),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1060),
.A2(n_1169),
.B(n_1049),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1102),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_1058),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1138),
.A2(n_1094),
.A3(n_1148),
.B(n_1141),
.Y(n_1236)
);

NAND3x1_ASAP7_75t_L g1237 ( 
.A(n_1075),
.B(n_1153),
.C(n_1151),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1152),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1104),
.A2(n_1144),
.B(n_1170),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1016),
.B(n_1147),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1117),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1113),
.A2(n_1036),
.B(n_1089),
.C(n_1137),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1072),
.B(n_1103),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1027),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1129),
.A2(n_1041),
.B(n_1065),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1159),
.A2(n_1139),
.B(n_1166),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1107),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1047),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1125),
.B(n_1132),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1032),
.A2(n_1109),
.B1(n_1073),
.B2(n_1078),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_SL g1252 ( 
.A1(n_1115),
.A2(n_1120),
.B(n_1136),
.C(n_1082),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1124),
.A2(n_1128),
.B(n_1087),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1105),
.A2(n_1031),
.B(n_1062),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1093),
.A2(n_1091),
.B1(n_1081),
.B2(n_1076),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1130),
.A2(n_1105),
.B(n_1081),
.C(n_1059),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1038),
.Y(n_1257)
);

AO22x2_ASAP7_75t_L g1258 ( 
.A1(n_1067),
.A2(n_1038),
.B1(n_1053),
.B2(n_1068),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1038),
.B(n_1053),
.Y(n_1259)
);

CKINVDCx8_ASAP7_75t_R g1260 ( 
.A(n_1053),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1068),
.B(n_1076),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1068),
.A2(n_1076),
.B1(n_1059),
.B2(n_1067),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1067),
.A2(n_1024),
.A3(n_1019),
.B(n_1064),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1030),
.B(n_691),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1030),
.B(n_691),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1054),
.A2(n_852),
.B(n_824),
.Y(n_1266)
);

AOI221x1_ASAP7_75t_L g1267 ( 
.A1(n_1156),
.A2(n_852),
.B1(n_1019),
.B2(n_1024),
.C(n_1146),
.Y(n_1267)
);

NAND3x1_ASAP7_75t_L g1268 ( 
.A(n_1085),
.B(n_661),
.C(n_536),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1054),
.A2(n_852),
.B(n_824),
.Y(n_1269)
);

BUFx4_ASAP7_75t_SL g1270 ( 
.A(n_1126),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1034),
.B(n_1101),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1030),
.B(n_691),
.Y(n_1272)
);

AOI221x1_ASAP7_75t_L g1273 ( 
.A1(n_1156),
.A2(n_852),
.B1(n_1019),
.B2(n_1024),
.C(n_1146),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1030),
.B(n_691),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1097),
.B(n_877),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1014),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1054),
.A2(n_852),
.B(n_824),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1063),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1063),
.B(n_557),
.Y(n_1280)
);

AO32x2_ASAP7_75t_L g1281 ( 
.A1(n_1146),
.A2(n_1017),
.A3(n_730),
.B1(n_961),
.B2(n_951),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1090),
.B(n_657),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1033),
.A2(n_852),
.B(n_691),
.C(n_661),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1030),
.B(n_691),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1162),
.A2(n_852),
.B(n_918),
.C(n_939),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1042),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1024),
.A2(n_1019),
.A3(n_1064),
.B(n_1077),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1014),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1023),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1033),
.A2(n_852),
.B(n_691),
.C(n_661),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1063),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1090),
.B(n_362),
.Y(n_1294)
);

AO22x2_ASAP7_75t_L g1295 ( 
.A1(n_1146),
.A2(n_1147),
.B1(n_727),
.B2(n_1096),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1030),
.B(n_691),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1030),
.B(n_691),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1033),
.A2(n_852),
.B(n_691),
.C(n_661),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1142),
.B(n_852),
.C(n_691),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1097),
.B(n_877),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1030),
.B(n_691),
.Y(n_1302)
);

AO32x2_ASAP7_75t_L g1303 ( 
.A1(n_1146),
.A2(n_1017),
.A3(n_730),
.B1(n_961),
.B2(n_951),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1097),
.B(n_877),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1028),
.A2(n_661),
.B1(n_657),
.B2(n_365),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1063),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1063),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1024),
.A2(n_1019),
.A3(n_1064),
.B(n_1077),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1033),
.A2(n_852),
.B(n_691),
.C(n_661),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1014),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1030),
.B(n_691),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1033),
.A2(n_852),
.B(n_691),
.C(n_661),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1014),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1107),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1097),
.A2(n_727),
.B1(n_691),
.B2(n_985),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1063),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1029),
.A2(n_987),
.B(n_1080),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1030),
.B(n_691),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1024),
.A2(n_1019),
.B(n_1161),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1030),
.B(n_691),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1033),
.A2(n_852),
.B(n_691),
.C(n_661),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1097),
.B(n_877),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1014),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1054),
.A2(n_852),
.B(n_824),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1030),
.B(n_691),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1014),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1023),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1028),
.A2(n_661),
.B1(n_657),
.B2(n_365),
.Y(n_1330)
);

NAND2xp33_ASAP7_75t_L g1331 ( 
.A(n_1112),
.B(n_852),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1090),
.B(n_362),
.Y(n_1332)
);

NOR2xp67_ASAP7_75t_SL g1333 ( 
.A(n_1063),
.B(n_830),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1118),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1240),
.A2(n_1300),
.B1(n_1295),
.B2(n_1331),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1268),
.A2(n_1297),
.B1(n_1296),
.B2(n_1302),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1229),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1295),
.A2(n_1282),
.B1(n_1317),
.B2(n_1305),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1242),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1292),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1248),
.Y(n_1341)
);

BUFx4f_ASAP7_75t_L g1342 ( 
.A(n_1271),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1330),
.A2(n_1294),
.B1(n_1332),
.B2(n_1207),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1215),
.A2(n_1265),
.B1(n_1312),
.B2(n_1285),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1315),
.Y(n_1345)
);

INVx6_ASAP7_75t_L g1346 ( 
.A(n_1221),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1306),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1221),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1264),
.A2(n_1275),
.B1(n_1272),
.B2(n_1327),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1320),
.A2(n_1322),
.B1(n_1201),
.B2(n_1177),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1334),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1280),
.B(n_1307),
.Y(n_1352)
);

BUFx4_ASAP7_75t_SL g1353 ( 
.A(n_1271),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1266),
.A2(n_1278),
.B(n_1326),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1277),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1277),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1276),
.B(n_1301),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1260),
.Y(n_1358)
);

BUFx8_ASAP7_75t_L g1359 ( 
.A(n_1244),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1304),
.B(n_1324),
.Y(n_1360)
);

BUFx8_ASAP7_75t_L g1361 ( 
.A(n_1203),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1289),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1289),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1181),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1222),
.A2(n_1241),
.B1(n_1328),
.B2(n_1325),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1222),
.A2(n_1311),
.B1(n_1325),
.B2(n_1328),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1311),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1194),
.A2(n_1182),
.B1(n_1219),
.B2(n_1214),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1238),
.A2(n_1279),
.B1(n_1213),
.B2(n_1173),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1204),
.B(n_1284),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1314),
.A2(n_1258),
.B1(n_1237),
.B2(n_1313),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1314),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1291),
.B(n_1299),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1187),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1200),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1270),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1287),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1245),
.B(n_1329),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1203),
.A2(n_1216),
.B1(n_1318),
.B2(n_1184),
.Y(n_1379)
);

BUFx5_ASAP7_75t_L g1380 ( 
.A(n_1234),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1310),
.A2(n_1323),
.B(n_1273),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1216),
.A2(n_1258),
.B1(n_1223),
.B2(n_1269),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1250),
.Y(n_1383)
);

INVx6_ASAP7_75t_L g1384 ( 
.A(n_1245),
.Y(n_1384)
);

INVx8_ASAP7_75t_L g1385 ( 
.A(n_1245),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1198),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_1224),
.Y(n_1387)
);

BUFx8_ASAP7_75t_SL g1388 ( 
.A(n_1224),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1329),
.B(n_1205),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1216),
.A2(n_1210),
.B1(n_1199),
.B2(n_1179),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1216),
.A2(n_1202),
.B1(n_1226),
.B2(n_1255),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1216),
.A2(n_1176),
.B1(n_1321),
.B2(n_1249),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1261),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1262),
.A2(n_1188),
.B1(n_1186),
.B2(n_1256),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1185),
.A2(n_1251),
.B1(n_1333),
.B2(n_1286),
.Y(n_1395)
);

BUFx8_ASAP7_75t_L g1396 ( 
.A(n_1178),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1259),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1178),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1218),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1192),
.A2(n_1247),
.B1(n_1239),
.B2(n_1246),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1218),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1329),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1257),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1243),
.A2(n_1171),
.B1(n_1235),
.B2(n_1193),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1206),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1206),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1211),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1321),
.A2(n_1197),
.B1(n_1190),
.B2(n_1220),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1267),
.B(n_1195),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1211),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1253),
.A2(n_1254),
.B1(n_1193),
.B2(n_1190),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1257),
.B(n_1290),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1290),
.Y(n_1413)
);

INVx5_ASAP7_75t_L g1414 ( 
.A(n_1211),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1231),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1217),
.A2(n_1233),
.B1(n_1191),
.B2(n_1231),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1220),
.A2(n_1303),
.B1(n_1281),
.B2(n_1212),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1281),
.B(n_1303),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1288),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1183),
.A2(n_1180),
.B1(n_1189),
.B2(n_1174),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1281),
.A2(n_1303),
.B1(n_1263),
.B2(n_1196),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1263),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1217),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1263),
.A2(n_1308),
.B1(n_1288),
.B2(n_1225),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1208),
.A2(n_1227),
.B1(n_1319),
.B2(n_1274),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1288),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1252),
.Y(n_1427)
);

BUFx4f_ASAP7_75t_SL g1428 ( 
.A(n_1236),
.Y(n_1428)
);

BUFx4f_ASAP7_75t_SL g1429 ( 
.A(n_1236),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_SL g1430 ( 
.A(n_1236),
.Y(n_1430)
);

NOR3xp33_ASAP7_75t_L g1431 ( 
.A(n_1316),
.B(n_1283),
.C(n_1298),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1308),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1228),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1232),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1308),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1175),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1225),
.B(n_1293),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1225),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1309),
.Y(n_1439)
);

BUFx2_ASAP7_75t_SL g1440 ( 
.A(n_1209),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1306),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1172),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1260),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1305),
.A2(n_657),
.B1(n_1330),
.B2(n_551),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1248),
.Y(n_1445)
);

AO22x1_ASAP7_75t_L g1446 ( 
.A1(n_1240),
.A2(n_661),
.B1(n_1085),
.B2(n_778),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1230),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1200),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1240),
.A2(n_657),
.B1(n_661),
.B2(n_1004),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1268),
.A2(n_852),
.B1(n_1300),
.B2(n_1265),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1264),
.B(n_1265),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1229),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1268),
.A2(n_852),
.B1(n_1300),
.B2(n_1265),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1268),
.A2(n_852),
.B1(n_1300),
.B2(n_1265),
.Y(n_1454)
);

BUFx8_ASAP7_75t_L g1455 ( 
.A(n_1229),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1248),
.Y(n_1456)
);

CKINVDCx6p67_ASAP7_75t_R g1457 ( 
.A(n_1229),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1230),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1240),
.A2(n_657),
.B1(n_661),
.B2(n_1004),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1276),
.B(n_1301),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1172),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1268),
.A2(n_852),
.B1(n_1300),
.B2(n_1265),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1268),
.A2(n_661),
.B1(n_852),
.B2(n_1317),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1292),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1305),
.A2(n_657),
.B1(n_1330),
.B2(n_551),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1240),
.A2(n_1300),
.B1(n_661),
.B2(n_727),
.Y(n_1466)
);

BUFx10_ASAP7_75t_L g1467 ( 
.A(n_1248),
.Y(n_1467)
);

CKINVDCx6p67_ASAP7_75t_R g1468 ( 
.A(n_1229),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1268),
.A2(n_852),
.B1(n_1300),
.B2(n_1265),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1260),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1240),
.A2(n_1300),
.B1(n_661),
.B2(n_727),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1268),
.A2(n_1240),
.B1(n_1300),
.B2(n_661),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1268),
.A2(n_1240),
.B1(n_1300),
.B2(n_661),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1306),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1287),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1347),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1463),
.A2(n_1473),
.B(n_1472),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1422),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1342),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1444),
.A2(n_1465),
.B1(n_1335),
.B2(n_1449),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1354),
.A2(n_1420),
.B(n_1425),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1437),
.A2(n_1439),
.B(n_1416),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1426),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1373),
.A2(n_1409),
.B(n_1450),
.Y(n_1484)
);

INVxp33_ASAP7_75t_L g1485 ( 
.A(n_1360),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1432),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1435),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1438),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1419),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1418),
.B(n_1372),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1380),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1436),
.A2(n_1424),
.B(n_1404),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1472),
.A2(n_1473),
.B(n_1471),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1355),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1466),
.A2(n_1450),
.B(n_1454),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1423),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1356),
.B(n_1362),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1350),
.B(n_1344),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1363),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1367),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1459),
.A2(n_1338),
.B1(n_1469),
.B2(n_1454),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1352),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1442),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1342),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1424),
.A2(n_1400),
.B(n_1411),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1384),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1396),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1446),
.B(n_1336),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1370),
.B(n_1371),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1461),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1341),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1453),
.A2(n_1469),
.B1(n_1462),
.B2(n_1343),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1434),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1430),
.Y(n_1514)
);

AOI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1453),
.A2(n_1462),
.B(n_1371),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1417),
.B(n_1397),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1430),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1433),
.B(n_1374),
.Y(n_1518)
);

AOI21xp33_ASAP7_75t_L g1519 ( 
.A1(n_1381),
.A2(n_1336),
.B(n_1395),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1417),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1384),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1428),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1421),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1421),
.Y(n_1524)
);

NAND2x1p5_ASAP7_75t_L g1525 ( 
.A(n_1395),
.B(n_1414),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1394),
.A2(n_1381),
.B(n_1366),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1349),
.A2(n_1369),
.B1(n_1368),
.B2(n_1451),
.C(n_1391),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1385),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1366),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1339),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1394),
.A2(n_1365),
.B(n_1440),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1429),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1376),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1447),
.Y(n_1534)
);

AOI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1365),
.A2(n_1399),
.B(n_1403),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1408),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1464),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1393),
.B(n_1357),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1441),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1460),
.B(n_1458),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1383),
.B(n_1474),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1390),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1345),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1427),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1382),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1359),
.A2(n_1427),
.B1(n_1348),
.B2(n_1340),
.Y(n_1546)
);

AO21x1_ASAP7_75t_L g1547 ( 
.A1(n_1431),
.A2(n_1401),
.B(n_1413),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1379),
.A2(n_1392),
.B(n_1364),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1427),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1412),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1414),
.B(n_1415),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1475),
.B(n_1386),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1389),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1378),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1414),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1475),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1377),
.B(n_1386),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1385),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1415),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1415),
.A2(n_1402),
.B(n_1410),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1398),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1398),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1406),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1346),
.A2(n_1358),
.B1(n_1470),
.B2(n_1443),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1353),
.A2(n_1396),
.B(n_1361),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1443),
.B(n_1361),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1405),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1443),
.A2(n_1387),
.B(n_1348),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1375),
.B(n_1448),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1407),
.A2(n_1359),
.B(n_1388),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1351),
.B(n_1468),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1337),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1337),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1455),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1452),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1452),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1457),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1455),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1467),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1496),
.B(n_1467),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1502),
.B(n_1445),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_SL g1582 ( 
.A1(n_1495),
.A2(n_1456),
.B(n_1493),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_SL g1583 ( 
.A1(n_1519),
.A2(n_1498),
.B(n_1477),
.C(n_1508),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1512),
.A2(n_1501),
.B(n_1480),
.C(n_1527),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1585)
);

BUFx10_ASAP7_75t_L g1586 ( 
.A(n_1557),
.Y(n_1586)
);

AO32x2_ASAP7_75t_L g1587 ( 
.A1(n_1520),
.A2(n_1484),
.A3(n_1523),
.B1(n_1524),
.B2(n_1516),
.Y(n_1587)
);

AND2x2_ASAP7_75t_SL g1588 ( 
.A(n_1496),
.B(n_1509),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1542),
.A2(n_1509),
.B1(n_1523),
.B2(n_1524),
.C(n_1520),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_R g1590 ( 
.A(n_1511),
.B(n_1543),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1526),
.A2(n_1542),
.B1(n_1545),
.B2(n_1525),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1545),
.B(n_1484),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_R g1593 ( 
.A(n_1574),
.B(n_1507),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1526),
.A2(n_1505),
.B(n_1531),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1550),
.B(n_1476),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1550),
.B(n_1556),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1546),
.A2(n_1485),
.B1(n_1525),
.B2(n_1479),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1505),
.A2(n_1531),
.B(n_1492),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1497),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1548),
.A2(n_1504),
.B(n_1479),
.C(n_1565),
.Y(n_1600)
);

INVx5_ASAP7_75t_L g1601 ( 
.A(n_1522),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1513),
.B(n_1532),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1538),
.B(n_1490),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1486),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1540),
.B(n_1516),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_SL g1606 ( 
.A(n_1564),
.B(n_1533),
.C(n_1568),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1540),
.B(n_1497),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_SL g1608 ( 
.A(n_1569),
.B(n_1558),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1479),
.A2(n_1504),
.B(n_1565),
.C(n_1560),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1537),
.A2(n_1552),
.B(n_1553),
.C(n_1579),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_SL g1612 ( 
.A(n_1535),
.B(n_1514),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1553),
.A2(n_1579),
.B(n_1529),
.C(n_1536),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1561),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1504),
.A2(n_1578),
.B1(n_1574),
.B2(n_1507),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1562),
.Y(n_1617)
);

NAND4xp25_ASAP7_75t_L g1618 ( 
.A(n_1577),
.B(n_1536),
.C(n_1529),
.D(n_1514),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1518),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1547),
.A2(n_1482),
.B(n_1481),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1577),
.A2(n_1572),
.B(n_1532),
.C(n_1573),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1522),
.B(n_1513),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1566),
.A2(n_1576),
.B1(n_1573),
.B2(n_1507),
.Y(n_1623)
);

O2A1O1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1576),
.A2(n_1517),
.B(n_1578),
.C(n_1566),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1517),
.B(n_1513),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1566),
.A2(n_1569),
.B1(n_1575),
.B2(n_1574),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1571),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1483),
.A2(n_1535),
.B(n_1478),
.Y(n_1629)
);

AO32x2_ASAP7_75t_L g1630 ( 
.A1(n_1506),
.A2(n_1521),
.A3(n_1528),
.B1(n_1558),
.B2(n_1478),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1549),
.B(n_1554),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1500),
.B(n_1510),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1578),
.A2(n_1506),
.B(n_1521),
.C(n_1544),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1486),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1584),
.B(n_1583),
.C(n_1600),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1634),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1598),
.B(n_1594),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1629),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1510),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1592),
.B(n_1503),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1604),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1582),
.A2(n_1570),
.B1(n_1578),
.B2(n_1571),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1598),
.B(n_1486),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1583),
.B(n_1563),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1594),
.B(n_1487),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1585),
.B(n_1503),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1599),
.B(n_1620),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1620),
.B(n_1488),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1612),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1630),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1587),
.B(n_1489),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1591),
.A2(n_1569),
.B(n_1571),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1587),
.B(n_1489),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1587),
.B(n_1489),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1630),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1591),
.A2(n_1551),
.B(n_1544),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1615),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1630),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1587),
.B(n_1491),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1628),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1588),
.A2(n_1570),
.B1(n_1534),
.B2(n_1530),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1650),
.B(n_1609),
.Y(n_1664)
);

NAND2x1p5_ASAP7_75t_L g1665 ( 
.A(n_1648),
.B(n_1601),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1635),
.A2(n_1589),
.B1(n_1618),
.B2(n_1597),
.C(n_1611),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1636),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1635),
.A2(n_1626),
.B(n_1610),
.C(n_1624),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1652),
.A2(n_1589),
.B1(n_1611),
.B2(n_1613),
.C(n_1606),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1650),
.B(n_1609),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1650),
.B(n_1609),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1639),
.B(n_1640),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1655),
.B(n_1614),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1652),
.A2(n_1606),
.B(n_1588),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1649),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1643),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1655),
.B(n_1614),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1652),
.A2(n_1627),
.B1(n_1616),
.B2(n_1605),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1636),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1641),
.Y(n_1680)
);

AND2x4_ASAP7_75t_SL g1681 ( 
.A(n_1663),
.B(n_1622),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.B(n_1614),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1658),
.B(n_1630),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1662),
.B(n_1595),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1637),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1601),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1646),
.B(n_1586),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1601),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1643),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1636),
.Y(n_1692)
);

OAI33xp33_ASAP7_75t_L g1693 ( 
.A1(n_1639),
.A2(n_1596),
.A3(n_1623),
.B1(n_1621),
.B2(n_1613),
.B3(n_1624),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1658),
.B(n_1607),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1640),
.B(n_1603),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1642),
.A2(n_1580),
.B1(n_1602),
.B2(n_1625),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1656),
.A2(n_1608),
.B(n_1625),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1659),
.B(n_1617),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1687),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1672),
.B(n_1686),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1687),
.B(n_1651),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1688),
.B(n_1645),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1687),
.B(n_1651),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1672),
.B(n_1660),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1687),
.B(n_1651),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1687),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1687),
.B(n_1653),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1667),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1688),
.B(n_1645),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1680),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1688),
.B(n_1645),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1676),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1684),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1684),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1679),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1683),
.B(n_1684),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1683),
.B(n_1653),
.Y(n_1718)
);

AND2x4_ASAP7_75t_SL g1719 ( 
.A(n_1688),
.B(n_1622),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1679),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1691),
.B(n_1638),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1692),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1664),
.B(n_1670),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1698),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1698),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1688),
.B(n_1690),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1707),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1723),
.B(n_1670),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1707),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1700),
.B(n_1693),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1728),
.B(n_1674),
.Y(n_1734)
);

NAND3xp33_ASAP7_75t_L g1735 ( 
.A(n_1704),
.B(n_1666),
.C(n_1668),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1704),
.B(n_1689),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1707),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1723),
.B(n_1671),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1711),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1709),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1709),
.Y(n_1741)
);

NAND2x1_ASAP7_75t_L g1742 ( 
.A(n_1728),
.B(n_1675),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1709),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1711),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1716),
.Y(n_1745)
);

NAND2x1_ASAP7_75t_SL g1746 ( 
.A(n_1728),
.B(n_1671),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1723),
.B(n_1728),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1717),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1723),
.Y(n_1749)
);

AOI21x1_ASAP7_75t_SL g1750 ( 
.A1(n_1728),
.A2(n_1682),
.B(n_1677),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1728),
.B(n_1690),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1725),
.B(n_1695),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1716),
.Y(n_1753)
);

NOR3xp33_ASAP7_75t_L g1754 ( 
.A(n_1699),
.B(n_1693),
.C(n_1666),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1694),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1725),
.B(n_1695),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1728),
.Y(n_1757)
);

OAI32xp33_ASAP7_75t_L g1758 ( 
.A1(n_1718),
.A2(n_1697),
.A3(n_1674),
.B1(n_1678),
.B2(n_1682),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1716),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1725),
.B(n_1644),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1719),
.B(n_1668),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1725),
.B(n_1685),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1720),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1719),
.B(n_1694),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1719),
.A2(n_1697),
.B1(n_1669),
.B2(n_1678),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1699),
.A2(n_1669),
.B1(n_1656),
.B2(n_1601),
.Y(n_1767)
);

INVxp33_ASAP7_75t_L g1768 ( 
.A(n_1699),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1717),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1720),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1726),
.B(n_1685),
.Y(n_1771)
);

AO221x1_ASAP7_75t_L g1772 ( 
.A1(n_1767),
.A2(n_1675),
.B1(n_1706),
.B2(n_1699),
.C(n_1722),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1746),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1739),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1749),
.B(n_1726),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1762),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1754),
.B(n_1621),
.C(n_1642),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1747),
.B(n_1724),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1770),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1730),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1753),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1733),
.B(n_1671),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1747),
.B(n_1724),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1729),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1732),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_1762),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1733),
.B(n_1673),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1737),
.Y(n_1789)
);

NAND4xp25_ASAP7_75t_L g1790 ( 
.A(n_1735),
.B(n_1696),
.C(n_1663),
.D(n_1656),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1730),
.B(n_1724),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1731),
.B(n_1726),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1761),
.B(n_1726),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1742),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1738),
.B(n_1724),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1740),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1736),
.B(n_1673),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1766),
.B(n_1673),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_L g1799 ( 
.A(n_1734),
.B(n_1570),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1744),
.B(n_1677),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1738),
.B(n_1677),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1734),
.B(n_1727),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1758),
.B(n_1586),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1741),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1743),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1734),
.B(n_1727),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1755),
.B(n_1682),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1777),
.B(n_1767),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1776),
.B(n_1765),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1787),
.A2(n_1764),
.B1(n_1768),
.B2(n_1751),
.C(n_1769),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1803),
.A2(n_1734),
.B1(n_1751),
.B2(n_1681),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1783),
.B(n_1752),
.Y(n_1812)
);

OAI21xp33_ASAP7_75t_L g1813 ( 
.A1(n_1788),
.A2(n_1756),
.B(n_1763),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1773),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1778),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1790),
.A2(n_1681),
.B(n_1649),
.C(n_1633),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1794),
.A2(n_1593),
.B(n_1751),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1798),
.A2(n_1757),
.B1(n_1681),
.B2(n_1665),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1781),
.B(n_1757),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_1771),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1773),
.A2(n_1757),
.B1(n_1690),
.B2(n_1712),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1778),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1799),
.B(n_1745),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1794),
.B(n_1590),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1782),
.B(n_1769),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

NOR2x1_ASAP7_75t_L g1827 ( 
.A(n_1782),
.B(n_1780),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1772),
.A2(n_1800),
.B(n_1797),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1772),
.A2(n_1781),
.B1(n_1806),
.B2(n_1802),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1802),
.B(n_1712),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1792),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1792),
.B(n_1748),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1779),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1814),
.B(n_1791),
.Y(n_1834)
);

NAND2x1_ASAP7_75t_L g1835 ( 
.A(n_1817),
.B(n_1823),
.Y(n_1835)
);

OAI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1808),
.A2(n_1827),
.B1(n_1828),
.B2(n_1820),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1809),
.B(n_1791),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1833),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1808),
.A2(n_1806),
.B(n_1804),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1824),
.A2(n_1829),
.B1(n_1816),
.B2(n_1811),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1824),
.B(n_1795),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1829),
.A2(n_1816),
.B1(n_1810),
.B2(n_1812),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1833),
.B(n_1795),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1831),
.A2(n_1768),
.B1(n_1807),
.B2(n_1775),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_SL g1845 ( 
.A1(n_1815),
.A2(n_1805),
.B(n_1785),
.C(n_1796),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1819),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1822),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1821),
.A2(n_1801),
.B1(n_1779),
.B2(n_1784),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1826),
.B(n_1784),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1825),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1832),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1813),
.Y(n_1852)
);

O2A1O1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1818),
.A2(n_1805),
.B(n_1796),
.C(n_1789),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1836),
.B(n_1793),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1834),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1838),
.Y(n_1856)
);

AOI221x1_ASAP7_75t_SL g1857 ( 
.A1(n_1836),
.A2(n_1789),
.B1(n_1786),
.B2(n_1785),
.C(n_1748),
.Y(n_1857)
);

XNOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1839),
.B(n_1581),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1849),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1842),
.B(n_1590),
.Y(n_1860)
);

OA211x2_ASAP7_75t_L g1861 ( 
.A1(n_1835),
.A2(n_1750),
.B(n_1631),
.C(n_1661),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1845),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1843),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1846),
.B(n_1786),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1841),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1863),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1860),
.B(n_1852),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1865),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1865),
.Y(n_1869)
);

AOI21xp33_ASAP7_75t_L g1870 ( 
.A1(n_1854),
.A2(n_1844),
.B(n_1853),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1854),
.B(n_1850),
.Y(n_1871)
);

OAI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1857),
.A2(n_1840),
.B1(n_1851),
.B2(n_1837),
.C(n_1848),
.Y(n_1872)
);

AOI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1860),
.A2(n_1844),
.B1(n_1847),
.B2(n_1830),
.C(n_1775),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1858),
.A2(n_1862),
.B1(n_1861),
.B2(n_1855),
.Y(n_1874)
);

NOR3xp33_ASAP7_75t_L g1875 ( 
.A(n_1859),
.B(n_1847),
.C(n_1793),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1864),
.B(n_1759),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1867),
.B(n_1856),
.Y(n_1877)
);

O2A1O1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1870),
.A2(n_1706),
.B(n_1760),
.C(n_1665),
.Y(n_1878)
);

NAND2x1_ASAP7_75t_L g1879 ( 
.A(n_1868),
.B(n_1706),
.Y(n_1879)
);

AOI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1872),
.A2(n_1871),
.B(n_1873),
.C(n_1875),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1869),
.A2(n_1706),
.B1(n_1665),
.B2(n_1657),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1866),
.Y(n_1882)
);

CKINVDCx16_ASAP7_75t_R g1883 ( 
.A(n_1877),
.Y(n_1883)
);

OAI21xp33_ASAP7_75t_L g1884 ( 
.A1(n_1880),
.A2(n_1874),
.B(n_1876),
.Y(n_1884)
);

AOI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1878),
.A2(n_1882),
.B(n_1881),
.C(n_1879),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1880),
.A2(n_1710),
.B1(n_1702),
.B2(n_1712),
.C(n_1703),
.Y(n_1886)
);

O2A1O1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1880),
.A2(n_1665),
.B(n_1703),
.C(n_1701),
.Y(n_1887)
);

AOI31xp33_ASAP7_75t_L g1888 ( 
.A1(n_1880),
.A2(n_1551),
.A3(n_1528),
.B(n_1567),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1883),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1885),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1888),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1886),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1887),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1889),
.B(n_1884),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1889),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1890),
.Y(n_1896)
);

OR2x6_ASAP7_75t_L g1897 ( 
.A(n_1894),
.B(n_1891),
.Y(n_1897)
);

AOI31xp33_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1895),
.A3(n_1896),
.B(n_1893),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1898),
.B(n_1892),
.Y(n_1899)
);

AO22x2_ASAP7_75t_SL g1900 ( 
.A1(n_1898),
.A2(n_1701),
.B1(n_1708),
.B2(n_1705),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1900),
.B(n_1899),
.Y(n_1901)
);

OAI22x1_ASAP7_75t_L g1902 ( 
.A1(n_1899),
.A2(n_1712),
.B1(n_1710),
.B2(n_1702),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1901),
.Y(n_1903)
);

OAI21x1_ASAP7_75t_L g1904 ( 
.A1(n_1902),
.A2(n_1714),
.B(n_1713),
.Y(n_1904)
);

OAI21x1_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1713),
.B(n_1714),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1905),
.A2(n_1903),
.B1(n_1904),
.B2(n_1715),
.Y(n_1906)
);

XNOR2xp5_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1602),
.Y(n_1907)
);

OAI221xp5_ASAP7_75t_R g1908 ( 
.A1(n_1907),
.A2(n_1712),
.B1(n_1710),
.B2(n_1702),
.C(n_1721),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1555),
.B(n_1559),
.C(n_1567),
.Y(n_1909)
);


endmodule