module fake_netlist_6_3220_n_843 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_843);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_843;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_55),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_16),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_19),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_62),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_104),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_51),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_30),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_99),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_112),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_133),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_48),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_71),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_61),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_78),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_50),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_165),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_82),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_28),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_25),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_52),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_53),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_32),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_13),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_123),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_105),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_146),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_151),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_14),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_13),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_100),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_20),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_0),
.B(n_1),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_181),
.A2(n_0),
.B(n_1),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_227),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_230),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

OAI22x1_ASAP7_75t_SL g255 ( 
.A1(n_205),
.A2(n_235),
.B1(n_236),
.B2(n_210),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

BUFx8_ASAP7_75t_SL g258 ( 
.A(n_206),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_2),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_176),
.B(n_21),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_184),
.A2(n_2),
.B(n_3),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_185),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_174),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_215),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_195),
.A2(n_4),
.B(n_5),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_197),
.Y(n_273)
);

OAI22x1_ASAP7_75t_L g274 ( 
.A1(n_198),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_201),
.B(n_6),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_177),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_211),
.A2(n_216),
.B(n_212),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_218),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_8),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_206),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_180),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_258),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_270),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_270),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_277),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_277),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_287),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_251),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_269),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_253),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_263),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_269),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_288),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_R g315 ( 
.A(n_244),
.B(n_182),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_183),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_288),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_288),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_255),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_250),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_271),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_267),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_284),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_249),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_249),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_249),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_265),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_264),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_275),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_264),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_241),
.B(n_278),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_261),
.B1(n_274),
.B2(n_219),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_241),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_241),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_322),
.B(n_193),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_286),
.C(n_276),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_326),
.B(n_186),
.Y(n_349)
);

BUFx6f_ASAP7_75t_SL g350 ( 
.A(n_290),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_241),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_329),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_241),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_328),
.B(n_188),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

AO221x1_ASAP7_75t_L g356 ( 
.A1(n_338),
.A2(n_274),
.B1(n_257),
.B2(n_272),
.C(n_266),
.Y(n_356)
);

NOR2x1p5_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_189),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_278),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_244),
.C(n_264),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_314),
.B(n_203),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_259),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_313),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_338),
.A2(n_279),
.B1(n_244),
.B2(n_207),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_318),
.B(n_320),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_306),
.B(n_319),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_262),
.Y(n_370)
);

CKINVDCx11_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_312),
.B(n_295),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_259),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_259),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_292),
.B(n_279),
.Y(n_375)
);

NAND2x1_ASAP7_75t_L g376 ( 
.A(n_298),
.B(n_262),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_268),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_316),
.B(n_259),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_316),
.B(n_259),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_299),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_296),
.B(n_204),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_308),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_268),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_297),
.B(n_208),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_298),
.B(n_260),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_L g389 ( 
.A(n_321),
.B(n_202),
.C(n_266),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_300),
.B(n_273),
.C(n_268),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_301),
.B(n_209),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_298),
.B(n_260),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_310),
.B(n_268),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_333),
.B(n_260),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_260),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_307),
.B(n_273),
.Y(n_397)
);

NOR2x1p5_ASAP7_75t_L g398 ( 
.A(n_289),
.B(n_214),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_291),
.B(n_217),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_330),
.B(n_262),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_260),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_322),
.B(n_222),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_262),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_322),
.B(n_223),
.Y(n_406)
);

NOR2x1p5_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_225),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_324),
.B(n_285),
.C(n_282),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

NAND2x1_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_262),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_243),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_407),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_243),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_226),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_410),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_352),
.B(n_273),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_273),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_360),
.B(n_272),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

BUFx6f_ASAP7_75t_SL g426 ( 
.A(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_383),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_345),
.B(n_229),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_356),
.A2(n_285),
.B1(n_282),
.B2(n_252),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_359),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_359),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_358),
.B(n_240),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_359),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

BUFx4f_ASAP7_75t_SL g442 ( 
.A(n_399),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_370),
.A2(n_231),
.B1(n_232),
.B2(n_239),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_361),
.B(n_240),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_371),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_361),
.B(n_248),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_348),
.B(n_346),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_376),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_367),
.B(n_248),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_364),
.B(n_252),
.Y(n_454)
);

CKINVDCx11_ASAP7_75t_R g455 ( 
.A(n_364),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_363),
.B(n_282),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_363),
.B(n_282),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_389),
.A2(n_285),
.B1(n_252),
.B2(n_257),
.Y(n_460)
);

CKINVDCx12_ASAP7_75t_R g461 ( 
.A(n_350),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_341),
.A2(n_285),
.B1(n_257),
.B2(n_280),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_349),
.B(n_23),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_354),
.B(n_24),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_344),
.B(n_280),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_351),
.B(n_280),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_364),
.B(n_9),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

AO22x1_ASAP7_75t_L g473 ( 
.A1(n_343),
.A2(n_281),
.B1(n_280),
.B2(n_11),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_403),
.B(n_406),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_353),
.B(n_280),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_357),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_395),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_365),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_384),
.B(n_281),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_400),
.A2(n_281),
.B1(n_10),
.B2(n_11),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_398),
.B(n_387),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_393),
.B(n_26),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_447),
.A2(n_392),
.B1(n_350),
.B2(n_373),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_374),
.B1(n_281),
.B2(n_95),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_281),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_419),
.B(n_9),
.Y(n_490)
);

O2A1O1Ixp5_ASAP7_75t_L g491 ( 
.A1(n_418),
.A2(n_464),
.B(n_411),
.C(n_477),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_435),
.A2(n_94),
.B(n_172),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_12),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_415),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_417),
.A2(n_93),
.B1(n_170),
.B2(n_168),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_465),
.B(n_466),
.Y(n_497)
);

CKINVDCx8_ASAP7_75t_R g498 ( 
.A(n_431),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_422),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_27),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_412),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_446),
.A2(n_92),
.B(n_167),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_428),
.B(n_12),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_420),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_412),
.B(n_14),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_435),
.A2(n_96),
.B(n_166),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_465),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_SL g509 ( 
.A(n_476),
.B(n_15),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_453),
.A2(n_97),
.B(n_29),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_416),
.B(n_17),
.Y(n_512)
);

BUFx12f_ASAP7_75t_L g513 ( 
.A(n_455),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_424),
.B(n_31),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_33),
.C(n_34),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_453),
.A2(n_449),
.B(n_446),
.Y(n_517)
);

A2O1A1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_452),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_452),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_449),
.A2(n_41),
.B(n_42),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_430),
.B(n_43),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_454),
.B(n_44),
.Y(n_523)
);

OR2x6_ASAP7_75t_SL g524 ( 
.A(n_456),
.B(n_45),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_467),
.A2(n_46),
.B(n_47),
.C(n_49),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_425),
.B(n_54),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_470),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_454),
.B(n_482),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_418),
.A2(n_56),
.B(n_57),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_478),
.A2(n_58),
.B(n_59),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_448),
.B(n_63),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_472),
.B(n_64),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_457),
.A2(n_65),
.B(n_66),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_471),
.Y(n_534)
);

BUFx2_ASAP7_75t_SL g535 ( 
.A(n_426),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_454),
.B(n_67),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_466),
.B(n_68),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_471),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_457),
.A2(n_69),
.B(n_72),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_479),
.B(n_73),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_459),
.A2(n_74),
.B(n_75),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_459),
.A2(n_77),
.B(n_81),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_471),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_501),
.Y(n_544)
);

AOI22x1_ASAP7_75t_L g545 ( 
.A1(n_502),
.A2(n_451),
.B1(n_483),
.B2(n_479),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_517),
.A2(n_491),
.B(n_483),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_468),
.B(n_475),
.Y(n_547)
);

CKINVDCx8_ASAP7_75t_R g548 ( 
.A(n_534),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_488),
.A2(n_432),
.B(n_414),
.Y(n_549)
);

OAI21x1_ASAP7_75t_SL g550 ( 
.A1(n_532),
.A2(n_529),
.B(n_492),
.Y(n_550)
);

AO21x2_ASAP7_75t_L g551 ( 
.A1(n_490),
.A2(n_468),
.B(n_475),
.Y(n_551)
);

BUFx4f_ASAP7_75t_SL g552 ( 
.A(n_513),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_506),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_487),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_485),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

INVx3_ASAP7_75t_SL g557 ( 
.A(n_497),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_540),
.A2(n_469),
.B(n_444),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_538),
.Y(n_559)
);

INVx6_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

BUFx2_ASAP7_75t_SL g561 ( 
.A(n_498),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_511),
.A2(n_458),
.B(n_463),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_493),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_507),
.A2(n_530),
.B(n_506),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_495),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_499),
.A2(n_423),
.B(n_480),
.Y(n_566)
);

INVx5_ASAP7_75t_SL g567 ( 
.A(n_493),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_521),
.A2(n_445),
.B(n_438),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_503),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_504),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_528),
.Y(n_571)
);

AOI22x1_ASAP7_75t_L g572 ( 
.A1(n_522),
.A2(n_479),
.B1(n_443),
.B2(n_441),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_533),
.A2(n_445),
.B(n_439),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_539),
.A2(n_440),
.B(n_433),
.Y(n_574)
);

OA21x2_ASAP7_75t_L g575 ( 
.A1(n_527),
.A2(n_414),
.B(n_423),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_500),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_541),
.A2(n_434),
.B(n_481),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_510),
.B(n_442),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_515),
.B(n_437),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_505),
.B(n_442),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_500),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_526),
.Y(n_583)
);

NAND2x1p5_ASAP7_75t_L g584 ( 
.A(n_537),
.B(n_461),
.Y(n_584)
);

BUFx8_ASAP7_75t_L g585 ( 
.A(n_523),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_514),
.A2(n_462),
.B1(n_426),
.B2(n_460),
.Y(n_586)
);

BUFx2_ASAP7_75t_SL g587 ( 
.A(n_500),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_509),
.Y(n_588)
);

INVx3_ASAP7_75t_SL g589 ( 
.A(n_536),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_500),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_578),
.A2(n_489),
.B(n_519),
.Y(n_591)
);

BUFx2_ASAP7_75t_R g592 ( 
.A(n_561),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_588),
.A2(n_508),
.B1(n_494),
.B2(n_520),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

OA21x2_ASAP7_75t_L g595 ( 
.A1(n_546),
.A2(n_545),
.B(n_564),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_553),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_557),
.A2(n_520),
.B1(n_524),
.B2(n_486),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_562),
.A2(n_542),
.B(n_496),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_557),
.A2(n_583),
.B1(n_586),
.B2(n_569),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_544),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_555),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_575),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_590),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_565),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_570),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_574),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_577),
.B(n_518),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_580),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_554),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_571),
.A2(n_516),
.B1(n_512),
.B2(n_531),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_577),
.B(n_525),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_556),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_550),
.A2(n_473),
.B(n_484),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_581),
.A2(n_484),
.B1(n_85),
.B2(n_86),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_568),
.A2(n_549),
.B(n_573),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_583),
.A2(n_484),
.B1(n_87),
.B2(n_88),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_549),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_556),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_588),
.A2(n_484),
.B1(n_89),
.B2(n_90),
.Y(n_622)
);

CKINVDCx6p67_ASAP7_75t_R g623 ( 
.A(n_589),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_572),
.A2(n_84),
.B(n_98),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_560),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx6_ASAP7_75t_L g627 ( 
.A(n_576),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_581),
.B(n_101),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_569),
.A2(n_589),
.B1(n_584),
.B2(n_579),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_579),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_560),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_566),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_584),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_600),
.B(n_559),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_601),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g636 ( 
.A1(n_618),
.A2(n_582),
.B(n_587),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_R g637 ( 
.A(n_600),
.B(n_552),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_610),
.B(n_563),
.Y(n_638)
);

AO31x2_ASAP7_75t_L g639 ( 
.A1(n_607),
.A2(n_547),
.A3(n_551),
.B(n_576),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_605),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_623),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_594),
.B(n_567),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_599),
.B(n_567),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_548),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_567),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_609),
.B(n_543),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_592),
.Y(n_647)
);

CKINVDCx16_ASAP7_75t_R g648 ( 
.A(n_610),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_585),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_597),
.B(n_547),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_613),
.A2(n_543),
.B1(n_585),
.B2(n_590),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g652 ( 
.A(n_612),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_606),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_596),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_611),
.B(n_543),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_SL g656 ( 
.A1(n_619),
.A2(n_590),
.B(n_558),
.C(n_560),
.Y(n_656)
);

CKINVDCx16_ASAP7_75t_R g657 ( 
.A(n_612),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_SL g658 ( 
.A(n_630),
.B(n_552),
.C(n_590),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_615),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_621),
.B(n_558),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_620),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_111),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_603),
.B(n_114),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_R g664 ( 
.A(n_603),
.B(n_115),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_631),
.B(n_116),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_R g666 ( 
.A(n_614),
.B(n_117),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_614),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_122),
.Y(n_668)
);

AO31x2_ASAP7_75t_L g669 ( 
.A1(n_607),
.A2(n_124),
.A3(n_125),
.B(n_127),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_603),
.B(n_129),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_R g671 ( 
.A(n_603),
.B(n_130),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_602),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_608),
.B(n_614),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_625),
.B(n_132),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_622),
.A2(n_608),
.B1(n_603),
.B2(n_624),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_608),
.B(n_134),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_617),
.A2(n_173),
.B1(n_137),
.B2(n_138),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_602),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_136),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_627),
.B(n_139),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_591),
.B(n_141),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_604),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_673),
.B(n_626),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_661),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_660),
.B(n_632),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_672),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_673),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_678),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_682),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_634),
.B(n_644),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_650),
.B(n_632),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_639),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_643),
.B(n_626),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_650),
.B(n_604),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_648),
.B(n_627),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_673),
.B(n_595),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_636),
.B(n_624),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_659),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_639),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_635),
.B(n_640),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_653),
.B(n_595),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_654),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_639),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_SL g704 ( 
.A1(n_649),
.A2(n_627),
.B1(n_616),
.B2(n_144),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_681),
.B(n_598),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_676),
.B(n_598),
.Y(n_706)
);

AOI211xp5_ASAP7_75t_L g707 ( 
.A1(n_679),
.A2(n_616),
.B(n_143),
.C(n_145),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_651),
.B(n_627),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_638),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_669),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_669),
.B(n_142),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_669),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_645),
.B(n_164),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_676),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_663),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_652),
.B(n_149),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_663),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_667),
.B(n_153),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_656),
.Y(n_719)
);

NOR4xp25_ASAP7_75t_SL g720 ( 
.A(n_666),
.B(n_647),
.C(n_658),
.D(n_664),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_SL g721 ( 
.A1(n_718),
.A2(n_651),
.B(n_667),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_694),
.B(n_675),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_698),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_694),
.B(n_685),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_686),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_686),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_688),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_700),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_700),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_714),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_688),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_707),
.A2(n_677),
.B1(n_704),
.B2(n_716),
.C(n_708),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_714),
.B(n_657),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_687),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_689),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_691),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_689),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_690),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_718),
.B(n_675),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_701),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_687),
.B(n_646),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_687),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_685),
.B(n_642),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_691),
.B(n_662),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_696),
.B(n_655),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_709),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_696),
.B(n_668),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_687),
.B(n_638),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_701),
.B(n_674),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_718),
.A2(n_677),
.B1(n_658),
.B2(n_641),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_693),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_739),
.B(n_687),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_725),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_745),
.B(n_683),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_730),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_726),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_739),
.B(n_718),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_745),
.B(n_709),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_724),
.B(n_683),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_734),
.B(n_683),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_736),
.B(n_706),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_724),
.B(n_683),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_723),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_722),
.B(n_692),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_751),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_744),
.B(n_706),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_722),
.B(n_703),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_731),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_735),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_684),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_740),
.B(n_703),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_737),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_738),
.B(n_705),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_727),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_757),
.A2(n_721),
.B1(n_732),
.B2(n_750),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_771),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_753),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_759),
.B(n_747),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_765),
.B(n_743),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_774),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_759),
.B(n_747),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_756),
.Y(n_782)
);

NOR2x1_ASAP7_75t_L g783 ( 
.A(n_763),
.B(n_719),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_771),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_757),
.A2(n_752),
.B1(n_748),
.B2(n_741),
.Y(n_785)
);

OAI32xp33_ASAP7_75t_L g786 ( 
.A1(n_752),
.A2(n_733),
.A3(n_716),
.B1(n_719),
.B2(n_729),
.Y(n_786)
);

O2A1O1Ixp5_ASAP7_75t_R g787 ( 
.A1(n_773),
.A2(n_720),
.B(n_743),
.C(n_746),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_762),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_762),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_777),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_775),
.A2(n_748),
.B1(n_741),
.B2(n_746),
.Y(n_791)
);

OA22x2_ASAP7_75t_L g792 ( 
.A1(n_785),
.A2(n_764),
.B1(n_767),
.B2(n_758),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_778),
.B(n_754),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_787),
.A2(n_748),
.B1(n_741),
.B2(n_760),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_786),
.A2(n_711),
.B(n_770),
.C(n_755),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_790),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_795),
.B(n_779),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_792),
.B(n_783),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_791),
.B(n_779),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_794),
.A2(n_760),
.B1(n_713),
.B2(n_695),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_793),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_SL g802 ( 
.A(n_797),
.B(n_637),
.C(n_711),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_801),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_796),
.Y(n_804)
);

AOI221x1_ASAP7_75t_L g805 ( 
.A1(n_799),
.A2(n_782),
.B1(n_769),
.B2(n_772),
.C(n_768),
.Y(n_805)
);

INVxp33_ASAP7_75t_L g806 ( 
.A(n_802),
.Y(n_806)
);

NOR2x1_ASAP7_75t_L g807 ( 
.A(n_804),
.B(n_798),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_803),
.B(n_800),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_R g809 ( 
.A(n_808),
.B(n_713),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_806),
.A2(n_805),
.B(n_680),
.C(n_780),
.Y(n_810)
);

NOR3x1_ASAP7_75t_L g811 ( 
.A(n_807),
.B(n_742),
.C(n_789),
.Y(n_811)
);

AOI211xp5_ASAP7_75t_L g812 ( 
.A1(n_806),
.A2(n_680),
.B(n_671),
.C(n_766),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_812),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_810),
.A2(n_742),
.B1(n_734),
.B2(n_760),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_809),
.B(n_780),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_811),
.B(n_788),
.Y(n_816)
);

NOR2x1p5_ASAP7_75t_L g817 ( 
.A(n_809),
.B(n_734),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_812),
.A2(n_767),
.B1(n_764),
.B2(n_749),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_817),
.Y(n_819)
);

XNOR2xp5_ASAP7_75t_L g820 ( 
.A(n_813),
.B(n_665),
.Y(n_820)
);

OAI222xp33_ASAP7_75t_L g821 ( 
.A1(n_814),
.A2(n_776),
.B1(n_784),
.B2(n_670),
.C1(n_710),
.C2(n_705),
.Y(n_821)
);

AND4x1_ASAP7_75t_L g822 ( 
.A(n_816),
.B(n_781),
.C(n_754),
.D(n_749),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_815),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_823),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_819),
.A2(n_818),
.B1(n_784),
.B2(n_776),
.Y(n_825)
);

AND3x4_ASAP7_75t_L g826 ( 
.A(n_822),
.B(n_670),
.C(n_715),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_820),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_824),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_825),
.A2(n_821),
.B1(n_717),
.B2(n_710),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_827),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_826),
.A2(n_821),
.B1(n_717),
.B2(n_728),
.Y(n_831)
);

HB1xp67_ASAP7_75t_SL g832 ( 
.A(n_824),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_832),
.Y(n_833)
);

AOI31xp33_ASAP7_75t_L g834 ( 
.A1(n_830),
.A2(n_715),
.A3(n_761),
.B(n_712),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_828),
.A2(n_717),
.B1(n_712),
.B2(n_699),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_829),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_SL g837 ( 
.A1(n_833),
.A2(n_831),
.B1(n_727),
.B2(n_702),
.Y(n_837)
);

INVxp33_ASAP7_75t_L g838 ( 
.A(n_835),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_837),
.A2(n_836),
.B1(n_834),
.B2(n_697),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_839),
.B(n_838),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_SL g841 ( 
.A1(n_840),
.A2(n_697),
.B1(n_692),
.B2(n_699),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_841),
.B(n_154),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_842),
.A2(n_155),
.B1(n_156),
.B2(n_161),
.Y(n_843)
);


endmodule