module fake_jpeg_31745_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_18),
.B1(n_2),
.B2(n_14),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_11),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_19),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_16),
.B1(n_18),
.B2(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_20),
.B(n_22),
.C(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_24),
.B(n_28),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_37),
.C(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_30),
.B1(n_32),
.B2(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_36),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_43),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_38),
.B(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.A3(n_24),
.B1(n_21),
.B2(n_13),
.C1(n_9),
.C2(n_0),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_13),
.B(n_0),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_49),
.B(n_0),
.Y(n_51)
);


endmodule