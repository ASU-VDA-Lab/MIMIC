module real_jpeg_11085_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_288;
wire n_176;
wire n_221;
wire n_166;
wire n_249;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_1),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_44),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_3),
.A2(n_27),
.B1(n_54),
.B2(n_55),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_68),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_70),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_7),
.B(n_25),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_140),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_3),
.A2(n_8),
.B(n_54),
.C(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_4),
.A2(n_10),
.B1(n_68),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_4),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_80),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_80),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_4),
.A2(n_41),
.B1(n_43),
.B2(n_80),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_7),
.A2(n_38),
.B(n_41),
.C(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_7),
.B(n_41),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_8),
.A2(n_41),
.B1(n_43),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_54),
.B(n_56),
.C(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_54),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_11),
.B1(n_33),
.B2(n_68),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_33),
.B1(n_41),
.B2(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_33),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_122),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_103),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_16),
.B(n_103),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_81),
.C(n_90),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_17),
.A2(n_18),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.C(n_63),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_19),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_20),
.B(n_36),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_21),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_22),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_23),
.A2(n_34),
.B(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_24),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_27),
.A2(n_39),
.B(n_43),
.C(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_27),
.B(n_37),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_27),
.B(n_35),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_27),
.A2(n_41),
.B(n_57),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_28),
.B(n_32),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_28),
.B(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_29),
.A2(n_35),
.B(n_130),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_30),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_34),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_34),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_45),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_37),
.A2(n_95),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_38),
.B(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_38),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_40),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_45),
.B(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_47),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_47),
.B(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_49),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_60),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_52),
.B(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_55),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_54),
.B(n_73),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_55),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_56),
.A2(n_61),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_58),
.B(n_139),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_59),
.B(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_59),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_61),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_71),
.B(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_67),
.B(n_76),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_71),
.B(n_72),
.C(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_72),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_69),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_79),
.Y(n_136)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_76),
.B(n_109),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_77),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_81),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_89),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_83),
.B(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_139),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_104),
.CI(n_120),
.CON(n_103),
.SN(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_93),
.A2(n_98),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_93),
.B(n_221),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_96),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_100),
.B(n_102),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_103),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_112),
.B2(n_113),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_135),
.C(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_115),
.B1(n_137),
.B2(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_283),
.B(n_289),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_271),
.B(n_282),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_176),
.B(n_253),
.C(n_270),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_162),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_126),
.B(n_162),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_142),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_128),
.B(n_134),
.C(n_142),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_129),
.B(n_132),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_133),
.B(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_136),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_152),
.B1(n_153),
.B2(n_161),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_151),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_144),
.B(n_151),
.C(n_152),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_163),
.A2(n_164),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.C(n_172),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_170),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_171),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_252),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_246),
.B(n_251),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_232),
.B(n_245),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_217),
.B(n_231),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_206),
.B(n_216),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_195),
.B(n_205),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_187),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_191),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_200),
.B(n_204),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_219),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_224),
.B1(n_225),
.B2(n_230),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_229),
.C(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_241),
.C(n_244),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_241),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_255),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_268),
.B2(n_269),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_259),
.C(n_269),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_281),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_279),
.C(n_281),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule