module fake_jpeg_5345_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_5),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_7),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_34),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_17),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_7),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_29),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_59),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_51),
.A2(n_54),
.B1(n_74),
.B2(n_76),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_63),
.Y(n_104)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_66),
.Y(n_112)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_19),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_29),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_39),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_27),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_87),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_27),
.C(n_15),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_59),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_92),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_39),
.A2(n_35),
.B1(n_26),
.B2(n_18),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_37),
.B(n_35),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_39),
.A2(n_26),
.B1(n_18),
.B2(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_27),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_15),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_100),
.B(n_111),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_59),
.B(n_15),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_117),
.B(n_54),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_124),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_58),
.A2(n_26),
.B(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_57),
.B(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_57),
.Y(n_153)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_65),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_138),
.B(n_160),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_134),
.B(n_139),
.Y(n_192)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

AO21x2_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_84),
.B(n_51),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_154),
.B1(n_120),
.B2(n_109),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_89),
.B1(n_95),
.B2(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_152),
.B1(n_163),
.B2(n_105),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_141),
.B(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_142),
.B(n_146),
.Y(n_198)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_101),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_78),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_122),
.B1(n_119),
.B2(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_SL g193 ( 
.A(n_153),
.B(n_83),
.C(n_67),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_90),
.B1(n_91),
.B2(n_56),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_62),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_159),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_61),
.B1(n_77),
.B2(n_70),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_62),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_138),
.C(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_191),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_168),
.B1(n_174),
.B2(n_197),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_105),
.B1(n_115),
.B2(n_120),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_194),
.B1(n_196),
.B2(n_65),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_107),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_53),
.C(n_128),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_107),
.B1(n_56),
.B2(n_79),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_187),
.B(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_195),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_133),
.A2(n_107),
.B(n_86),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_142),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_154),
.B1(n_152),
.B2(n_140),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_159),
.B1(n_139),
.B2(n_134),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_52),
.B1(n_66),
.B2(n_63),
.Y(n_197)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_128),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_208),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_129),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_211),
.B(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_136),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_131),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_145),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_0),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_198),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_17),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_0),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_225),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_170),
.B(n_10),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_53),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_222),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_128),
.C(n_0),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_190),
.B(n_13),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_1),
.B(n_3),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_219),
.B(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_167),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_212),
.C(n_225),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_182),
.Y(n_236)
);

AO32x1_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_201),
.A3(n_214),
.B1(n_209),
.B2(n_203),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_175),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_184),
.Y(n_262)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_185),
.B1(n_194),
.B2(n_189),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_202),
.B1(n_205),
.B2(n_215),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_194),
.B1(n_189),
.B2(n_192),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_193),
.C(n_170),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_247),
.C(n_176),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_248),
.A2(n_226),
.B1(n_246),
.B2(n_233),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_255),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_257),
.B(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_220),
.C(n_203),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_254),
.C(n_231),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_201),
.C(n_222),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_211),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_213),
.B(n_200),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_223),
.B1(n_186),
.B2(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_210),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_197),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_262),
.B(n_263),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_199),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_249),
.C(n_259),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_247),
.B(n_230),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_172),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_275),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_230),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_240),
.B1(n_226),
.B2(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_233),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_250),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_283),
.B(n_288),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_253),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_281),
.C(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_260),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_246),
.C(n_242),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_280),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_271),
.B(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_237),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_294),
.B(n_265),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_237),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_276),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_296),
.B(n_272),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_299),
.B(n_302),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_297),
.B(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_245),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_307),
.B(n_195),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_295),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_303),
.A3(n_281),
.B1(n_228),
.B2(n_297),
.C1(n_171),
.C2(n_184),
.Y(n_308)
);

AOI321xp33_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_309),
.A3(n_228),
.B1(n_304),
.B2(n_171),
.C(n_6),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_1),
.Y(n_311)
);


endmodule