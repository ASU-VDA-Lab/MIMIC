module fake_jpeg_25804_n_253 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_52),
.Y(n_76)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_59),
.Y(n_93)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_15),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_2),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_37),
.C(n_27),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_65),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_24),
.B1(n_37),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_63),
.A2(n_71),
.B1(n_29),
.B2(n_22),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_37),
.C(n_20),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_77),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_24),
.B1(n_36),
.B2(n_34),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_78),
.A3(n_40),
.B1(n_45),
.B2(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_91),
.B(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_30),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_34),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_31),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_99),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_21),
.B(n_31),
.C(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_51),
.B1(n_50),
.B2(n_30),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_120),
.B1(n_123),
.B2(n_80),
.Y(n_138)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_111),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_30),
.B(n_29),
.C(n_22),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_117),
.C(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_29),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_118),
.Y(n_132)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_3),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_93),
.C(n_62),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_145),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_67),
.B1(n_75),
.B2(n_72),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_65),
.B1(n_93),
.B2(n_67),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_142),
.B1(n_150),
.B2(n_103),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_72),
.B1(n_90),
.B2(n_81),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_61),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_108),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_61),
.B1(n_45),
.B2(n_40),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_105),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_74),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_96),
.B(n_110),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_74),
.B1(n_76),
.B2(n_5),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_99),
.B1(n_116),
.B2(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_96),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_157),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_121),
.B1(n_119),
.B2(n_113),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_162),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_113),
.B1(n_118),
.B2(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_115),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_94),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_101),
.B1(n_100),
.B2(n_95),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_130),
.B1(n_141),
.B2(n_124),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_117),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_3),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_170),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_173),
.B1(n_143),
.B2(n_128),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_150),
.B1(n_127),
.B2(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_14),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_12),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_133),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_182),
.B(n_193),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_130),
.B1(n_141),
.B2(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_174),
.B1(n_165),
.B2(n_159),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_132),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_143),
.B1(n_139),
.B2(n_126),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_12),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_194),
.Y(n_201)
);

OAI322xp33_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_166),
.A3(n_174),
.B1(n_153),
.B2(n_154),
.C1(n_170),
.C2(n_173),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_178),
.C(n_189),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_199),
.B(n_208),
.Y(n_213)
);

AOI221xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_174),
.B1(n_155),
.B2(n_165),
.C(n_153),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_200),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_163),
.B1(n_153),
.B2(n_171),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_166),
.A3(n_151),
.B1(n_163),
.B2(n_167),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_175),
.C(n_152),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_207),
.C(n_181),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_127),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_139),
.B(n_126),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_179),
.B(n_177),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_222),
.Y(n_231)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_217),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_183),
.B1(n_181),
.B2(n_180),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_219),
.B1(n_204),
.B2(n_198),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_183),
.B1(n_182),
.B2(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_221),
.A2(n_204),
.B1(n_200),
.B2(n_210),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_207),
.C(n_206),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_228),
.C(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_226),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_210),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_200),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_220),
.C(n_213),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_216),
.B(n_213),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_234),
.B(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_236),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_214),
.B(n_219),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_215),
.C(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_211),
.Y(n_238)
);

OAI221xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_201),
.B1(n_176),
.B2(n_178),
.C(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_176),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_242),
.B(n_194),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_227),
.B(n_229),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_191),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_239),
.A2(n_233),
.B(n_228),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_225),
.C(n_13),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_249),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_13),
.Y(n_253)
);


endmodule