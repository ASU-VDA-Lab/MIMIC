module real_aes_14235_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_723, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_723;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g569 ( .A(n_0), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_0), .A2(n_46), .B1(n_636), .B2(n_647), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_1), .Y(n_658) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_2), .A2(n_41), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g169 ( .A(n_2), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_3), .B(n_198), .Y(n_270) );
INVx1_ASAP7_75t_L g659 ( .A(n_3), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_4), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g711 ( .A(n_4), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_5), .B(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g497 ( .A(n_6), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_7), .B(n_156), .Y(n_205) );
INVx3_ASAP7_75t_L g542 ( .A(n_8), .Y(n_542) );
INVx1_ASAP7_75t_L g501 ( .A(n_9), .Y(n_501) );
INVx2_ASAP7_75t_L g513 ( .A(n_9), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_10), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_11), .B(n_145), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_12), .B(n_269), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_13), .Y(n_185) );
INVx1_ASAP7_75t_L g533 ( .A(n_14), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_14), .A2(n_63), .B1(n_590), .B2(n_594), .Y(n_589) );
INVx1_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
BUFx3_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_16), .B(n_220), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_17), .Y(n_143) );
BUFx10_ASAP7_75t_L g686 ( .A(n_18), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_19), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g669 ( .A(n_20), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_21), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_22), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_23), .B(n_238), .Y(n_241) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_24), .Y(n_667) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_25), .Y(n_585) );
INVx1_ASAP7_75t_L g609 ( .A(n_25), .Y(n_609) );
INVxp33_ASAP7_75t_L g622 ( .A(n_25), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_26), .B(n_220), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g273 ( .A(n_27), .B(n_157), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_28), .A2(n_175), .B(n_177), .C(n_179), .Y(n_174) );
INVx1_ASAP7_75t_L g88 ( .A(n_29), .Y(n_88) );
INVx2_ASAP7_75t_L g549 ( .A(n_30), .Y(n_549) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_31), .A2(n_522), .B(n_526), .Y(n_521) );
INVx1_ASAP7_75t_L g576 ( .A(n_31), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_32), .B(n_224), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_33), .B(n_92), .Y(n_119) );
INVx1_ASAP7_75t_L g664 ( .A(n_33), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_34), .B(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_35), .Y(n_551) );
INVx2_ASAP7_75t_L g556 ( .A(n_35), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_35), .B(n_609), .Y(n_608) );
AO221x1_ASAP7_75t_L g245 ( .A1(n_36), .A2(n_65), .B1(n_187), .B2(n_238), .C(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_37), .B(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_37), .Y(n_721) );
AND2x4_ASAP7_75t_L g87 ( .A(n_38), .B(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_38), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g225 ( .A(n_39), .B(n_179), .C(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g500 ( .A(n_40), .Y(n_500) );
INVx1_ASAP7_75t_L g512 ( .A(n_40), .Y(n_512) );
INVx1_ASAP7_75t_L g168 ( .A(n_41), .Y(n_168) );
INVx1_ASAP7_75t_L g131 ( .A(n_42), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g109 ( .A1(n_43), .A2(n_110), .B(n_112), .C(n_114), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_44), .Y(n_183) );
INVx2_ASAP7_75t_L g113 ( .A(n_45), .Y(n_113) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_46), .A2(n_74), .B1(n_601), .B2(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_47), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g529 ( .A(n_48), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g699 ( .A(n_49), .B(n_489), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_50), .B(n_200), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_51), .A2(n_76), .B1(n_594), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_51), .A2(n_69), .B1(n_626), .B2(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g670 ( .A(n_52), .Y(n_670) );
AND2x2_ASAP7_75t_L g206 ( .A(n_53), .B(n_160), .Y(n_206) );
INVx1_ASAP7_75t_L g254 ( .A(n_54), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_55), .A2(n_63), .B1(n_494), .B2(n_502), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_55), .A2(n_64), .B1(n_596), .B2(n_599), .Y(n_595) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_56), .Y(n_661) );
OAI222xp33_ASAP7_75t_L g544 ( .A1(n_57), .A2(n_58), .B1(n_69), .B2(n_545), .C1(n_552), .C2(n_559), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_57), .A2(n_76), .B1(n_633), .B2(n_636), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_58), .A2(n_74), .B1(n_626), .B2(n_629), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g250 ( .A1(n_59), .A2(n_62), .B1(n_121), .B2(n_198), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_60), .B(n_179), .Y(n_222) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_61), .A2(n_64), .B1(n_506), .B2(n_514), .C(n_520), .Y(n_505) );
OAI211xp5_ASAP7_75t_L g566 ( .A1(n_61), .A2(n_567), .B(n_568), .C(n_580), .Y(n_566) );
AND2x2_ASAP7_75t_L g127 ( .A(n_66), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
INVx1_ASAP7_75t_L g116 ( .A(n_67), .Y(n_116) );
BUFx3_ASAP7_75t_L g151 ( .A(n_67), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_68), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_70), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g548 ( .A(n_71), .Y(n_548) );
AND2x2_ASAP7_75t_L g558 ( .A(n_71), .B(n_549), .Y(n_558) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_71), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_72), .B(n_148), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_73), .B(n_160), .Y(n_274) );
INVx2_ASAP7_75t_L g539 ( .A(n_75), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_77), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_98), .B(n_487), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
BUFx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_89), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_84), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx3_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
BUFx6f_ASAP7_75t_SL g158 ( .A(n_87), .Y(n_158) );
INVx2_ASAP7_75t_L g172 ( .A(n_87), .Y(n_172) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_88), .Y(n_682) );
AO21x2_ASAP7_75t_L g718 ( .A1(n_89), .A2(n_707), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g111 ( .A(n_93), .Y(n_111) );
INVx2_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
INVx2_ASAP7_75t_L g226 ( .A(n_93), .Y(n_226) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
INVx2_ASAP7_75t_SL g95 ( .A(n_96), .Y(n_95) );
AOI21xp5_ASAP7_75t_SL g196 ( .A1(n_96), .A2(n_197), .B(n_199), .Y(n_196) );
BUFx3_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g126 ( .A(n_97), .Y(n_126) );
INVxp67_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
NAND4xp75_ASAP7_75t_L g100 ( .A(n_101), .B(n_386), .C(n_439), .D(n_473), .Y(n_100) );
AND4x1_ASAP7_75t_L g101 ( .A(n_102), .B(n_309), .C(n_342), .D(n_364), .Y(n_101) );
NOR2xp33_ASAP7_75t_SL g102 ( .A(n_103), .B(n_278), .Y(n_102) );
OAI222xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_212), .B1(n_256), .B2(n_259), .C1(n_275), .C2(n_723), .Y(n_103) );
NOR2x1_ASAP7_75t_L g104 ( .A(n_105), .B(n_207), .Y(n_104) );
NOR2x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_161), .Y(n_105) );
OR2x2_ASAP7_75t_L g256 ( .A(n_106), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_137), .Y(n_106) );
INVx1_ASAP7_75t_L g281 ( .A(n_107), .Y(n_281) );
OR2x2_ASAP7_75t_L g418 ( .A(n_107), .B(n_163), .Y(n_418) );
AND2x2_ASAP7_75t_L g429 ( .A(n_107), .B(n_163), .Y(n_429) );
AND2x2_ASAP7_75t_L g470 ( .A(n_107), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g211 ( .A(n_108), .Y(n_211) );
AND2x2_ASAP7_75t_L g293 ( .A(n_108), .B(n_163), .Y(n_293) );
INVx1_ASAP7_75t_L g307 ( .A(n_108), .Y(n_307) );
OR2x2_ASAP7_75t_L g321 ( .A(n_108), .B(n_192), .Y(n_321) );
AND2x2_ASAP7_75t_L g332 ( .A(n_108), .B(n_191), .Y(n_332) );
AND2x2_ASAP7_75t_L g354 ( .A(n_108), .B(n_190), .Y(n_354) );
AO21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_117), .B(n_132), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_110), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_111), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_115), .A2(n_272), .B(n_273), .Y(n_271) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g249 ( .A(n_116), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_127), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_121), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g269 ( .A(n_122), .Y(n_269) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_125), .A2(n_153), .B(n_155), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_125), .A2(n_203), .B(n_205), .Y(n_202) );
BUFx10_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI21xp33_ASAP7_75t_L g132 ( .A1(n_127), .A2(n_133), .B(n_135), .Y(n_132) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx2_ASAP7_75t_L g134 ( .A(n_130), .Y(n_134) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
INVx1_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_133), .B(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx3_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
AND2x4_ASAP7_75t_L g194 ( .A(n_135), .B(n_195), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_135), .A2(n_267), .B(n_271), .Y(n_266) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_136), .B(n_160), .Y(n_243) );
NOR2xp33_ASAP7_75t_R g251 ( .A(n_136), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g210 ( .A(n_137), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g282 ( .A(n_137), .B(n_164), .Y(n_282) );
OR2x2_ASAP7_75t_L g317 ( .A(n_137), .B(n_190), .Y(n_317) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g277 ( .A(n_138), .Y(n_277) );
AND2x2_ASAP7_75t_L g297 ( .A(n_138), .B(n_192), .Y(n_297) );
INVx1_ASAP7_75t_L g370 ( .A(n_138), .Y(n_370) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g308 ( .A(n_139), .B(n_192), .Y(n_308) );
INVxp33_ASAP7_75t_L g471 ( .A(n_139), .Y(n_471) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_159), .Y(n_139) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_152), .B(n_158), .Y(n_141) );
O2A1O1Ixp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_147), .C(n_150), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_145), .B(n_185), .Y(n_184) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_146), .Y(n_238) );
INVx2_ASAP7_75t_SL g200 ( .A(n_148), .Y(n_200) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g198 ( .A(n_149), .Y(n_198) );
INVx2_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_150), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_150), .A2(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx2_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
INVx2_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
INVx3_ASAP7_75t_L g246 ( .A(n_157), .Y(n_246) );
INVx2_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_160), .Y(n_234) );
INVx1_ASAP7_75t_L g265 ( .A(n_160), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_190), .Y(n_161) );
BUFx2_ASAP7_75t_SL g335 ( .A(n_162), .Y(n_335) );
INVx2_ASAP7_75t_L g384 ( .A(n_162), .Y(n_384) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_164), .B(n_307), .Y(n_306) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_173), .B(n_180), .Y(n_164) );
AO21x1_ASAP7_75t_SL g258 ( .A1(n_165), .A2(n_173), .B(n_180), .Y(n_258) );
INVxp67_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
OAI21x1_ASAP7_75t_SL g180 ( .A1(n_166), .A2(n_181), .B(n_188), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
INVx2_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .Y(n_167) );
AOI21x1_ASAP7_75t_L g252 ( .A1(n_168), .A2(n_169), .B(n_170), .Y(n_252) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_184), .B(n_186), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_186), .A2(n_237), .B(n_239), .Y(n_236) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_190), .B(n_211), .Y(n_385) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g209 ( .A(n_192), .Y(n_209) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
NAND2x1_ASAP7_75t_L g193 ( .A(n_194), .B(n_196), .Y(n_193) );
AOI21x1_ASAP7_75t_L g201 ( .A1(n_194), .A2(n_202), .B(n_206), .Y(n_201) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_194), .A2(n_217), .B(n_221), .C(n_227), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_207), .A2(n_461), .B1(n_485), .B2(n_486), .Y(n_484) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g276 ( .A(n_209), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_210), .Y(n_485) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_212), .A2(n_325), .B1(n_330), .B2(n_331), .Y(n_324) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_229), .Y(n_213) );
NOR2x1_ASAP7_75t_L g303 ( .A(n_214), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g346 ( .A(n_214), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_214), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g452 ( .A(n_214), .B(n_291), .Y(n_452) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_SL g260 ( .A(n_215), .Y(n_260) );
AND2x2_ASAP7_75t_L g287 ( .A(n_215), .B(n_263), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_215), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g328 ( .A(n_215), .Y(n_328) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_225), .Y(n_221) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g329 ( .A(n_229), .Y(n_329) );
AND2x2_ASAP7_75t_L g372 ( .A(n_229), .B(n_314), .Y(n_372) );
AND2x4_ASAP7_75t_L g382 ( .A(n_229), .B(n_287), .Y(n_382) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_244), .Y(n_229) );
INVx2_ASAP7_75t_L g302 ( .A(n_230), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_230), .B(n_328), .Y(n_339) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g291 ( .A(n_231), .B(n_263), .Y(n_291) );
OR2x2_ASAP7_75t_L g304 ( .A(n_231), .B(n_244), .Y(n_304) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_231), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_231), .B(n_263), .Y(n_376) );
AND2x2_ASAP7_75t_L g420 ( .A(n_231), .B(n_262), .Y(n_420) );
AND2x4_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_240), .B(n_243), .Y(n_235) );
OR2x2_ASAP7_75t_L g261 ( .A(n_244), .B(n_262), .Y(n_261) );
BUFx3_ASAP7_75t_L g285 ( .A(n_244), .Y(n_285) );
INVx2_ASAP7_75t_SL g290 ( .A(n_244), .Y(n_290) );
AND2x2_ASAP7_75t_L g359 ( .A(n_244), .B(n_302), .Y(n_359) );
AND2x2_ASAP7_75t_L g377 ( .A(n_244), .B(n_328), .Y(n_377) );
AND2x2_ASAP7_75t_L g421 ( .A(n_244), .B(n_327), .Y(n_421) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .A3(n_251), .B(n_253), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_268), .B(n_270), .Y(n_267) );
INVx2_ASAP7_75t_L g255 ( .A(n_252), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_257), .B(n_276), .Y(n_275) );
INVx5_ASAP7_75t_L g316 ( .A(n_257), .Y(n_316) );
AND2x2_ASAP7_75t_L g347 ( .A(n_257), .B(n_285), .Y(n_347) );
AND2x2_ASAP7_75t_L g389 ( .A(n_257), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g451 ( .A(n_257), .B(n_354), .Y(n_451) );
AND2x4_ASAP7_75t_SL g458 ( .A(n_257), .B(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVxp67_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_259), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NOR2x1_ASAP7_75t_SL g434 ( .A(n_260), .B(n_261), .Y(n_434) );
AND2x2_ASAP7_75t_L g476 ( .A(n_260), .B(n_291), .Y(n_476) );
OR2x2_ASAP7_75t_L g414 ( .A(n_261), .B(n_339), .Y(n_414) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
INVx1_ASAP7_75t_L g338 ( .A(n_263), .Y(n_338) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B(n_274), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OAI33xp33_ASAP7_75t_L g333 ( .A1(n_276), .A2(n_286), .A3(n_334), .B1(n_336), .B2(n_340), .B3(n_341), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_276), .B(n_316), .Y(n_340) );
INVx1_ASAP7_75t_L g438 ( .A(n_276), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_276), .A2(n_474), .B(n_477), .Y(n_473) );
OR2x2_ASAP7_75t_L g362 ( .A(n_277), .B(n_321), .Y(n_362) );
INVx1_ASAP7_75t_L g402 ( .A(n_277), .Y(n_402) );
OAI221xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_283), .B1(n_288), .B2(n_292), .C(n_294), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_280), .A2(n_446), .B1(n_449), .B2(n_452), .Y(n_445) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_281), .B(n_379), .Y(n_444) );
OAI321xp33_ASAP7_75t_L g477 ( .A1(n_281), .A2(n_379), .A3(n_478), .B1(n_480), .B2(n_481), .C(n_484), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_282), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g437 ( .A(n_282), .Y(n_437) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_285), .B(n_291), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_285), .A2(n_388), .B(n_391), .C(n_394), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_285), .B(n_379), .C(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_285), .Y(n_404) );
INVx2_ASAP7_75t_L g427 ( .A(n_285), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_286), .A2(n_454), .B1(n_460), .B2(n_462), .C(n_465), .Y(n_453) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g322 ( .A(n_287), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_287), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g301 ( .A(n_290), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_290), .B(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g356 ( .A(n_291), .Y(n_356) );
NOR2xp33_ASAP7_75t_SL g463 ( .A(n_292), .B(n_317), .Y(n_463) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_293), .B(n_297), .Y(n_330) );
AND2x2_ASAP7_75t_L g361 ( .A(n_293), .B(n_308), .Y(n_361) );
AOI32xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .A3(n_301), .B1(n_303), .B2(n_305), .Y(n_294) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_295), .Y(n_371) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_297), .A2(n_431), .B(n_432), .C(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g436 ( .A(n_297), .Y(n_436) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g314 ( .A(n_299), .Y(n_314) );
OR2x2_ASAP7_75t_L g408 ( .A(n_299), .B(n_304), .Y(n_408) );
AND2x2_ASAP7_75t_L g472 ( .A(n_301), .B(n_314), .Y(n_472) );
INVx1_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
INVx1_ASAP7_75t_L g448 ( .A(n_304), .Y(n_448) );
INVx2_ASAP7_75t_L g459 ( .A(n_304), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_306), .Y(n_397) );
INVx4_ASAP7_75t_L g380 ( .A(n_308), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_324), .C(n_333), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .B(n_318), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_313), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_314), .B(n_323), .Y(n_443) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g319 ( .A(n_316), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_354), .Y(n_353) );
NAND2x1_ASAP7_75t_L g378 ( .A(n_316), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g411 ( .A(n_316), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g469 ( .A(n_316), .B(n_470), .Y(n_469) );
OAI322xp33_ASAP7_75t_L g343 ( .A1(n_317), .A2(n_344), .A3(n_348), .B1(n_350), .B2(n_351), .C1(n_352), .C2(n_355), .Y(n_343) );
INVx1_ASAP7_75t_L g412 ( .A(n_317), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
INVx1_ASAP7_75t_L g468 ( .A(n_320), .Y(n_468) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g363 ( .A(n_322), .Y(n_363) );
OR2x2_ASAP7_75t_L g425 ( .A(n_323), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_326), .B(n_420), .Y(n_480) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g393 ( .A(n_332), .B(n_384), .Y(n_393) );
AND2x2_ASAP7_75t_L g401 ( .A(n_332), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g424 ( .A(n_332), .Y(n_424) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g483 ( .A(n_335), .B(n_385), .Y(n_483) );
INVx1_ASAP7_75t_L g431 ( .A(n_336), .Y(n_431) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx2_ASAP7_75t_L g349 ( .A(n_338), .Y(n_349) );
INVx2_ASAP7_75t_L g406 ( .A(n_339), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_341), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_357), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_346), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g398 ( .A(n_349), .Y(n_398) );
AND2x4_ASAP7_75t_L g405 ( .A(n_349), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g479 ( .A(n_356), .B(n_377), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_362), .B2(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_371), .B(n_372), .C(n_373), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_381), .B2(n_383), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_374), .A2(n_423), .B1(n_425), .B2(n_428), .Y(n_422) );
INVx4_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AND2x4_ASAP7_75t_L g461 ( .A(n_377), .B(n_420), .Y(n_461) );
INVx6_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_380), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI211x1_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_398), .B(n_399), .C(n_409), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2x1_ASAP7_75t_SL g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g407 ( .A(n_393), .Y(n_407) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B1(n_407), .B2(n_408), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g423 ( .A(n_402), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_410), .B(n_430), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_415), .B2(n_419), .C(n_422), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_428), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .C(n_438), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_440), .B(n_453), .Y(n_439) );
OAI21xp33_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_444), .B(n_445), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g464 ( .A(n_450), .Y(n_464) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx4_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_469), .B(n_472), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g486 ( .A(n_480), .Y(n_486) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_675), .B1(n_699), .B2(n_700), .C(n_709), .Y(n_487) );
XNOR2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_652), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
XOR2xp5_ASAP7_75t_L g710 ( .A(n_490), .B(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_543), .C(n_623), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_505), .B(n_535), .Y(n_492) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g508 ( .A(n_495), .Y(n_508) );
AND2x4_ASAP7_75t_L g534 ( .A(n_495), .B(n_524), .Y(n_534) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g641 ( .A(n_496), .B(n_538), .Y(n_641) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g504 ( .A(n_497), .Y(n_504) );
AND2x4_ASAP7_75t_L g651 ( .A(n_497), .B(n_538), .Y(n_651) );
OR2x2_ASAP7_75t_L g688 ( .A(n_497), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g698 ( .A(n_497), .B(n_689), .Y(n_698) );
OR2x2_ASAP7_75t_L g502 ( .A(n_498), .B(n_503), .Y(n_502) );
INVx8_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AND2x4_ASAP7_75t_L g518 ( .A(n_500), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g528 ( .A(n_501), .Y(n_528) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g527 ( .A(n_504), .B(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g530 ( .A(n_504), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x6_ASAP7_75t_L g515 ( .A(n_508), .B(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g628 ( .A(n_510), .Y(n_628) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
AND2x4_ASAP7_75t_L g525 ( .A(n_511), .B(n_519), .Y(n_525) );
INVx1_ASAP7_75t_L g532 ( .A(n_511), .Y(n_532) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g635 ( .A(n_512), .B(n_513), .Y(n_635) );
INVx2_ASAP7_75t_L g519 ( .A(n_513), .Y(n_519) );
CKINVDCx14_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx12f_ASAP7_75t_L g631 ( .A(n_518), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_534), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_524), .Y(n_638) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .B1(n_530), .B2(n_533), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_528), .B(n_685), .C(n_687), .Y(n_684) );
AND2x4_ASAP7_75t_L g695 ( .A(n_528), .B(n_696), .Y(n_695) );
AOI222xp33_ASAP7_75t_L g568 ( .A1(n_529), .A2(n_569), .B1(n_570), .B2(n_574), .C1(n_576), .C2(n_577), .Y(n_568) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_540), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g689 ( .A(n_539), .Y(n_689) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g586 ( .A(n_541), .Y(n_586) );
INVx1_ASAP7_75t_L g606 ( .A(n_541), .Y(n_606) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND3x1_ASAP7_75t_L g620 ( .A(n_542), .B(n_621), .C(n_622), .Y(n_620) );
INVx2_ASAP7_75t_L g640 ( .A(n_542), .Y(n_640) );
INVx1_ASAP7_75t_L g650 ( .A(n_542), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_566), .B(n_582), .C(n_587), .Y(n_543) );
OR2x2_ASAP7_75t_SL g545 ( .A(n_546), .B(n_550), .Y(n_545) );
OR2x6_ASAP7_75t_L g567 ( .A(n_546), .B(n_554), .Y(n_567) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x4_ASAP7_75t_L g564 ( .A(n_548), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g573 ( .A(n_548), .Y(n_573) );
INVx2_ASAP7_75t_L g565 ( .A(n_549), .Y(n_565) );
INVx2_ASAP7_75t_L g572 ( .A(n_549), .Y(n_572) );
INVx3_ASAP7_75t_R g561 ( .A(n_550), .Y(n_561) );
AND2x4_ASAP7_75t_L g581 ( .A(n_550), .B(n_571), .Y(n_581) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g574 ( .A(n_555), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_SL g577 ( .A(n_555), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g621 ( .A(n_555), .Y(n_621) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx12f_ASAP7_75t_SL g598 ( .A(n_557), .Y(n_598) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_558), .Y(n_616) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx4_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_564), .Y(n_602) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_565), .Y(n_575) );
INVx1_ASAP7_75t_L g593 ( .A(n_565), .Y(n_593) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx2_ASAP7_75t_L g594 ( .A(n_571), .Y(n_594) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g592 ( .A(n_579), .B(n_593), .Y(n_592) );
CKINVDCx8_ASAP7_75t_R g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_610), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_595), .C(n_603), .Y(n_588) );
INVx4_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
INVx5_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .C(n_617), .Y(n_610) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_642), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_632), .C(n_639), .Y(n_624) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g645 ( .A(n_631), .Y(n_645) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g648 ( .A(n_634), .Y(n_648) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x6_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .C(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x6_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
XOR2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_666), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_664), .B2(n_665), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_655) );
INVx1_ASAP7_75t_L g662 ( .A(n_656), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_659), .Y(n_660) );
INVx2_ASAP7_75t_L g663 ( .A(n_661), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_664), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_673), .B2(n_674), .Y(n_666) );
INVx1_ASAP7_75t_L g673 ( .A(n_667), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_668), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_669), .Y(n_672) );
INVx1_ASAP7_75t_L g671 ( .A(n_670), .Y(n_671) );
BUFx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x6_ASAP7_75t_L g677 ( .A(n_678), .B(n_690), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_683), .Y(n_678) );
INVxp67_ASAP7_75t_L g716 ( .A(n_679), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g708 ( .A(n_680), .Y(n_708) );
INVx1_ASAP7_75t_L g720 ( .A(n_681), .Y(n_720) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g707 ( .A(n_682), .Y(n_707) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_684), .B(n_694), .Y(n_717) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
CKINVDCx11_ASAP7_75t_R g692 ( .A(n_686), .Y(n_692) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
INVx3_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_704), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g719 ( .A(n_708), .B(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B1(n_718), .B2(n_721), .Y(n_709) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx4f_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx4_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
endmodule