module real_jpeg_4152_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_0),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_0),
.B(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_0),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_0),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_0),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_0),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_0),
.B(n_108),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_1),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_1),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_1),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_1),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_2),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_2),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_2),
.B(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_4),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_4),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_4),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_4),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_5),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_5),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_5),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_5),
.B(n_203),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_5),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_5),
.B(n_196),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_8),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_8),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_8),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_8),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_8),
.B(n_356),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_8),
.B(n_99),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_8),
.B(n_295),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_9),
.Y(n_531)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_10),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_10),
.Y(n_373)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_12),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_14),
.B(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_14),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_14),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_14),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_14),
.B(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_14),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_15),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_15),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_15),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_15),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_15),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_15),
.B(n_183),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_15),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_15),
.B(n_359),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_16),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_16),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_16),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_16),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_16),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_16),
.B(n_391),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_16),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_17),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_17),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_17),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_17),
.B(n_99),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_17),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_17),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_17),
.B(n_313),
.Y(n_417)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_19),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_19),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_19),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_19),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_19),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_529),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_22),
.Y(n_530)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_43),
.B(n_78),
.C(n_528),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_51),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_27),
.B(n_51),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.C(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_29),
.A2(n_33),
.B1(n_42),
.B2(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_31),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_55),
.C(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_35),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_40),
.Y(n_152)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_74),
.C(n_76),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_63),
.C(n_64),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_60),
.B1(n_70),
.B2(n_111),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_57),
.Y(n_278)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_58),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.C(n_70),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_64),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_66),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_68),
.Y(n_286)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_70),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_72),
.Y(n_208)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_72),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_72),
.Y(n_412)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_122),
.B(n_527),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_119),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_80),
.B(n_119),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_116),
.C(n_117),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_81),
.A2(n_82),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_104),
.C(n_112),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_83),
.A2(n_84),
.B1(n_504),
.B2(n_506),
.Y(n_503)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_90),
.C(n_93),
.Y(n_116)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_92),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_100),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_94),
.B(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_494)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_104),
.A2(n_112),
.B1(n_113),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_104),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.C(n_111),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_105),
.B(n_500),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_106),
.A2(n_107),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_107),
.B(n_191),
.C(n_195),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_116),
.B(n_117),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_521),
.B(n_526),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_487),
.B(n_518),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_298),
.B(n_486),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_248),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_126),
.B(n_248),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_188),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_127),
.B(n_189),
.C(n_225),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_162),
.C(n_171),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_128),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_149),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_129),
.B(n_471),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_133),
.C(n_136),
.Y(n_170)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_131),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_147),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_141),
.B(n_147),
.Y(n_461)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_144),
.B(n_461),
.Y(n_460)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_149),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_150),
.B(n_154),
.C(n_159),
.Y(n_245)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_157),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_157),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_158),
.B(n_195),
.C(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_158),
.A2(n_159),
.B1(n_195),
.B2(n_198),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_171),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_170),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_168),
.C(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_166),
.A2(n_169),
.B1(n_237),
.B2(n_241),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_169),
.B(n_230),
.C(n_241),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_182),
.C(n_184),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_172),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_180),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_173),
.B(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_177),
.B(n_180),
.Y(n_260)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_182),
.B(n_184),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_225),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_199),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_190),
.B(n_200),
.C(n_209),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_195),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_209),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.C(n_206),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_206),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_204),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g356 ( 
.A(n_208),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_222),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_211),
.B(n_217),
.C(n_222),
.Y(n_502)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_216),
.Y(n_360)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_242),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_227),
.B(n_229),
.C(n_242),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.C(n_246),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_255),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_250),
.B(n_253),
.Y(n_481)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_255),
.B(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_279),
.C(n_282),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_257),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.C(n_267),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_258),
.A2(n_259),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_261),
.A2(n_262),
.B(n_265),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_261),
.B(n_267),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.C(n_276),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_429)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_276),
.B(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_277),
.B(n_372),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_282),
.Y(n_475)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_291),
.C(n_294),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_284),
.B(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_285),
.B(n_441),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_287),
.Y(n_442)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_291),
.B(n_294),
.Y(n_463)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_479),
.B(n_485),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_466),
.B(n_478),
.Y(n_299)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_448),
.B(n_465),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_422),
.B(n_447),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_396),
.B(n_421),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_364),
.B(n_395),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_345),
.B(n_363),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_326),
.B(n_344),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_320),
.B(n_325),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_316),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_316),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_312),
.Y(n_327)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_328),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_336),
.B2(n_337),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_339),
.C(n_341),
.Y(n_362)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_334),
.Y(n_353)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_362),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_362),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_353),
.C(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_351),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_384),
.C(n_385),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_367),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_382),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_383),
.C(n_386),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_371),
.C(n_374),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

INVx4_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_377),
.B1(n_378),
.B2(n_381),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_375),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_381),
.Y(n_405)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_392),
.C(n_393),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_390),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_392),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_420),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_420),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_407),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_406),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_406),
.C(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_405),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_436),
.C(n_437),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_413),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_415),
.C(n_418),
.Y(n_425)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_408),
.Y(n_532)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_410),
.CI(n_411),
.CON(n_408),
.SN(n_408)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_410),
.C(n_411),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_418),
.B2(n_419),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_417),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_445),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_445),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_434),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_426),
.C(n_434),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_457),
.C(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_438),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_439),
.C(n_444),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_443),
.B2(n_444),
.Y(n_438)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_439),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_464),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_464),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_455),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_454),
.C(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_452),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_455),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_460),
.C(n_462),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_476),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_476),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_483),
.C(n_484),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_482),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_480),
.B(n_482),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_515),
.Y(n_487)
);

OAI21xp33_ASAP7_75t_L g518 ( 
.A1(n_488),
.A2(n_519),
.B(n_520),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_508),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_508),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_491),
.B1(n_497),
.B2(n_507),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_490),
.B(n_498),
.C(n_503),
.Y(n_525)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.C(n_495),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_510),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_493),
.A2(n_495),
.B1(n_496),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_503),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.C(n_502),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_513),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_502),
.Y(n_513)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_504),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_512),
.C(n_514),
.Y(n_508)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_509),
.B(n_512),
.CI(n_514),
.CON(n_516),
.SN(n_516)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_517),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_516),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_525),
.Y(n_526)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_523),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);


endmodule