module fake_jpeg_29176_n_483 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_483);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_483;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_50),
.B(n_54),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_86),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_22),
.C(n_35),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_81),
.C(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_68),
.Y(n_149)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_8),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_10),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_79),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_76),
.B(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_24),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_10),
.B(n_14),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_10),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_87),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_29),
.B1(n_23),
.B2(n_41),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_101),
.A2(n_129),
.B1(n_11),
.B2(n_15),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_104),
.A2(n_106),
.B1(n_113),
.B2(n_118),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_77),
.B1(n_84),
.B2(n_85),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_37),
.B1(n_26),
.B2(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_81),
.B(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_133),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_67),
.A2(n_37),
.B1(n_26),
.B2(n_43),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_36),
.Y(n_119)
);

OR2x4_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_73),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_74),
.A2(n_24),
.B1(n_41),
.B2(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_121),
.A2(n_134),
.B1(n_151),
.B2(n_96),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_30),
.B1(n_34),
.B2(n_31),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_47),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_83),
.A2(n_44),
.B1(n_42),
.B2(n_45),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_88),
.B(n_47),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_42),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_34),
.B1(n_31),
.B2(n_44),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_62),
.B(n_40),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_153),
.B(n_159),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_148),
.C(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_100),
.B(n_82),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_155),
.B(n_170),
.Y(n_234)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_156),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_99),
.A2(n_123),
.A3(n_124),
.B1(n_102),
.B2(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_160),
.B(n_162),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_78),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_164),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_90),
.B1(n_80),
.B2(n_95),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_166),
.A2(n_198),
.B1(n_201),
.B2(n_110),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_78),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_169),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_102),
.B(n_12),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_44),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_176),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_36),
.B(n_33),
.C(n_32),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_178),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_181),
.C(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_103),
.B(n_45),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_45),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_180),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_36),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_45),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_120),
.B(n_65),
.Y(n_181)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_143),
.B1(n_131),
.B2(n_130),
.Y(n_237)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_45),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_192),
.Y(n_226)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_125),
.A2(n_57),
.B(n_92),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_112),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_94),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx9p33_ASAP7_75t_R g191 ( 
.A(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_109),
.B(n_11),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_146),
.B(n_11),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_14),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_195),
.A2(n_104),
.B1(n_113),
.B2(n_118),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_130),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_137),
.A2(n_33),
.B1(n_32),
.B2(n_2),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_135),
.B(n_143),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_132),
.A2(n_33),
.B1(n_6),
.B2(n_2),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_144),
.B1(n_122),
.B2(n_108),
.Y(n_224)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_203),
.B(n_233),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_154),
.B(n_172),
.C(n_191),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_147),
.B1(n_140),
.B2(n_110),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_238),
.B(n_199),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_211),
.A2(n_213),
.B1(n_222),
.B2(n_240),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_157),
.B1(n_160),
.B2(n_178),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_155),
.A2(n_147),
.B1(n_140),
.B2(n_108),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_221),
.B1(n_235),
.B2(n_238),
.Y(n_246)
);

AOI22x1_ASAP7_75t_SL g235 ( 
.A1(n_164),
.A2(n_144),
.B1(n_122),
.B2(n_135),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_179),
.B(n_187),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_241),
.B1(n_168),
.B2(n_198),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_163),
.A2(n_171),
.B1(n_182),
.B2(n_161),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_182),
.A2(n_131),
.B1(n_6),
.B2(n_4),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_153),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_243),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_186),
.B1(n_176),
.B2(n_177),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_252),
.B1(n_277),
.B2(n_224),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_246),
.A2(n_229),
.B1(n_230),
.B2(n_216),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_247),
.A2(n_248),
.B(n_253),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_158),
.B1(n_185),
.B2(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_251),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_159),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_170),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_256),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_212),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_209),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_234),
.B(n_158),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_274),
.C(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_263),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_189),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_202),
.B(n_201),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_200),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_158),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_221),
.A2(n_198),
.B1(n_197),
.B2(n_168),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_231),
.B1(n_232),
.B2(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_206),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_226),
.B(n_174),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_209),
.A2(n_174),
.B(n_169),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_204),
.B(n_229),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_210),
.A2(n_197),
.B1(n_165),
.B2(n_156),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_280),
.A2(n_300),
.B(n_302),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_281),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_254),
.B(n_203),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_270),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_304),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_247),
.A2(n_213),
.B1(n_204),
.B2(n_211),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_207),
.B1(n_218),
.B2(n_230),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_229),
.C(n_218),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_303),
.C(n_305),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_246),
.A2(n_231),
.B1(n_228),
.B2(n_232),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_236),
.B(n_228),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_214),
.B(n_219),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_264),
.A2(n_219),
.B1(n_215),
.B2(n_214),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_233),
.B(n_215),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_219),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_183),
.B1(n_173),
.B2(n_0),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_4),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_274),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_313),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_245),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_316),
.C(n_325),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_328),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_242),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_319),
.B(n_330),
.Y(n_367)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_255),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_279),
.B(n_251),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_279),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_329),
.B(n_335),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_262),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_333),
.B(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_337),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_288),
.B(n_272),
.Y(n_335)
);

NOR2x1_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_272),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_267),
.C(n_273),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_345),
.C(n_299),
.Y(n_362)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_341),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_269),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_257),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_343),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_291),
.B(n_258),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_344),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_280),
.B(n_249),
.C(n_244),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_289),
.B1(n_290),
.B2(n_292),
.Y(n_346)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_268),
.B1(n_248),
.B2(n_313),
.Y(n_351)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_337),
.B1(n_297),
.B2(n_336),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_354),
.A2(n_358),
.B1(n_371),
.B2(n_372),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_320),
.A2(n_337),
.B1(n_336),
.B2(n_326),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_322),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_341),
.Y(n_382)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_302),
.C(n_283),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_360),
.B(n_332),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_338),
.C(n_324),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_318),
.A2(n_312),
.B1(n_304),
.B2(n_253),
.Y(n_364)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_340),
.A2(n_301),
.B1(n_300),
.B2(n_277),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_312),
.B1(n_296),
.B2(n_253),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_305),
.Y(n_373)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_318),
.A2(n_271),
.B1(n_285),
.B2(n_283),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_271),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_324),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_376),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_352),
.B(n_316),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_356),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_377),
.B(n_353),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g401 ( 
.A1(n_381),
.A2(n_367),
.B(n_349),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_382),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_389),
.C(n_391),
.Y(n_400)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g387 ( 
.A(n_347),
.B(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_387),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_397),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_345),
.C(n_315),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_325),
.C(n_314),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_314),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_399),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_361),
.A2(n_317),
.B(n_334),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_393),
.A2(n_398),
.B(n_355),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_331),
.C(n_327),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_355),
.C(n_357),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_285),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_401),
.B(n_402),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_383),
.B(n_385),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_404),
.A2(n_393),
.B(n_392),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_378),
.A2(n_369),
.B1(n_349),
.B2(n_359),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

BUFx12_ASAP7_75t_L g410 ( 
.A(n_387),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_387),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_412),
.C(n_413),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_372),
.C(n_357),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_353),
.C(n_364),
.Y(n_413)
);

A2O1A1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_361),
.B(n_368),
.C(n_363),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_374),
.B1(n_371),
.B2(n_363),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_416),
.A2(n_419),
.B1(n_382),
.B2(n_397),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_399),
.A2(n_370),
.B1(n_368),
.B2(n_339),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_420),
.B(n_426),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_391),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_403),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_425),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_394),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_411),
.B(n_395),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_435),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_419),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_406),
.A2(n_386),
.B1(n_408),
.B2(n_380),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_430),
.A2(n_406),
.B1(n_414),
.B2(n_410),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_396),
.B1(n_388),
.B2(n_370),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_433),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_415),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_423),
.B(n_400),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_438),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_309),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_423),
.B(n_400),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_440),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_421),
.A2(n_389),
.B(n_410),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_443),
.B(n_444),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_432),
.A2(n_417),
.B(n_416),
.C(n_409),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_432),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_311),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_403),
.C(n_409),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_448),
.C(n_422),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_376),
.C(n_298),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_441),
.A2(n_421),
.B(n_429),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_450),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_449),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_431),
.C(n_426),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_456),
.Y(n_469)
);

AOI21x1_ASAP7_75t_SL g454 ( 
.A1(n_437),
.A2(n_428),
.B(n_420),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_454),
.A2(n_263),
.B(n_275),
.C(n_278),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_445),
.A2(n_298),
.B(n_309),
.Y(n_455)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_455),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_SL g457 ( 
.A(n_448),
.B(n_311),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_275),
.B(n_5),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_460),
.B(n_461),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_442),
.Y(n_461)
);

NOR2x1_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_444),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_465),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_452),
.A2(n_439),
.B(n_260),
.Y(n_467)
);

AO21x1_ASAP7_75t_L g473 ( 
.A1(n_467),
.A2(n_468),
.B(n_470),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_451),
.C(n_453),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_472),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_469),
.B(n_458),
.Y(n_474)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_474),
.A2(n_475),
.B(n_462),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_459),
.Y(n_475)
);

AOI21xp33_ASAP7_75t_L g480 ( 
.A1(n_477),
.A2(n_478),
.B(n_5),
.Y(n_480)
);

AOI321xp33_ASAP7_75t_SL g478 ( 
.A1(n_471),
.A2(n_466),
.A3(n_455),
.B1(n_468),
.B2(n_13),
.C(n_15),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_466),
.C(n_473),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_479),
.A2(n_480),
.B(n_12),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

O2A1O1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_0),
.B(n_15),
.C(n_464),
.Y(n_483)
);


endmodule