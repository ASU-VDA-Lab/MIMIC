module fake_jpeg_22567_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_8),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_24),
.B1(n_31),
.B2(n_26),
.Y(n_70)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_45),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_21),
.B1(n_25),
.B2(n_22),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_45),
.B(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_69),
.B1(n_24),
.B2(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_49),
.C(n_20),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_37),
.B1(n_25),
.B2(n_31),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_102),
.B1(n_30),
.B2(n_32),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_39),
.C(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_40),
.C(n_46),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_83),
.B1(n_100),
.B2(n_28),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_51),
.B1(n_47),
.B2(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_41),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_85),
.Y(n_135)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_90),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_51),
.B1(n_42),
.B2(n_37),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_30),
.B1(n_20),
.B2(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_18),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_38),
.B(n_39),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_97),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_103),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_39),
.B1(n_38),
.B2(n_59),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_119),
.B1(n_126),
.B2(n_127),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_39),
.B1(n_59),
.B2(n_50),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_99),
.B1(n_84),
.B2(n_92),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_100),
.C(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_80),
.B1(n_83),
.B2(n_74),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_54),
.B1(n_60),
.B2(n_68),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_80),
.A2(n_63),
.B1(n_67),
.B2(n_19),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_19),
.B1(n_23),
.B2(n_27),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_146),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_160),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_144),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_78),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_149),
.C(n_160),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_97),
.CI(n_92),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_73),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_157),
.B1(n_165),
.B2(n_121),
.Y(n_196)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_150),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_108),
.B(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_46),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_164),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_0),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_129),
.B(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_156),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_103),
.B1(n_105),
.B2(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_130),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_40),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_91),
.C(n_40),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_136),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_116),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_19),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_117),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_46),
.C(n_36),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_95),
.B1(n_91),
.B2(n_71),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVxp67_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_200),
.B(n_144),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_170),
.B(n_187),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_35),
.B(n_12),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_110),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_176),
.B(n_132),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_118),
.B1(n_113),
.B2(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_143),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_33),
.C(n_2),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_123),
.B1(n_133),
.B2(n_124),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_195),
.B1(n_196),
.B2(n_156),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_117),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_198),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_138),
.A2(n_112),
.B1(n_113),
.B2(n_118),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_145),
.B1(n_164),
.B2(n_138),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_36),
.B1(n_71),
.B2(n_19),
.Y(n_215)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_9),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_112),
.B(n_32),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_202),
.B(n_227),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_210),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_142),
.B(n_152),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_173),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_214),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_135),
.A3(n_72),
.B1(n_79),
.B2(n_81),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_132),
.B1(n_71),
.B2(n_34),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_36),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_171),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_29),
.B1(n_27),
.B2(n_23),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_29),
.B1(n_27),
.B2(n_23),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_29),
.B1(n_23),
.B2(n_35),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_229),
.B1(n_192),
.B2(n_199),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_225),
.C(n_226),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_33),
.A3(n_8),
.B1(n_9),
.B2(n_16),
.C1(n_15),
.C2(n_14),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_184),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_33),
.C(n_2),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_33),
.C(n_2),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_16),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_1),
.C(n_2),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_179),
.C(n_178),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_177),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_252),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_243),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_206),
.B1(n_195),
.B2(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_169),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_181),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_213),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_167),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_256),
.C(n_257),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_205),
.B(n_174),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_185),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_174),
.C(n_186),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_186),
.C(n_188),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_270),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_212),
.B1(n_203),
.B2(n_215),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_233),
.B1(n_234),
.B2(n_239),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_223),
.C(n_214),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_228),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_204),
.C(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_247),
.B1(n_235),
.B2(n_218),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_230),
.B(n_188),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_220),
.B(n_230),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_205),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_279),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_238),
.B1(n_236),
.B2(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_295),
.B1(n_270),
.B2(n_265),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_268),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_249),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_296),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_297),
.B(n_279),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_277),
.B(n_253),
.Y(n_291)
);

OAI221xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_293),
.B1(n_264),
.B2(n_278),
.C(n_258),
.Y(n_302)
);

OA21x2_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_245),
.B(n_251),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_234),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_265),
.C(n_258),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_304),
.C(n_306),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_303),
.B(n_5),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_286),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_300),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_302),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_269),
.C(n_239),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_273),
.C(n_243),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_9),
.B1(n_16),
.B2(n_14),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_216),
.C(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.C(n_284),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_1),
.C(n_4),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_294),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_298),
.B(n_311),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_323),
.B(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_319),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_296),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_322),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_10),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_325),
.B(n_328),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_309),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_309),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_317),
.B(n_10),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_324),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_335),
.B(n_339),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_327),
.A2(n_316),
.B(n_11),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_337),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_326),
.A2(n_316),
.B1(n_11),
.B2(n_14),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_6),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_6),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_329),
.C(n_6),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_341),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

AO21x2_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_343),
.B(n_342),
.Y(n_346)
);

AOI31xp33_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_338),
.A3(n_344),
.B(n_334),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_6),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_348),
.A2(n_7),
.B(n_172),
.Y(n_349)
);


endmodule