module fake_netlist_6_4246_n_1021 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1021);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1021;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_575;
wire n_368;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_643;
wire n_349;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_608;
wire n_261;
wire n_474;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_273;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_550;
wire n_487;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_672;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_515;
wire n_315;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_385;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_663;
wire n_361;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_82),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_157),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_149),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_108),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_146),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_122),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_59),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_5),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_142),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_88),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_20),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_114),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_86),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_119),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_75),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_92),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_90),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_94),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_121),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_91),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_41),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_197),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_155),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_70),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_83),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_117),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_39),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_21),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_178),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_65),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_72),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_20),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_125),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_30),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_29),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_200),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_128),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_154),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_67),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_143),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_179),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_89),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_141),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_100),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_172),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_93),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_165),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_24),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_147),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_81),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_223),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_139),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_156),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_145),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_104),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_152),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_189),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_102),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_133),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_182),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_151),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_38),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_217),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_214),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_161),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_57),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_60),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_130),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_137),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_221),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_18),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_211),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_44),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_53),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_77),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_69),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_129),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_47),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_203),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_168),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_76),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_80),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_124),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_135),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_73),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_113),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_170),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_103),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_66),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_195),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_111),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_207),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_169),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_191),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_31),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_175),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_63),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_224),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_11),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_118),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_192),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_29),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_213),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_19),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_212),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_49),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_115),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_159),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_4),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_140),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_183),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_148),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_225),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_131),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_54),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_204),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_40),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_144),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_173),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_171),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_181),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_180),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_0),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_55),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_43),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_64),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_79),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_127),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_153),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_134),
.Y(n_383)
);

BUFx8_ASAP7_75t_SL g384 ( 
.A(n_107),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_193),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_187),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_84),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_48),
.B(n_97),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_61),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_245),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_250),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_252),
.B(n_0),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_271),
.B(n_1),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_290),
.B(n_1),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_250),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_250),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_262),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_5),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_279),
.Y(n_399)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_245),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_305),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_291),
.B(n_6),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_321),
.B(n_287),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_7),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_276),
.B(n_8),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_259),
.A2(n_278),
.B(n_263),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_245),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_303),
.A2(n_45),
.B(n_42),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_245),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_262),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_266),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_239),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_286),
.B(n_9),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_9),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_235),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_262),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_242),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_272),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_244),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_384),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_294),
.B(n_319),
.Y(n_421)
);

AOI22x1_ASAP7_75t_SL g422 ( 
.A1(n_229),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_319),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_262),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_304),
.A2(n_50),
.B(n_46),
.Y(n_425)
);

OAI22x1_ASAP7_75t_SL g426 ( 
.A1(n_247),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_262),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_345),
.B(n_13),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_266),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_347),
.B(n_15),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g431 ( 
.A(n_277),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_230),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_306),
.B(n_17),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_306),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_262),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_306),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_306),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_231),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_369),
.B(n_18),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_280),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_372),
.B(n_19),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_227),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_316),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_316),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_282),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_316),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_316),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_228),
.A2(n_52),
.B(n_51),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_236),
.B(n_21),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_232),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_241),
.A2(n_22),
.B(n_23),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_233),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_243),
.B(n_23),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_296),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_298),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_378),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_353),
.B(n_25),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_254),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_56),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_378),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_256),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_258),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_234),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_310),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_237),
.Y(n_469)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_346),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_267),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_226),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_322),
.B(n_32),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_268),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_270),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_360),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_275),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_283),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_285),
.Y(n_479)
);

AOI22x1_ASAP7_75t_SL g480 ( 
.A1(n_350),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_238),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_288),
.A2(n_160),
.B(n_220),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_297),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_240),
.Y(n_484)
);

BUFx8_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_302),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_323),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_376),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_324),
.A2(n_163),
.B(n_219),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_327),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_246),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_333),
.A2(n_36),
.B(n_37),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_334),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_335),
.B(n_37),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_341),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_260),
.B(n_38),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_281),
.B(n_62),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_248),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_348),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_362),
.B(n_71),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_249),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_251),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_253),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_255),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_373),
.B(n_74),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_438),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_472),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_488),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_454),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_443),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_469),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_491),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_501),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_502),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_395),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_396),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_432),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_452),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_484),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_431),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_445),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_R g528 ( 
.A(n_440),
.B(n_292),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_498),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_403),
.B(n_320),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_R g532 ( 
.A(n_456),
.B(n_357),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_485),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_503),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_503),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_444),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_504),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_485),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_444),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_448),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_504),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_467),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_481),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_R g548 ( 
.A(n_457),
.B(n_365),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_415),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_449),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_415),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_417),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_419),
.Y(n_554)
);

AND3x2_ASAP7_75t_L g555 ( 
.A(n_430),
.B(n_377),
.C(n_375),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_470),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_470),
.B(n_382),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_399),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_476),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_459),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_476),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_401),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_497),
.B(n_371),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_496),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_493),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_471),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_R g570 ( 
.A(n_442),
.B(n_257),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_471),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_398),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_397),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_418),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_483),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_573),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_523),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_564),
.B(n_394),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_531),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_574),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_553),
.B(n_505),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_544),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_542),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_512),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_567),
.B(n_461),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_528),
.A2(n_500),
.B(n_482),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_512),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_520),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_509),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_553),
.B(n_390),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_563),
.B(n_405),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_533),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_514),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_530),
.B(n_390),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_536),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_571),
.B(n_428),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_524),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_506),
.B(n_390),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_400),
.Y(n_599)
);

BUFx6f_ASAP7_75t_SL g600 ( 
.A(n_510),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_546),
.B(n_400),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_532),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_547),
.B(n_400),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_560),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_511),
.B(n_413),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_560),
.B(n_411),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_562),
.B(n_411),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_562),
.B(n_411),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_513),
.B(n_367),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_543),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_568),
.B(n_434),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_575),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_555),
.B(n_392),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_518),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_548),
.B(n_528),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_508),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_548),
.B(n_392),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_572),
.A2(n_473),
.B1(n_468),
.B2(n_433),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_517),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_558),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_515),
.B(n_393),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_551),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_529),
.B(n_434),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_535),
.B(n_437),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_538),
.B(n_437),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_570),
.B(n_463),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_517),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_540),
.B(n_447),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_554),
.B(n_466),
.C(n_465),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_521),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_545),
.B(n_458),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_522),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_557),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_570),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_525),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_576),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_584),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_604),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_581),
.B(n_451),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_608),
.B(n_451),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_SL g646 ( 
.A(n_622),
.B(n_527),
.C(n_526),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_612),
.B(n_639),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_616),
.B(n_402),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_635),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_583),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_591),
.B(n_455),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_604),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_593),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_635),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_587),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_602),
.B(n_556),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_594),
.B(n_494),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_621),
.B(n_566),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_598),
.B(n_404),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_623),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_595),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_635),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_637),
.B(n_404),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_625),
.B(n_559),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_615),
.B(n_601),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_578),
.B(n_552),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_637),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_607),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_637),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_582),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_606),
.B(n_414),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_624),
.B(n_414),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_632),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_618),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_632),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_624),
.B(n_561),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_577),
.Y(n_679)
);

XOR2xp5_ASAP7_75t_L g680 ( 
.A(n_589),
.B(n_565),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_624),
.B(n_439),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_632),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_579),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_619),
.B(n_510),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_640),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_596),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_585),
.B(n_441),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_617),
.B(n_516),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_590),
.B(n_441),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_588),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_617),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_597),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_626),
.B(n_534),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_631),
.A2(n_264),
.B1(n_265),
.B2(n_261),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_627),
.B(n_479),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_600),
.B(n_541),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_603),
.B(n_269),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_605),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_620),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_610),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_599),
.B(n_463),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_586),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_611),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_634),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_628),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_645),
.B(n_629),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_663),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_670),
.B(n_453),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_L g713 ( 
.A1(n_672),
.A2(n_495),
.B(n_499),
.C(n_487),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_651),
.A2(n_492),
.B1(n_273),
.B2(n_274),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_674),
.A2(n_489),
.B(n_450),
.Y(n_715)
);

AO32x2_ASAP7_75t_L g716 ( 
.A1(n_686),
.A2(n_422),
.A3(n_480),
.B1(n_426),
.B2(n_406),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_644),
.B(n_630),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_657),
.B(n_633),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_687),
.A2(n_425),
.B(n_408),
.C(n_462),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_702),
.A2(n_475),
.B(n_486),
.C(n_462),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_654),
.B(n_636),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_685),
.B(n_284),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_669),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_412),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_668),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_649),
.B(n_670),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_647),
.B(n_289),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_641),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_684),
.B(n_293),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_641),
.B(n_295),
.Y(n_730)
);

AOI21xp33_ASAP7_75t_L g731 ( 
.A1(n_667),
.A2(n_300),
.B(n_299),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_689),
.B(n_301),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_702),
.A2(n_486),
.B(n_475),
.C(n_424),
.Y(n_733)
);

INVx5_ASAP7_75t_L g734 ( 
.A(n_664),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_671),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_681),
.A2(n_458),
.B(n_416),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_695),
.B(n_307),
.Y(n_737)
);

AOI21x1_ASAP7_75t_L g738 ( 
.A1(n_705),
.A2(n_427),
.B(n_410),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_662),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_SL g740 ( 
.A1(n_707),
.A2(n_435),
.B(n_389),
.C(n_387),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_658),
.B(n_309),
.C(n_308),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_691),
.Y(n_742)
);

INVx6_ASAP7_75t_L g743 ( 
.A(n_653),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_655),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_666),
.A2(n_351),
.B1(n_312),
.B2(n_313),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_642),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_692),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_677),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_704),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_706),
.A2(n_708),
.B1(n_664),
.B2(n_659),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_703),
.B(n_311),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_701),
.B(n_474),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_655),
.Y(n_753)
);

NOR3xp33_ASAP7_75t_L g754 ( 
.A(n_693),
.B(n_315),
.C(n_314),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_648),
.A2(n_356),
.B(n_325),
.C(n_326),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_675),
.B(n_478),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_678),
.A2(n_328),
.B(n_318),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_706),
.A2(n_330),
.B(n_329),
.Y(n_758)
);

OAI22x1_ASAP7_75t_L g759 ( 
.A1(n_680),
.A2(n_386),
.B1(n_385),
.B2(n_383),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_643),
.A2(n_336),
.B(n_332),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_709),
.B(n_337),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_652),
.A2(n_339),
.B(n_338),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_709),
.B(n_661),
.Y(n_763)
);

INVx5_ASAP7_75t_SL g764 ( 
.A(n_748),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_739),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_749),
.Y(n_766)
);

BUFx5_ASAP7_75t_L g767 ( 
.A(n_728),
.Y(n_767)
);

AOI21x1_ASAP7_75t_L g768 ( 
.A1(n_715),
.A2(n_673),
.B(n_676),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_746),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_725),
.Y(n_770)
);

BUFx8_ASAP7_75t_L g771 ( 
.A(n_716),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_711),
.Y(n_772)
);

OA21x2_ASAP7_75t_L g773 ( 
.A1(n_719),
.A2(n_736),
.B(n_713),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_724),
.Y(n_774)
);

AOI22x1_ASAP7_75t_L g775 ( 
.A1(n_712),
.A2(n_699),
.B1(n_700),
.B2(n_679),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_738),
.A2(n_683),
.B(n_694),
.Y(n_776)
);

BUFx8_ASAP7_75t_L g777 ( 
.A(n_716),
.Y(n_777)
);

AO21x2_ASAP7_75t_L g778 ( 
.A1(n_750),
.A2(n_665),
.B(n_646),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_734),
.B(n_690),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_735),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_734),
.B(n_698),
.Y(n_781)
);

OAI21x1_ASAP7_75t_L g782 ( 
.A1(n_763),
.A2(n_656),
.B(n_697),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_744),
.A2(n_688),
.B(n_704),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_743),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_744),
.A2(n_682),
.B(n_660),
.Y(n_786)
);

AO21x2_ASAP7_75t_L g787 ( 
.A1(n_710),
.A2(n_342),
.B(n_340),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_743),
.B(n_696),
.Y(n_788)
);

BUFx2_ASAP7_75t_SL g789 ( 
.A(n_726),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_752),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_749),
.Y(n_791)
);

INVx6_ASAP7_75t_L g792 ( 
.A(n_748),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_742),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_753),
.A2(n_85),
.B(n_87),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_733),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_722),
.B(n_490),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_717),
.A2(n_381),
.B(n_380),
.Y(n_798)
);

INVx8_ASAP7_75t_L g799 ( 
.A(n_721),
.Y(n_799)
);

AOI21xp33_ASAP7_75t_L g800 ( 
.A1(n_729),
.A2(n_366),
.B(n_344),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_748),
.Y(n_801)
);

INVxp33_ASAP7_75t_L g802 ( 
.A(n_759),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_718),
.B(n_343),
.Y(n_803)
);

AO21x2_ASAP7_75t_L g804 ( 
.A1(n_714),
.A2(n_379),
.B(n_374),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_730),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_721),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_720),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_756),
.Y(n_808)
);

AO21x2_ASAP7_75t_L g809 ( 
.A1(n_732),
.A2(n_370),
.B(n_368),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_751),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_761),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_740),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_785),
.Y(n_813)
);

NAND2x1p5_ASAP7_75t_L g814 ( 
.A(n_791),
.B(n_727),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_784),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_771),
.A2(n_731),
.B1(n_754),
.B2(n_741),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_767),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_793),
.Y(n_818)
);

BUFx4f_ASAP7_75t_SL g819 ( 
.A(n_801),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_766),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_766),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_769),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_766),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_780),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_767),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_774),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_792),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_807),
.Y(n_828)
);

AO21x1_ASAP7_75t_L g829 ( 
.A1(n_812),
.A2(n_757),
.B(n_758),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_810),
.B(n_745),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_807),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_772),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_767),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_790),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_796),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_805),
.B(n_755),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_796),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_783),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_794),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_768),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_786),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_811),
.B(n_737),
.Y(n_842)
);

BUFx4f_ASAP7_75t_SL g843 ( 
.A(n_770),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_779),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_764),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_778),
.A2(n_760),
.B(n_762),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_788),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_776),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_775),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_779),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_797),
.B(n_349),
.Y(n_851)
);

AOI21x1_ASAP7_75t_L g852 ( 
.A1(n_773),
.A2(n_364),
.B(n_363),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_777),
.A2(n_361),
.B1(n_358),
.B2(n_354),
.Y(n_853)
);

BUFx2_ASAP7_75t_R g854 ( 
.A(n_789),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_781),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_775),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_773),
.A2(n_352),
.B(n_98),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_845),
.B(n_765),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_845),
.Y(n_859)
);

AO31x2_ASAP7_75t_L g860 ( 
.A1(n_840),
.A2(n_803),
.A3(n_804),
.B(n_778),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_835),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_R g862 ( 
.A(n_813),
.B(n_788),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_815),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_826),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_832),
.B(n_799),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_830),
.B(n_781),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_837),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_SL g868 ( 
.A1(n_836),
.A2(n_800),
.B(n_802),
.C(n_806),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_830),
.B(n_764),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_R g870 ( 
.A(n_847),
.B(n_795),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_834),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_828),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_831),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_851),
.B(n_808),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_843),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_SL g876 ( 
.A(n_842),
.B(n_809),
.C(n_787),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_822),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_SL g878 ( 
.A(n_836),
.B(n_809),
.C(n_787),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_824),
.B(n_798),
.Y(n_879)
);

BUFx4f_ASAP7_75t_SL g880 ( 
.A(n_827),
.Y(n_880)
);

XNOR2xp5_ASAP7_75t_L g881 ( 
.A(n_853),
.B(n_798),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_819),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_844),
.B(n_782),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_838),
.Y(n_884)
);

CKINVDCx16_ASAP7_75t_R g885 ( 
.A(n_823),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_820),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_843),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_850),
.B(n_96),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_855),
.B(n_99),
.Y(n_889)
);

AO21x2_ASAP7_75t_L g890 ( 
.A1(n_852),
.A2(n_105),
.B(n_106),
.Y(n_890)
);

BUFx4f_ASAP7_75t_SL g891 ( 
.A(n_820),
.Y(n_891)
);

AO31x2_ASAP7_75t_L g892 ( 
.A1(n_848),
.A2(n_109),
.A3(n_110),
.B(n_112),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

BUFx4f_ASAP7_75t_L g894 ( 
.A(n_821),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_816),
.B(n_116),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_818),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_861),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_867),
.B(n_817),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_866),
.B(n_839),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_887),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_884),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_869),
.B(n_839),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_871),
.B(n_817),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_872),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_874),
.B(n_877),
.Y(n_905)
);

BUFx4f_ASAP7_75t_SL g906 ( 
.A(n_875),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_873),
.B(n_825),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_863),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_896),
.B(n_833),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_864),
.B(n_833),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_884),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_879),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_SL g913 ( 
.A1(n_858),
.A2(n_856),
.B1(n_849),
.B2(n_846),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_SL g914 ( 
.A1(n_889),
.A2(n_846),
.B1(n_854),
.B2(n_814),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_883),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_860),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_860),
.B(n_841),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_862),
.B(n_885),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_892),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_870),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_892),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_892),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_868),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_888),
.B(n_821),
.Y(n_924)
);

AO21x2_ASAP7_75t_L g925 ( 
.A1(n_878),
.A2(n_857),
.B(n_841),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_881),
.B(n_829),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_876),
.B(n_895),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_886),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_893),
.Y(n_929)
);

BUFx6f_ASAP7_75t_SL g930 ( 
.A(n_859),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_911),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_920),
.B(n_865),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_897),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_901),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_912),
.B(n_890),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_902),
.B(n_905),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_901),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_929),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_904),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_926),
.B(n_890),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_908),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_899),
.B(n_882),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_903),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_914),
.A2(n_894),
.B1(n_891),
.B2(n_880),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_898),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_900),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_915),
.B(n_126),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_L g948 ( 
.A(n_923),
.B(n_913),
.C(n_927),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_916),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_910),
.B(n_132),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_927),
.B(n_136),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_916),
.B(n_919),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_918),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_907),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_918),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_924),
.B(n_218),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_943),
.B(n_917),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_953),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_941),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_931),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_955),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_940),
.B(n_921),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_936),
.B(n_922),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_933),
.B(n_917),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_949),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_946),
.B(n_914),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_932),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_937),
.B(n_909),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_939),
.B(n_925),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_942),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_945),
.B(n_925),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_934),
.B(n_935),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_949),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_954),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_960),
.Y(n_975)
);

OAI31xp33_ASAP7_75t_L g976 ( 
.A1(n_966),
.A2(n_944),
.A3(n_951),
.B(n_948),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_964),
.B(n_952),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_964),
.B(n_952),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_958),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_970),
.B(n_930),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_965),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_938),
.Y(n_982)
);

OAI222xp33_ASAP7_75t_L g983 ( 
.A1(n_961),
.A2(n_947),
.B1(n_950),
.B2(n_906),
.C1(n_938),
.C2(n_956),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_975),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_976),
.B(n_967),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_977),
.B(n_972),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_983),
.A2(n_969),
.B(n_971),
.Y(n_987)
);

AOI22x1_ASAP7_75t_L g988 ( 
.A1(n_979),
.A2(n_973),
.B1(n_974),
.B2(n_959),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_980),
.A2(n_957),
.B1(n_963),
.B2(n_968),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_977),
.A2(n_963),
.B1(n_962),
.B2(n_930),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_984),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_986),
.B(n_978),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_985),
.A2(n_982),
.B(n_981),
.Y(n_993)
);

AOI21xp33_ASAP7_75t_L g994 ( 
.A1(n_987),
.A2(n_990),
.B(n_988),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_989),
.B(n_938),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_991),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_995),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_997),
.A2(n_994),
.B(n_993),
.Y(n_998)
);

NOR2x1_ASAP7_75t_L g999 ( 
.A(n_996),
.B(n_992),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_998),
.B(n_928),
.C(n_929),
.Y(n_1000)
);

AND4x1_ASAP7_75t_L g1001 ( 
.A(n_999),
.B(n_158),
.C(n_162),
.D(n_164),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_1001),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_1000),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_1002),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_1003),
.B(n_167),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_1005),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_1004),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_1007),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1006),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1008),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_1009),
.Y(n_1011)
);

AOI22x1_ASAP7_75t_L g1012 ( 
.A1(n_1011),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1010),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1013),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1015),
.B(n_1014),
.Y(n_1016)
);

XNOR2xp5_ASAP7_75t_L g1017 ( 
.A(n_1015),
.B(n_1012),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_1016),
.A2(n_194),
.B1(n_196),
.B2(n_198),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_SL g1019 ( 
.A1(n_1017),
.A2(n_199),
.B1(n_202),
.B2(n_205),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_1019),
.B(n_206),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_1018),
.B1(n_209),
.B2(n_210),
.Y(n_1021)
);


endmodule