module fake_jpeg_25801_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_1),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_18),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_11),
.Y(n_22)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_24),
.B1(n_17),
.B2(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_11),
.B1(n_13),
.B2(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_13),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_14),
.B(n_12),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_25),
.B(n_28),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_24),
.B(n_27),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_21),
.C(n_9),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_26),
.B(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_5),
.B1(n_18),
.B2(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_33),
.B(n_30),
.Y(n_40)
);

NOR4xp25_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_39),
.C(n_32),
.D(n_29),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_31),
.B(n_34),
.C(n_26),
.Y(n_42)
);


endmodule