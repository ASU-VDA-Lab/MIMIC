module real_aes_15650_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g116 ( .A(n_0), .B(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_1), .A2(n_4), .B1(n_214), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_2), .A2(n_45), .B1(n_152), .B2(n_154), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_3), .A2(n_25), .B1(n_154), .B2(n_178), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_5), .A2(n_16), .B1(n_195), .B2(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_6), .A2(n_62), .B1(n_180), .B2(n_252), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_7), .A2(n_17), .B1(n_152), .B2(n_199), .Y(n_521) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_9), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_10), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_11), .A2(n_18), .B1(n_197), .B2(n_251), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_12), .A2(n_66), .B1(n_822), .B2(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_12), .Y(n_822) );
OR2x2_ASAP7_75t_L g112 ( .A(n_13), .B(n_40), .Y(n_112) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_15), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_19), .A2(n_101), .B1(n_195), .B2(n_214), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_20), .A2(n_488), .B(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_21), .A2(n_41), .B1(n_228), .B2(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_22), .B(n_196), .Y(n_269) );
OAI22x1_ASAP7_75t_SL g819 ( .A1(n_23), .A2(n_820), .B1(n_821), .B2(n_824), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_23), .Y(n_824) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_24), .A2(n_60), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_26), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_27), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_28), .B(n_158), .Y(n_545) );
INVx4_ASAP7_75t_R g534 ( .A(n_29), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_30), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_31), .A2(n_49), .B1(n_160), .B2(n_162), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_32), .A2(n_56), .B1(n_162), .B2(n_195), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_33), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_34), .B(n_228), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_35), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_36), .B(n_154), .Y(n_552) );
INVx1_ASAP7_75t_L g600 ( .A(n_37), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_SL g581 ( .A1(n_38), .A2(n_152), .B(n_164), .C(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_39), .A2(n_57), .B1(n_152), .B2(n_162), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_42), .A2(n_89), .B1(n_152), .B2(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_43), .A2(n_55), .B1(n_137), .B2(n_138), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_43), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_44), .A2(n_48), .B1(n_152), .B2(n_199), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_46), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_47), .A2(n_61), .B1(n_195), .B2(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g549 ( .A(n_50), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_51), .B(n_152), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_52), .Y(n_562) );
INVx2_ASAP7_75t_L g122 ( .A(n_53), .Y(n_122) );
BUFx3_ASAP7_75t_L g111 ( .A(n_54), .Y(n_111) );
INVx1_ASAP7_75t_L g132 ( .A(n_54), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_55), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_58), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_59), .A2(n_90), .B1(n_152), .B2(n_162), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_63), .A2(n_78), .B1(n_160), .B2(n_217), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_64), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_65), .A2(n_80), .B1(n_152), .B2(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g823 ( .A(n_66), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_67), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_68), .A2(n_100), .B1(n_195), .B2(n_197), .Y(n_194) );
AND2x4_ASAP7_75t_L g148 ( .A(n_69), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g169 ( .A(n_70), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_71), .A2(n_92), .B1(n_160), .B2(n_162), .Y(n_596) );
AO22x1_ASAP7_75t_L g510 ( .A1(n_72), .A2(n_79), .B1(n_229), .B2(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g149 ( .A(n_73), .Y(n_149) );
AND2x2_ASAP7_75t_L g584 ( .A(n_74), .B(n_166), .Y(n_584) );
CKINVDCx14_ASAP7_75t_R g126 ( .A(n_75), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_75), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_76), .B(n_180), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_77), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_81), .B(n_154), .Y(n_563) );
INVx2_ASAP7_75t_L g158 ( .A(n_82), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_83), .B(n_166), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_84), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_85), .A2(n_99), .B1(n_162), .B2(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_86), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_87), .B(n_187), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_88), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_91), .B(n_166), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_93), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_94), .B(n_166), .Y(n_559) );
INVx1_ASAP7_75t_L g115 ( .A(n_95), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_95), .B(n_131), .Y(n_130) );
NAND2xp33_ASAP7_75t_L g272 ( .A(n_96), .B(n_196), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_97), .A2(n_180), .B(n_182), .C(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g536 ( .A(n_98), .B(n_537), .Y(n_536) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_102), .B(n_161), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_118), .B(n_833), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_107), .Y(n_835) );
BUFx12f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_113), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g832 ( .A(n_110), .B(n_817), .Y(n_832) );
NOR2x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g497 ( .A(n_111), .Y(n_497) );
INVx1_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g817 ( .A(n_115), .Y(n_817) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_491), .Y(n_118) );
NOR2x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
BUFx8_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g495 ( .A(n_122), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_122), .B(n_831), .Y(n_830) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_483), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_134), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
CKINVDCx8_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g487 ( .A(n_129), .Y(n_487) );
INVx5_ASAP7_75t_L g490 ( .A(n_129), .Y(n_490) );
AND2x6_ASAP7_75t_SL g129 ( .A(n_130), .B(n_133), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_133), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AOI21xp33_ASAP7_75t_SL g483 ( .A1(n_135), .A2(n_484), .B(n_488), .Y(n_483) );
XNOR2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_139), .Y(n_135) );
OAI22x1_ASAP7_75t_L g500 ( .A1(n_139), .A2(n_501), .B1(n_815), .B2(n_818), .Y(n_500) );
NOR2x1p5_ASAP7_75t_L g139 ( .A(n_140), .B(n_393), .Y(n_139) );
NAND4xp75_ASAP7_75t_L g140 ( .A(n_141), .B(n_338), .C(n_358), .D(n_374), .Y(n_140) );
NOR2x1p5_ASAP7_75t_SL g141 ( .A(n_142), .B(n_308), .Y(n_141) );
NAND4xp75_ASAP7_75t_L g142 ( .A(n_143), .B(n_244), .C(n_285), .D(n_294), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_205), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_172), .Y(n_144) );
AND2x4_ASAP7_75t_L g418 ( .A(n_145), .B(n_345), .Y(n_418) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_146), .Y(n_261) );
INVx2_ASAP7_75t_L g279 ( .A(n_146), .Y(n_279) );
AND2x2_ASAP7_75t_L g302 ( .A(n_146), .B(n_264), .Y(n_302) );
OR2x2_ASAP7_75t_L g357 ( .A(n_146), .B(n_173), .Y(n_357) );
AO31x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .A3(n_165), .B(n_170), .Y(n_146) );
INVx2_ASAP7_75t_L g202 ( .A(n_147), .Y(n_202) );
AO31x2_ASAP7_75t_L g225 ( .A1(n_147), .A2(n_174), .A3(n_226), .B(n_234), .Y(n_225) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_147), .A2(n_191), .A3(n_249), .B(n_255), .Y(n_248) );
AO31x2_ASAP7_75t_L g519 ( .A1(n_147), .A2(n_222), .A3(n_520), .B(n_523), .Y(n_519) );
BUFx10_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
INVx1_ASAP7_75t_L g517 ( .A(n_148), .Y(n_517) );
BUFx10_ASAP7_75t_L g554 ( .A(n_148), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B1(n_159), .B2(n_163), .Y(n_150) );
INVx1_ASAP7_75t_L g197 ( .A(n_152), .Y(n_197) );
INVx4_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
INVx1_ASAP7_75t_L g217 ( .A(n_152), .Y(n_217) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_153), .Y(n_154) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
INVx2_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx1_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
INVx1_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
INVx1_ASAP7_75t_L g230 ( .A(n_153), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_153), .Y(n_233) );
INVx1_ASAP7_75t_L g253 ( .A(n_153), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_154), .B(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_155), .A2(n_163), .B1(n_213), .B2(n_216), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_155), .A2(n_163), .B1(n_227), .B2(n_231), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_155), .A2(n_163), .B1(n_240), .B2(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g513 ( .A(n_156), .Y(n_513) );
BUFx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g565 ( .A(n_157), .Y(n_565) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx8_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
INVx1_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
INVx1_ASAP7_75t_L g548 ( .A(n_158), .Y(n_548) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g228 ( .A(n_161), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_161), .A2(n_233), .B1(n_534), .B2(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_162), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g598 ( .A(n_162), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_163), .A2(n_176), .B1(n_179), .B2(n_181), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_163), .A2(n_194), .B1(n_198), .B2(n_200), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_163), .A2(n_200), .B1(n_250), .B2(n_254), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_163), .A2(n_271), .B(n_272), .Y(n_270) );
OAI22x1_ASAP7_75t_L g520 ( .A1(n_163), .A2(n_181), .B1(n_521), .B2(n_522), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_163), .A2(n_513), .B1(n_588), .B2(n_589), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_163), .A2(n_181), .B1(n_596), .B2(n_597), .Y(n_595) );
INVx6_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g267 ( .A1(n_164), .A2(n_199), .B(n_268), .C(n_269), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_164), .A2(n_510), .B(n_512), .C(n_516), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_164), .A2(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_164), .B(n_510), .Y(n_612) );
AO31x2_ASAP7_75t_L g586 ( .A1(n_165), .A2(n_554), .A3(n_587), .B(n_590), .Y(n_586) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_166), .B(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_167), .B(n_171), .Y(n_170) );
BUFx3_ASAP7_75t_L g174 ( .A(n_167), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_167), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_167), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_SL g265 ( .A(n_167), .Y(n_265) );
AND2x2_ASAP7_75t_L g553 ( .A(n_167), .B(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
AND2x2_ASAP7_75t_L g275 ( .A(n_172), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g425 ( .A(n_172), .B(n_302), .Y(n_425) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_189), .Y(n_172) );
OR2x2_ASAP7_75t_L g262 ( .A(n_173), .B(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g293 ( .A(n_173), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_173), .B(n_190), .Y(n_299) );
INVx1_ASAP7_75t_L g317 ( .A(n_173), .Y(n_317) );
INVx2_ASAP7_75t_L g346 ( .A(n_173), .Y(n_346) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .A3(n_183), .B(n_185), .Y(n_173) );
INVx2_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_178), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_181), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_SL g200 ( .A(n_182), .Y(n_200) );
AO31x2_ASAP7_75t_L g238 ( .A1(n_183), .A2(n_218), .A3(n_239), .B(n_242), .Y(n_238) );
AO31x2_ASAP7_75t_L g594 ( .A1(n_183), .A2(n_191), .A3(n_595), .B(n_599), .Y(n_594) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_SL g273 ( .A(n_184), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
INVx2_ASAP7_75t_L g219 ( .A(n_186), .Y(n_219) );
NOR2xp33_ASAP7_75t_SL g255 ( .A(n_186), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g192 ( .A(n_187), .Y(n_192) );
INVx2_ASAP7_75t_L g222 ( .A(n_187), .Y(n_222) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_187), .A2(n_515), .B(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g322 ( .A(n_189), .Y(n_322) );
INVx2_ASAP7_75t_L g327 ( .A(n_189), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_189), .B(n_278), .Y(n_332) );
AND2x2_ASAP7_75t_L g355 ( .A(n_189), .B(n_334), .Y(n_355) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_189), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_189), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g344 ( .A(n_190), .Y(n_344) );
AND2x2_ASAP7_75t_L g392 ( .A(n_190), .B(n_346), .Y(n_392) );
AO31x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .A3(n_201), .B(n_203), .Y(n_190) );
AOI21x1_ASAP7_75t_L g573 ( .A1(n_191), .A2(n_574), .B(n_584), .Y(n_573) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_192), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g537 ( .A(n_192), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_192), .B(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_192), .B(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_196), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_199), .A2(n_562), .B(n_563), .C(n_564), .Y(n_561) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_201), .A2(n_212), .A3(n_218), .B(n_220), .Y(n_211) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_202), .A2(n_529), .B(n_532), .Y(n_528) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_223), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_207), .B(n_336), .Y(n_383) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_208), .B(n_336), .Y(n_380) );
INVx1_ASAP7_75t_L g481 ( .A(n_208), .Y(n_481) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g431 ( .A(n_209), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
OR2x2_ASAP7_75t_L g365 ( .A(n_210), .B(n_237), .Y(n_365) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g307 ( .A(n_211), .Y(n_307) );
AND2x4_ASAP7_75t_L g313 ( .A(n_211), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_215), .B(n_579), .Y(n_578) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_218), .A2(n_528), .B(n_536), .Y(n_527) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_222), .B(n_243), .Y(n_242) );
AOI32xp33_ASAP7_75t_L g451 ( .A1(n_223), .A2(n_354), .A3(n_452), .B1(n_454), .B2(n_455), .Y(n_451) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g400 ( .A(n_224), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_236), .Y(n_224) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_225), .Y(n_246) );
OR2x2_ASAP7_75t_L g282 ( .A(n_225), .B(n_238), .Y(n_282) );
INVx1_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
AND2x2_ASAP7_75t_L g306 ( .A(n_225), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g312 ( .A(n_225), .Y(n_312) );
INVx2_ASAP7_75t_L g337 ( .A(n_225), .Y(n_337) );
AND2x2_ASAP7_75t_L g456 ( .A(n_225), .B(n_248), .Y(n_456) );
OAI21xp33_ASAP7_75t_SL g544 ( .A1(n_229), .A2(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_236), .B(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g247 ( .A(n_238), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
INVx2_ASAP7_75t_L g314 ( .A(n_238), .Y(n_314) );
AND2x4_ASAP7_75t_L g336 ( .A(n_238), .B(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_238), .Y(n_428) );
AOI22x1_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_257), .B1(n_275), .B2(n_280), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND4xp25_ASAP7_75t_L g405 ( .A(n_247), .B(n_406), .C(n_407), .D(n_408), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_247), .B(n_306), .Y(n_436) );
INVx4_ASAP7_75t_SL g289 ( .A(n_248), .Y(n_289) );
BUFx2_ASAP7_75t_L g352 ( .A(n_248), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_248), .B(n_297), .Y(n_415) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_253), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g377 ( .A(n_259), .B(n_326), .Y(n_377) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g300 ( .A(n_263), .B(n_278), .Y(n_300) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_264), .B(n_279), .Y(n_324) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_274), .Y(n_264) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_265), .A2(n_266), .B(n_274), .Y(n_319) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_273), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_276), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g342 ( .A(n_276), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g381 ( .A(n_277), .B(n_299), .Y(n_381) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g424 ( .A(n_279), .B(n_334), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_280), .A2(n_397), .B1(n_399), .B2(n_402), .C(n_404), .Y(n_396) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g290 ( .A(n_282), .Y(n_290) );
OR2x2_ASAP7_75t_L g390 ( .A(n_282), .B(n_329), .Y(n_390) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_286), .A2(n_412), .B1(n_416), .B2(n_419), .Y(n_411) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
AND2x4_ASAP7_75t_L g335 ( .A(n_287), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g447 ( .A(n_287), .B(n_365), .Y(n_447) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g295 ( .A(n_289), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_289), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g370 ( .A(n_289), .B(n_307), .Y(n_370) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_289), .Y(n_387) );
INVx1_ASAP7_75t_L g401 ( .A(n_289), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_289), .B(n_314), .Y(n_444) );
AND2x4_ASAP7_75t_L g351 ( .A(n_290), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g349 ( .A(n_292), .Y(n_349) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_293), .B(n_334), .Y(n_333) );
NAND2x1_ASAP7_75t_L g453 ( .A(n_293), .B(n_355), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .B1(n_301), .B2(n_303), .Y(n_294) );
AND2x2_ASAP7_75t_L g320 ( .A(n_295), .B(n_313), .Y(n_320) );
INVx1_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
AND2x2_ASAP7_75t_L g468 ( .A(n_295), .B(n_329), .Y(n_468) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x2_ASAP7_75t_L g301 ( .A(n_299), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g441 ( .A(n_299), .Y(n_441) );
AND2x2_ASAP7_75t_L g458 ( .A(n_299), .B(n_318), .Y(n_458) );
AND2x2_ASAP7_75t_L g474 ( .A(n_299), .B(n_424), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_300), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g397 ( .A(n_300), .B(n_398), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_300), .A2(n_390), .B1(n_405), .B2(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
AND2x2_ASAP7_75t_L g391 ( .A(n_302), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_302), .B(n_398), .Y(n_420) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g426 ( .A(n_306), .B(n_427), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_306), .A2(n_330), .B1(n_435), .B2(n_437), .Y(n_434) );
INVx3_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
AND2x2_ASAP7_75t_L g461 ( .A(n_307), .B(n_314), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_325), .Y(n_308) );
AOI32xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_315), .A3(n_318), .B1(n_320), .B2(n_321), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_312), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_312), .Y(n_432) );
INVx3_ASAP7_75t_L g388 ( .A(n_313), .Y(n_388) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_316), .A2(n_464), .B1(n_465), .B2(n_466), .C(n_467), .Y(n_463) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g440 ( .A(n_318), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g476 ( .A(n_318), .B(n_437), .Y(n_476) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_321), .B(n_349), .Y(n_348) );
AO22x1_ASAP7_75t_L g378 ( .A1(n_321), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_321), .B(n_349), .Y(n_482) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g398 ( .A(n_322), .Y(n_398) );
INVx1_ASAP7_75t_L g408 ( .A(n_322), .Y(n_408) );
AND2x2_ASAP7_75t_L g328 ( .A(n_323), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_324), .Y(n_410) );
INVx1_ASAP7_75t_L g450 ( .A(n_324), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_330), .C(n_335), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2x1p5_ASAP7_75t_L g437 ( .A(n_327), .B(n_357), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_328), .B(n_387), .Y(n_464) );
AOI31xp33_ASAP7_75t_L g347 ( .A1(n_329), .A2(n_348), .A3(n_350), .B(n_353), .Y(n_347) );
INVx4_ASAP7_75t_L g406 ( .A(n_329), .Y(n_406) );
OR2x2_ASAP7_75t_L g443 ( .A(n_329), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x4_ASAP7_75t_L g345 ( .A(n_334), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_336), .Y(n_341) );
AND2x2_ASAP7_75t_L g372 ( .A(n_336), .B(n_370), .Y(n_372) );
NOR2xp67_ASAP7_75t_L g338 ( .A(n_339), .B(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g465 ( .A(n_342), .Y(n_465) );
INVx1_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g403 ( .A(n_344), .Y(n_403) );
AND2x2_ASAP7_75t_L g402 ( .A(n_345), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .A3(n_362), .B1(n_366), .B2(n_369), .C1(n_371), .C2(n_373), .Y(n_359) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI211x1_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_378), .C(n_384), .Y(n_374) );
INVx1_ASAP7_75t_L g479 ( .A(n_375), .Y(n_479) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B(n_391), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx2_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp33_ASAP7_75t_L g449 ( .A(n_392), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_462), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_429), .C(n_445), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_411), .C(n_421), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_398), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_402), .A2(n_458), .B(n_459), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_406), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_406), .B(n_456), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_407), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_408), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_418), .A2(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_434), .C(n_438), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_440), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_444), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_451), .C(n_457), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_456), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g477 ( .A(n_456), .Y(n_477) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g473 ( .A(n_461), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .C(n_478), .Y(n_462) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI21xp33_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_475), .B(n_477), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AOI21xp33_ASAP7_75t_R g478 ( .A1(n_479), .A2(n_480), .B(n_482), .Y(n_478) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_498), .B(n_826), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
BUFx12f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x6_ASAP7_75t_SL g494 ( .A(n_495), .B(n_496), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_819), .B2(n_825), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_725), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_654), .C(n_696), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_628), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_538), .B1(n_603), .B2(n_614), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_525), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_507), .A2(n_648), .B(n_650), .Y(n_647) );
AOI21xp33_ASAP7_75t_L g720 ( .A1(n_507), .A2(n_721), .B(n_722), .Y(n_720) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
INVx2_ASAP7_75t_L g640 ( .A(n_508), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_508), .B(n_519), .Y(n_670) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g611 ( .A(n_512), .Y(n_611) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_513), .A2(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g613 ( .A(n_516), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_517), .A2(n_575), .B(n_581), .Y(n_574) );
AND2x2_ASAP7_75t_L g710 ( .A(n_518), .B(n_557), .Y(n_710) );
INVx1_ASAP7_75t_L g743 ( .A(n_518), .Y(n_743) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g605 ( .A(n_519), .B(n_558), .Y(n_605) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g645 ( .A(n_519), .Y(n_645) );
OR2x2_ASAP7_75t_L g664 ( .A(n_519), .B(n_527), .Y(n_664) );
AND2x2_ASAP7_75t_L g679 ( .A(n_519), .B(n_527), .Y(n_679) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_526), .B(n_678), .Y(n_721) );
OR2x2_ASAP7_75t_L g809 ( .A(n_526), .B(n_670), .Y(n_809) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g637 ( .A(n_527), .Y(n_637) );
AND2x2_ASAP7_75t_L g646 ( .A(n_527), .B(n_609), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_527), .B(n_558), .Y(n_649) );
AND2x2_ASAP7_75t_L g668 ( .A(n_527), .B(n_557), .Y(n_668) );
AND2x4_ASAP7_75t_L g687 ( .A(n_527), .B(n_610), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_555), .B(n_592), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_539), .B(n_682), .Y(n_785) );
CKINVDCx14_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_541), .B(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g618 ( .A(n_541), .Y(n_618) );
OR2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_541), .B(n_619), .Y(n_651) );
AND2x2_ASAP7_75t_L g676 ( .A(n_541), .B(n_594), .Y(n_676) );
AND2x2_ASAP7_75t_L g694 ( .A(n_541), .B(n_624), .Y(n_694) );
INVx1_ASAP7_75t_L g733 ( .A(n_541), .Y(n_733) );
AND2x2_ASAP7_75t_L g735 ( .A(n_541), .B(n_736), .Y(n_735) );
NAND2x1p5_ASAP7_75t_SL g754 ( .A(n_541), .B(n_675), .Y(n_754) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_550), .B(n_553), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_548), .Y(n_580) );
INVx1_ASAP7_75t_L g570 ( .A(n_554), .Y(n_570) );
OAI32xp33_ASAP7_75t_L g638 ( .A1(n_555), .A2(n_630), .A3(n_639), .B1(n_641), .B2(n_643), .Y(n_638) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_571), .Y(n_555) );
INVx1_ASAP7_75t_L g678 ( .A(n_556), .Y(n_678) );
AND2x2_ASAP7_75t_L g686 ( .A(n_556), .B(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g685 ( .A(n_557), .B(n_609), .Y(n_685) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx3_ASAP7_75t_L g635 ( .A(n_558), .Y(n_635) );
AND2x2_ASAP7_75t_L g644 ( .A(n_558), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g750 ( .A(n_558), .Y(n_750) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_566), .B(n_569), .Y(n_560) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g620 ( .A(n_571), .Y(n_620) );
OR2x2_ASAP7_75t_L g630 ( .A(n_571), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g752 ( .A(n_571), .Y(n_752) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_585), .Y(n_571) );
AND2x2_ASAP7_75t_L g653 ( .A(n_572), .B(n_586), .Y(n_653) );
INVx2_ASAP7_75t_L g675 ( .A(n_572), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_572), .B(n_594), .Y(n_695) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g602 ( .A(n_573), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B(n_580), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_585), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g684 ( .A(n_585), .Y(n_684) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g624 ( .A(n_586), .Y(n_624) );
OR2x2_ASAP7_75t_L g690 ( .A(n_586), .B(n_594), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_586), .B(n_594), .Y(n_723) );
INVx2_ASAP7_75t_L g671 ( .A(n_592), .Y(n_671) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_601), .Y(n_592) );
OR2x2_ASAP7_75t_L g658 ( .A(n_593), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g736 ( .A(n_593), .Y(n_736) );
INVx1_ASAP7_75t_L g619 ( .A(n_594), .Y(n_619) );
INVx1_ASAP7_75t_L g627 ( .A(n_594), .Y(n_627) );
INVx1_ASAP7_75t_L g642 ( .A(n_594), .Y(n_642) );
OR2x2_ASAP7_75t_L g746 ( .A(n_601), .B(n_723), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_602), .B(n_618), .Y(n_659) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_602), .Y(n_661) );
OR2x2_ASAP7_75t_L g760 ( .A(n_602), .B(n_684), .Y(n_760) );
INVxp67_ASAP7_75t_L g784 ( .A(n_602), .Y(n_784) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_605), .B(n_646), .Y(n_713) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g662 ( .A(n_607), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g775 ( .A(n_608), .Y(n_775) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g804 ( .A(n_609), .B(n_637), .Y(n_804) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g730 ( .A(n_610), .B(n_637), .Y(n_730) );
AOI21x1_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B(n_613), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_617), .B(n_653), .Y(n_767) );
AND2x4_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx2_ASAP7_75t_L g631 ( .A(n_618), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_618), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_618), .B(n_675), .Y(n_724) );
OR2x2_ASAP7_75t_L g796 ( .A(n_618), .B(n_683), .Y(n_796) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g716 ( .A(n_622), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx2_ASAP7_75t_L g707 ( .A(n_623), .Y(n_707) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g697 ( .A(n_626), .B(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_626), .Y(n_708) );
OR2x2_ASAP7_75t_L g759 ( .A(n_626), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g814 ( .A(n_626), .Y(n_814) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_632), .B(n_638), .C(n_647), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g703 ( .A(n_631), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_631), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g776 ( .A(n_631), .B(n_653), .Y(n_776) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_634), .B(n_679), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g718 ( .A(n_634), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g786 ( .A(n_634), .B(n_787), .Y(n_786) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g729 ( .A(n_635), .Y(n_729) );
AND2x2_ASAP7_75t_L g757 ( .A(n_636), .B(n_685), .Y(n_757) );
INVx2_ASAP7_75t_L g780 ( .A(n_636), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_636), .B(n_678), .Y(n_812) );
AND2x4_ASAP7_75t_SL g766 ( .A(n_639), .B(n_644), .Y(n_766) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g719 ( .A(n_640), .B(n_645), .Y(n_719) );
OR2x2_ASAP7_75t_L g771 ( .A(n_640), .B(n_664), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_641), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_641), .B(n_653), .Y(n_807) );
BUFx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g755 ( .A(n_642), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g738 ( .A(n_644), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_644), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g788 ( .A(n_645), .Y(n_788) );
BUFx2_ASAP7_75t_L g656 ( .A(n_646), .Y(n_656) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g774 ( .A(n_649), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g698 ( .A(n_653), .Y(n_698) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_653), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_665), .C(n_680), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_657), .B1(n_660), .B2(n_662), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI222xp33_ASAP7_75t_L g768 ( .A1(n_662), .A2(n_688), .B1(n_769), .B2(n_772), .C1(n_774), .C2(n_776), .Y(n_768) );
AND2x2_ASAP7_75t_L g800 ( .A(n_663), .B(n_749), .Y(n_800) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g748 ( .A(n_664), .B(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_671), .B1(n_672), .B2(n_677), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx2_ASAP7_75t_SL g744 ( .A(n_668), .Y(n_744) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
AND2x2_ASAP7_75t_L g731 ( .A(n_673), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g689 ( .A(n_674), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g683 ( .A(n_675), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g798 ( .A(n_676), .Y(n_798) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_679), .B(n_775), .Y(n_794) );
INVx1_ASAP7_75t_L g811 ( .A(n_679), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B1(n_686), .B2(n_688), .C1(n_691), .C2(n_692), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_687), .Y(n_691) );
AND2x2_ASAP7_75t_L g709 ( .A(n_687), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g740 ( .A(n_687), .Y(n_740) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g704 ( .A(n_690), .Y(n_704) );
OR2x2_ASAP7_75t_L g773 ( .A(n_690), .B(n_754), .Y(n_773) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_702), .C(n_711), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_709), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_703), .A2(n_741), .B1(n_790), .B2(n_793), .C(n_795), .Y(n_789) );
AND2x4_ASAP7_75t_L g732 ( .A(n_704), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g763 ( .A(n_710), .Y(n_763) );
AOI211x1_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_716), .C(n_720), .Y(n_711) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g781 ( .A(n_719), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_722), .B(n_770), .C(n_771), .Y(n_769) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g805 ( .A(n_723), .Y(n_805) );
NOR2x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_777), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g726 ( .A(n_727), .B(n_734), .C(n_756), .D(n_768), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_731), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g787 ( .A(n_730), .B(n_788), .Y(n_787) );
AOI221x1_ASAP7_75t_L g756 ( .A1(n_732), .A2(n_757), .B1(n_758), .B2(n_761), .C(n_764), .Y(n_756) );
AND2x2_ASAP7_75t_L g782 ( .A(n_732), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g792 ( .A(n_733), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B1(n_741), .B2(n_745), .C(n_747), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_739), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_744), .A2(n_748), .B1(n_751), .B2(n_753), .Y(n_747) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_748), .A2(n_765), .B(n_767), .Y(n_764) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g770 ( .A(n_750), .Y(n_770) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVxp67_ASAP7_75t_L g791 ( .A(n_760), .Y(n_791) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_773), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_789), .C(n_801), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_782), .B1(n_785), .B2(n_786), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g797 ( .A(n_784), .B(n_798), .Y(n_797) );
NAND2x1_ASAP7_75t_L g813 ( .A(n_784), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B(n_799), .Y(n_795) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_805), .B1(n_806), .B2(n_808), .C(n_810), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx3_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
INVx4_ASAP7_75t_L g818 ( .A(n_815), .Y(n_818) );
BUFx12f_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_819), .Y(n_825) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
BUFx10_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_SL g833 ( .A(n_834), .B(n_835), .Y(n_833) );
endmodule