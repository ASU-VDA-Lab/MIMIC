module fake_ariane_3149_n_1563 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1563);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1563;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_2),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_8),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_59),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_54),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_39),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_35),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_31),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_17),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_21),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_8),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_37),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_58),
.Y(n_172)
);

BUFx8_ASAP7_75t_SL g173 ( 
.A(n_127),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_69),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_43),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_49),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_67),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_12),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_26),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_29),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_55),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_88),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_19),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_12),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_48),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_52),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_63),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_46),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_56),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_50),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_42),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_46),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_87),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_75),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_62),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_39),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_138),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_94),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_66),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_5),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_21),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_102),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_47),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_98),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_28),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_36),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_130),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_31),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_19),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_60),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_105),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_30),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_77),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_107),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_68),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_76),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_22),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_72),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_117),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_85),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_65),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_80),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_0),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_40),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_115),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_91),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_96),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_73),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_89),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_42),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_139),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_23),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_53),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_16),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_15),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_51),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_95),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_29),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_37),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_122),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_22),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_90),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_48),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_109),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_148),
.B(n_1),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_147),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_192),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_1),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_173),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_187),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_204),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_150),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_189),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_171),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_192),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_151),
.B(n_4),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_212),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_183),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_147),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_159),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_170),
.B(n_180),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_216),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_188),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_194),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_159),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_175),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_162),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_199),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_154),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_175),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_203),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_206),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_196),
.B(n_4),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_195),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_216),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_195),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_154),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_202),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_217),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_202),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_243),
.B(n_5),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_223),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_244),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_210),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_226),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_228),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_274),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_163),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_166),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_160),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_230),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_167),
.B(n_6),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_144),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_144),
.Y(n_348)
);

BUFx6f_ASAP7_75t_SL g349 ( 
.A(n_189),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_216),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_292),
.B(n_189),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_198),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_299),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_292),
.B(n_262),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_284),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_304),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_286),
.B(n_262),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_305),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_312),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_313),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_319),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_R g373 ( 
.A(n_293),
.B(n_296),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_328),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_336),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_295),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_294),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_302),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_337),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_301),
.B(n_212),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_341),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

BUFx10_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_298),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_301),
.B(n_145),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_309),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_303),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_310),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_281),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_316),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_301),
.B(n_246),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_294),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_347),
.B(n_153),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_320),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_321),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_306),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_348),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_348),
.B(n_164),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_306),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_311),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_366),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_329),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_366),
.B(n_330),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_360),
.B(n_274),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_342),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_372),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_394),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_333),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

NOR3xp33_ASAP7_75t_L g432 ( 
.A(n_362),
.B(n_300),
.C(n_283),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_361),
.B(n_338),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_396),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_398),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_356),
.B(n_318),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_413),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_387),
.B(n_339),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_387),
.B(n_343),
.Y(n_442)
);

NOR2x1p5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_340),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_345),
.Y(n_444)
);

BUFx4f_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_307),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_401),
.A2(n_322),
.B1(n_349),
.B2(n_287),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_323),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

NOR2x1p5_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_408),
.Y(n_453)
);

INVx4_ASAP7_75t_SL g454 ( 
.A(n_381),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_403),
.Y(n_455)
);

OAI21xp33_ASAP7_75t_SL g456 ( 
.A1(n_352),
.A2(n_332),
.B(n_287),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_368),
.B(n_169),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_352),
.B(n_323),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_383),
.B(n_344),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_332),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_369),
.B(n_315),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_369),
.B(n_176),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_165),
.C(n_161),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_374),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_399),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_378),
.B(n_177),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g474 ( 
.A1(n_351),
.A2(n_197),
.B1(n_267),
.B2(n_186),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_382),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_382),
.B(n_325),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_385),
.B(n_311),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_363),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_364),
.B(n_314),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_391),
.A2(n_197),
.B1(n_177),
.B2(n_267),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_392),
.B(n_184),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_R g485 ( 
.A(n_367),
.B(n_161),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_392),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_393),
.B(n_325),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_376),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_393),
.B(n_327),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_376),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_376),
.A2(n_346),
.B1(n_275),
.B2(n_234),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_380),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_409),
.B(n_193),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_370),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_390),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_381),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_L g499 ( 
.A1(n_406),
.A2(n_218),
.B1(n_165),
.B2(n_263),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_380),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_406),
.B(n_346),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_412),
.B(n_331),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_389),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_380),
.B(n_331),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_358),
.A2(n_259),
.B1(n_239),
.B2(n_279),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

OR2x6_ASAP7_75t_SL g508 ( 
.A(n_371),
.B(n_263),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_389),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_411),
.B(n_334),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_389),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_353),
.A2(n_248),
.B1(n_265),
.B2(n_213),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_412),
.B(n_334),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_353),
.B(n_317),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_389),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_389),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_353),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g519 ( 
.A1(n_354),
.A2(n_201),
.B(n_237),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_386),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_404),
.B(n_335),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_404),
.B(n_354),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_411),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_395),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_395),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_355),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_355),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_404),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_404),
.B(n_200),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_404),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_414),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_397),
.B(n_207),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_410),
.B(n_155),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_241),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_416),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_416),
.A2(n_269),
.B1(n_261),
.B2(n_262),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_377),
.B(n_211),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_379),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_388),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_359),
.B(n_246),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_352),
.B(n_214),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_357),
.B(n_225),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_362),
.B(n_251),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_359),
.B(n_276),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_366),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_SL g550 ( 
.A(n_394),
.B(n_253),
.C(n_278),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_523),
.B(n_155),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_442),
.B(n_276),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_523),
.B(n_156),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_459),
.B(n_157),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_417),
.A2(n_264),
.B1(n_158),
.B2(n_233),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_420),
.B(n_252),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_426),
.A2(n_280),
.B1(n_193),
.B2(n_256),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_418),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_482),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_462),
.B(n_158),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_417),
.B(n_549),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_264),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_545),
.B(n_272),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_466),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_426),
.A2(n_503),
.B1(n_511),
.B2(n_432),
.Y(n_571)
);

INVx8_ASAP7_75t_L g572 ( 
.A(n_422),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_445),
.B(n_227),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_423),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_501),
.B(n_273),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_445),
.B(n_229),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_430),
.B(n_232),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_425),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_434),
.B(n_277),
.Y(n_579)
);

NAND4xp25_ASAP7_75t_SL g580 ( 
.A(n_483),
.B(n_235),
.C(n_245),
.D(n_271),
.Y(n_580)
);

AND3x1_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_280),
.C(n_9),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_501),
.B(n_146),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_437),
.B(n_149),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_453),
.B(n_185),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_501),
.B(n_152),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_428),
.B(n_168),
.Y(n_587)
);

NOR2x1p5_ASAP7_75t_L g588 ( 
.A(n_428),
.B(n_172),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_468),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_434),
.B(n_7),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_440),
.B(n_7),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_424),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_424),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_444),
.B(n_9),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_468),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_485),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_446),
.B(n_10),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_419),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_424),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_450),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_421),
.B(n_174),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_480),
.B(n_10),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_503),
.B(n_179),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_442),
.A2(n_270),
.B1(n_260),
.B2(n_258),
.Y(n_604)
);

INVxp33_ASAP7_75t_SL g605 ( 
.A(n_496),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_438),
.B(n_11),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_490),
.B(n_221),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_460),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_222),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_488),
.B(n_514),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_476),
.A2(n_481),
.B(n_477),
.C(n_475),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_511),
.A2(n_250),
.B1(n_182),
.B2(n_181),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_524),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_525),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_511),
.A2(n_219),
.B1(n_190),
.B2(n_191),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_451),
.B(n_11),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_449),
.B(n_236),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_456),
.B(n_238),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_516),
.A2(n_242),
.B(n_255),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_544),
.B(n_13),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_466),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_544),
.B(n_205),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_547),
.B(n_14),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_427),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_544),
.B(n_208),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_533),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_511),
.B(n_15),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_461),
.B(n_541),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_457),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_548),
.B(n_249),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_443),
.B(n_16),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_541),
.B(n_20),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_548),
.A2(n_247),
.B1(n_215),
.B2(n_209),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_536),
.B(n_257),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_548),
.B(n_185),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_433),
.B(n_24),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_497),
.B(n_257),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_497),
.B(n_257),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_505),
.A2(n_185),
.B1(n_240),
.B2(n_216),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_485),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_476),
.B(n_521),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_467),
.B(n_185),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_433),
.B(n_25),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_520),
.Y(n_649)
);

BUFx12f_ASAP7_75t_SL g650 ( 
.A(n_538),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_543),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_439),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_479),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_494),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_466),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_452),
.B(n_25),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_486),
.B(n_257),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_489),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_536),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g661 ( 
.A1(n_474),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_470),
.B(n_240),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_486),
.B(n_240),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_491),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_493),
.A2(n_500),
.B1(n_519),
.B2(n_538),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_486),
.B(n_240),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_519),
.A2(n_240),
.B1(n_216),
.B2(n_38),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_531),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_458),
.B(n_240),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_531),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_499),
.B(n_506),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_542),
.B(n_33),
.C(n_34),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_431),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_458),
.B(n_240),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_535),
.B(n_507),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_463),
.B(n_216),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_507),
.B(n_517),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_429),
.B(n_216),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_463),
.B(n_38),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_484),
.B(n_40),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_484),
.B(n_44),
.C(n_45),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_546),
.B(n_44),
.Y(n_682)
);

O2A1O1Ixp5_ASAP7_75t_L g683 ( 
.A1(n_546),
.A2(n_45),
.B(n_57),
.C(n_78),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_539),
.B(n_141),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_507),
.B(n_83),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_436),
.B(n_137),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_517),
.B(n_512),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_534),
.B(n_84),
.C(n_108),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_517),
.B(n_512),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_538),
.A2(n_114),
.B1(n_116),
.B2(n_119),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_536),
.B(n_120),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_436),
.B(n_125),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_529),
.A2(n_129),
.B1(n_131),
.B2(n_135),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_536),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_448),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_504),
.B(n_512),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_513),
.B(n_540),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_508),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_590),
.A2(n_529),
.B(n_504),
.C(n_534),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_644),
.B(n_504),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_567),
.A2(n_522),
.B(n_515),
.C(n_509),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_610),
.B(n_492),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_574),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_632),
.B(n_571),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_632),
.B(n_502),
.Y(n_705)
);

NAND2x1_ASAP7_75t_L g706 ( 
.A(n_695),
.B(n_441),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_571),
.B(n_471),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_569),
.B(n_471),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_587),
.B(n_447),
.Y(n_709)
);

BUFx8_ASAP7_75t_SL g710 ( 
.A(n_564),
.Y(n_710)
);

CKINVDCx10_ASAP7_75t_R g711 ( 
.A(n_584),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_677),
.A2(n_689),
.B(n_687),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_578),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_614),
.B(n_498),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_687),
.A2(n_495),
.B(n_528),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_636),
.A2(n_528),
.B1(n_530),
.B2(n_510),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_554),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_636),
.B(n_579),
.C(n_661),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_605),
.B(n_510),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_689),
.A2(n_530),
.B(n_498),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_695),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_651),
.A2(n_473),
.B1(n_498),
.B2(n_466),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_696),
.A2(n_498),
.B(n_473),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_570),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_696),
.A2(n_473),
.B(n_455),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_678),
.A2(n_473),
.B(n_455),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_579),
.A2(n_494),
.B1(n_464),
.B2(n_527),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_609),
.A2(n_518),
.B1(n_464),
.B2(n_527),
.Y(n_728)
);

BUFx4f_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_611),
.A2(n_597),
.B(n_619),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_597),
.A2(n_518),
.B(n_526),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

OR2x6_ASAP7_75t_L g733 ( 
.A(n_647),
.B(n_532),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_600),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_565),
.B(n_526),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_658),
.A2(n_478),
.B(n_532),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_627),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_555),
.Y(n_738)
);

INVx5_ASAP7_75t_L g739 ( 
.A(n_647),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_556),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_663),
.A2(n_478),
.B(n_537),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_666),
.A2(n_478),
.B(n_454),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_631),
.A2(n_591),
.B(n_594),
.C(n_619),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_671),
.A2(n_478),
.B(n_494),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_557),
.A2(n_454),
.B1(n_494),
.B2(n_561),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_612),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_561),
.B(n_454),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_562),
.A2(n_494),
.B(n_563),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_654),
.B(n_551),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_570),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_596),
.B(n_608),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_553),
.B(n_591),
.Y(n_752)
);

INVxp67_ASAP7_75t_SL g753 ( 
.A(n_623),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_592),
.A2(n_633),
.B(n_599),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_593),
.A2(n_616),
.B(n_628),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_673),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_606),
.B(n_649),
.Y(n_757)
);

NOR2x1_ASAP7_75t_L g758 ( 
.A(n_588),
.B(n_584),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_631),
.B(n_614),
.C(n_634),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_667),
.A2(n_594),
.B1(n_623),
.B2(n_613),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_684),
.A2(n_642),
.B(n_641),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_615),
.A2(n_617),
.B1(n_630),
.B2(n_568),
.Y(n_762)
);

AOI21xp33_ASAP7_75t_L g763 ( 
.A1(n_601),
.A2(n_602),
.B(n_629),
.Y(n_763)
);

AO32x1_ASAP7_75t_L g764 ( 
.A1(n_659),
.A2(n_664),
.A3(n_668),
.B1(n_670),
.B2(n_660),
.Y(n_764)
);

NAND2x1_ASAP7_75t_L g765 ( 
.A(n_570),
.B(n_624),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_697),
.B(n_607),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_685),
.A2(n_682),
.B(n_679),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_559),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_573),
.A2(n_576),
.B(n_694),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_573),
.A2(n_576),
.B(n_638),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_638),
.A2(n_577),
.B(n_685),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_552),
.B(n_577),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_680),
.A2(n_657),
.B(n_648),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_552),
.B(n_626),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_580),
.A2(n_603),
.B1(n_575),
.B2(n_566),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_602),
.B(n_582),
.Y(n_776)
);

BUFx4f_ASAP7_75t_L g777 ( 
.A(n_556),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_572),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_589),
.B(n_595),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_586),
.B(n_625),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_640),
.B(n_657),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_640),
.B(n_648),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_683),
.A2(n_665),
.B(n_686),
.Y(n_783)
);

BUFx12f_ASAP7_75t_SL g784 ( 
.A(n_584),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_R g785 ( 
.A(n_655),
.B(n_624),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_570),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_656),
.B(n_622),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_652),
.B(n_604),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_653),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_665),
.A2(n_620),
.B1(n_650),
.B2(n_681),
.Y(n_790)
);

O2A1O1Ixp5_ASAP7_75t_L g791 ( 
.A1(n_621),
.A2(n_646),
.B(n_583),
.C(n_639),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_643),
.A2(n_672),
.B(n_690),
.C(n_637),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_558),
.B(n_618),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_656),
.A2(n_692),
.B(n_691),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_572),
.B(n_656),
.Y(n_795)
);

OAI21xp33_ASAP7_75t_L g796 ( 
.A1(n_635),
.A2(n_643),
.B(n_581),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_656),
.A2(n_674),
.B(n_669),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_676),
.A2(n_690),
.B(n_688),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_572),
.B(n_662),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_693),
.A2(n_655),
.B(n_698),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_655),
.B(n_598),
.Y(n_801)
);

AOI21x1_ASAP7_75t_L g802 ( 
.A1(n_655),
.A2(n_678),
.B(n_522),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_571),
.B(n_437),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_636),
.A2(n_560),
.B1(n_571),
.B2(n_590),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_570),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_647),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_644),
.B(n_284),
.Y(n_808)
);

NOR2x1_ASAP7_75t_L g809 ( 
.A(n_588),
.B(n_453),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_564),
.B(n_438),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_636),
.A2(n_560),
.B1(n_571),
.B2(n_590),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_564),
.B(n_438),
.Y(n_812)
);

OR2x6_ASAP7_75t_SL g813 ( 
.A(n_596),
.B(n_428),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_610),
.B(n_459),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_571),
.B(n_437),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_644),
.B(n_284),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_564),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_610),
.A2(n_611),
.B(n_597),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_686),
.A2(n_692),
.B(n_684),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_644),
.B(n_284),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_636),
.B(n_428),
.C(n_398),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_570),
.Y(n_824)
);

OA22x2_ASAP7_75t_L g825 ( 
.A1(n_596),
.A2(n_483),
.B1(n_608),
.B2(n_549),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_570),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_570),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_554),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_610),
.B(n_459),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_574),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_570),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_574),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_627),
.B(n_437),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_610),
.B(n_459),
.Y(n_835)
);

AOI21x1_ASAP7_75t_L g836 ( 
.A1(n_678),
.A2(n_522),
.B(n_658),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_570),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_574),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_590),
.A2(n_636),
.B(n_691),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_647),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_610),
.A2(n_611),
.B(n_597),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_571),
.B(n_437),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_571),
.B(n_437),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_610),
.A2(n_611),
.B(n_597),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_695),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_644),
.B(n_284),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_574),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_610),
.B(n_459),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_852)
);

BUFx2_ASAP7_75t_SL g853 ( 
.A(n_627),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_610),
.A2(n_645),
.B(n_675),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_574),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_610),
.B(n_459),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_610),
.B(n_459),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_695),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_636),
.A2(n_560),
.B1(n_571),
.B2(n_590),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_610),
.A2(n_611),
.B(n_597),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_686),
.A2(n_692),
.B(n_684),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_816),
.B(n_830),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_835),
.B(n_851),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_805),
.A2(n_811),
.B(n_859),
.C(n_743),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_SL g865 ( 
.A(n_784),
.B(n_807),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_723),
.A2(n_725),
.B(n_720),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_836),
.A2(n_821),
.B(n_861),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_856),
.B(n_857),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_704),
.B(n_766),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_810),
.B(n_812),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_715),
.A2(n_748),
.B(n_741),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_819),
.B(n_757),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_710),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_736),
.A2(n_802),
.B(n_742),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_739),
.B(n_840),
.Y(n_875)
);

OA22x2_ASAP7_75t_L g876 ( 
.A1(n_803),
.A2(n_843),
.B1(n_817),
.B2(n_842),
.Y(n_876)
);

AO31x2_ASAP7_75t_L g877 ( 
.A1(n_760),
.A2(n_846),
.A3(n_847),
.B(n_844),
.Y(n_877)
);

OA21x2_ASAP7_75t_L g878 ( 
.A1(n_783),
.A2(n_730),
.B(n_767),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_853),
.B(n_807),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_852),
.A2(n_854),
.B(n_712),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_798),
.A2(n_699),
.A3(n_792),
.B(n_728),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_808),
.B(n_818),
.Y(n_882)
);

CKINVDCx8_ASAP7_75t_R g883 ( 
.A(n_711),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_730),
.A2(n_860),
.B(n_845),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_820),
.A2(n_860),
.B(n_845),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_820),
.A2(n_841),
.B(n_718),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_841),
.A2(n_773),
.B(n_793),
.C(n_782),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_702),
.B(n_749),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_752),
.B(n_781),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_705),
.B(n_753),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_729),
.B(n_777),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_786),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_703),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_707),
.B(n_713),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_732),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_744),
.A2(n_731),
.B(n_769),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_739),
.B(n_840),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_773),
.A2(n_759),
.B(n_796),
.C(n_767),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_734),
.B(n_746),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_829),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_776),
.A2(n_709),
.B(n_763),
.C(n_722),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_831),
.B(n_833),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_714),
.A2(n_744),
.B(n_770),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_731),
.A2(n_726),
.B(n_755),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_838),
.B(n_850),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_855),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_762),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_708),
.A2(n_754),
.B(n_735),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_717),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_739),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_780),
.B(n_858),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_765),
.A2(n_701),
.B(n_791),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_738),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_727),
.A2(n_716),
.B(n_747),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_789),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_706),
.A2(n_745),
.B(n_788),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_800),
.A2(n_837),
.B(n_750),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_700),
.A2(n_772),
.B(n_801),
.Y(n_918)
);

INVx6_ASAP7_75t_L g919 ( 
.A(n_739),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_822),
.B(n_849),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_786),
.B(n_827),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_774),
.A2(n_775),
.B(n_848),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_721),
.Y(n_923)
);

AOI21xp33_ASAP7_75t_L g924 ( 
.A1(n_825),
.A2(n_823),
.B(n_790),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_764),
.A2(n_795),
.B(n_785),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_826),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_756),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_SL g928 ( 
.A1(n_733),
.A2(n_785),
.B(n_828),
.Y(n_928)
);

NOR2x1_ASAP7_75t_SL g929 ( 
.A(n_733),
.B(n_840),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_799),
.A2(n_824),
.B(n_724),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_764),
.A2(n_719),
.B(n_837),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_832),
.A2(n_758),
.B(n_779),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_733),
.A2(n_825),
.B1(n_840),
.B2(n_778),
.Y(n_933)
);

OAI22x1_ASAP7_75t_L g934 ( 
.A1(n_751),
.A2(n_737),
.B1(n_809),
.B2(n_813),
.Y(n_934)
);

OAI21x1_ASAP7_75t_SL g935 ( 
.A1(n_764),
.A2(n_786),
.B(n_806),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_740),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_806),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_806),
.A2(n_827),
.B(n_828),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_827),
.A2(n_828),
.B(n_834),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_703),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_819),
.B(n_428),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_786),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_768),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_805),
.A2(n_811),
.B1(n_859),
.B2(n_743),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_816),
.B(n_830),
.Y(n_946)
);

OAI21x1_ASAP7_75t_SL g947 ( 
.A1(n_730),
.A2(n_839),
.B(n_841),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_810),
.B(n_427),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_L g950 ( 
.A(n_743),
.B(n_781),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_703),
.Y(n_951)
);

O2A1O1Ixp5_ASAP7_75t_L g952 ( 
.A1(n_730),
.A2(n_743),
.B(n_841),
.C(n_820),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_804),
.A2(n_815),
.B(n_814),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_729),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_768),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_956)
);

AO21x2_ASAP7_75t_L g957 ( 
.A1(n_783),
.A2(n_730),
.B(n_839),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_804),
.A2(n_815),
.B(n_814),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_959)
);

O2A1O1Ixp5_ASAP7_75t_L g960 ( 
.A1(n_730),
.A2(n_743),
.B(n_841),
.C(n_820),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_805),
.A2(n_859),
.B(n_811),
.C(n_743),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_962)
);

AOI221xp5_ASAP7_75t_L g963 ( 
.A1(n_718),
.A2(n_661),
.B1(n_811),
.B2(n_859),
.C(n_805),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_810),
.B(n_812),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_794),
.A2(n_771),
.B(n_761),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_819),
.B(n_428),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_816),
.B(n_830),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_819),
.B(n_428),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_739),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_804),
.A2(n_815),
.B(n_814),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_810),
.B(n_812),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_739),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_810),
.B(n_812),
.Y(n_975)
);

OAI22x1_ASAP7_75t_L g976 ( 
.A1(n_805),
.A2(n_859),
.B1(n_811),
.B2(n_483),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_805),
.B(n_811),
.Y(n_977)
);

AO21x2_ASAP7_75t_L g978 ( 
.A1(n_783),
.A2(n_730),
.B(n_839),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_794),
.A2(n_787),
.B(n_797),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_928),
.B(n_875),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_927),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_889),
.B(n_869),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_870),
.B(n_964),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_889),
.B(n_869),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_875),
.B(n_897),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_862),
.B(n_863),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_899),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_890),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_899),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_897),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_862),
.B(n_863),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_879),
.B(n_954),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_883),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_902),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_972),
.Y(n_995)
);

AND2x2_ASAP7_75t_SL g996 ( 
.A(n_963),
.B(n_865),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_902),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_975),
.B(n_872),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_868),
.B(n_946),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_868),
.B(n_946),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_905),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_967),
.B(n_888),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_910),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_967),
.B(n_888),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_882),
.B(n_920),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_948),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_887),
.B(n_977),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_900),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_953),
.A2(n_971),
.B(n_958),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_905),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_942),
.B(n_966),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_963),
.B(n_968),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_909),
.B(n_895),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_906),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_976),
.B(n_944),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_893),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_910),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_955),
.B(n_936),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_941),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_879),
.B(n_929),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_921),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_L g1022 ( 
.A(n_934),
.B(n_892),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_864),
.A2(n_961),
.B(n_898),
.C(n_945),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_873),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_951),
.B(n_915),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_910),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_891),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_923),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_924),
.B(n_911),
.Y(n_1029)
);

NOR2xp67_ASAP7_75t_L g1030 ( 
.A(n_892),
.B(n_943),
.Y(n_1030)
);

BUFx4_ASAP7_75t_SL g1031 ( 
.A(n_937),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_945),
.A2(n_884),
.B1(n_885),
.B2(n_886),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_970),
.Y(n_1033)
);

HAxp5_ASAP7_75t_L g1034 ( 
.A(n_952),
.B(n_960),
.CON(n_1034),
.SN(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_886),
.B(n_884),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_921),
.Y(n_1036)
);

CKINVDCx14_ASAP7_75t_R g1037 ( 
.A(n_921),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_924),
.B(n_911),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_926),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_913),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_890),
.B(n_907),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_921),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_974),
.Y(n_1043)
);

INVx4_ASAP7_75t_SL g1044 ( 
.A(n_921),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_933),
.B(n_943),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_876),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_974),
.B(n_932),
.Y(n_1047)
);

AND2x6_ASAP7_75t_L g1048 ( 
.A(n_894),
.B(n_876),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_922),
.B(n_933),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_922),
.B(n_878),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_947),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_919),
.B(n_939),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_878),
.B(n_957),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_901),
.A2(n_916),
.B(n_931),
.C(n_925),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_930),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_930),
.B(n_938),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_957),
.B(n_978),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_978),
.B(n_877),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_918),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_914),
.A2(n_903),
.B1(n_908),
.B2(n_935),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_917),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_914),
.A2(n_896),
.B(n_925),
.Y(n_1062)
);

AND2x4_ASAP7_75t_SL g1063 ( 
.A(n_912),
.B(n_881),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_874),
.B(n_904),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_965),
.A2(n_871),
.B1(n_866),
.B2(n_867),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_940),
.B(n_949),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_956),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_959),
.B(n_962),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_979),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_969),
.B(n_973),
.Y(n_1070)
);

AOI21xp33_ASAP7_75t_SL g1071 ( 
.A1(n_942),
.A2(n_428),
.B(n_422),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_899),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_880),
.A2(n_814),
.B(n_804),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_882),
.B(n_428),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_883),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_927),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_899),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_910),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_883),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_870),
.B(n_964),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_950),
.A2(n_814),
.B(n_804),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_945),
.A2(n_743),
.B(n_884),
.C(n_952),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_889),
.B(n_869),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_889),
.B(n_869),
.Y(n_1084)
);

INVx3_ASAP7_75t_SL g1085 ( 
.A(n_873),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_945),
.B(n_784),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_899),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_875),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_864),
.A2(n_961),
.B1(n_945),
.B2(n_887),
.Y(n_1089)
);

BUFx2_ASAP7_75t_SL g1090 ( 
.A(n_883),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_882),
.A2(n_421),
.B1(n_811),
.B2(n_805),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_879),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_899),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1036),
.Y(n_1094)
);

BUFx2_ASAP7_75t_SL g1095 ( 
.A(n_1075),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1026),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1034),
.B(n_1057),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1013),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1025),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1032),
.B(n_1035),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1032),
.B(n_1035),
.Y(n_1101)
);

BUFx2_ASAP7_75t_R g1102 ( 
.A(n_1090),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_996),
.A2(n_1012),
.B1(n_1091),
.B2(n_1029),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1044),
.B(n_980),
.Y(n_1104)
);

OR2x6_ASAP7_75t_L g1105 ( 
.A(n_980),
.B(n_1049),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1019),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_995),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1014),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1016),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1005),
.B(n_986),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_981),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1044),
.B(n_980),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1048),
.A2(n_1086),
.B1(n_1089),
.B2(n_1038),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_1020),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1050),
.B(n_1053),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1086),
.A2(n_1074),
.B1(n_1011),
.B2(n_983),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1040),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_SL g1118 ( 
.A1(n_1048),
.A2(n_1089),
.B1(n_1046),
.B2(n_1037),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1015),
.B(n_1023),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1044),
.B(n_985),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1007),
.A2(n_999),
.B1(n_991),
.B2(n_1000),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_1018),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_981),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1080),
.A2(n_982),
.B1(n_984),
.B2(n_1084),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1048),
.A2(n_1007),
.B1(n_1045),
.B2(n_988),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_998),
.B(n_1076),
.Y(n_1126)
);

INVx11_ASAP7_75t_L g1127 ( 
.A(n_1048),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1028),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1039),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1002),
.A2(n_1004),
.B1(n_984),
.B2(n_1084),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_993),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_987),
.Y(n_1132)
);

INVx11_ASAP7_75t_L g1133 ( 
.A(n_1031),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_1079),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_982),
.A2(n_1083),
.B1(n_1076),
.B2(n_986),
.Y(n_1135)
);

AO21x1_ASAP7_75t_SL g1136 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1051),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1002),
.A2(n_1004),
.B1(n_1083),
.B2(n_1000),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1021),
.B(n_1042),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_989),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_991),
.B(n_999),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_994),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1056),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1093),
.A2(n_997),
.B1(n_1072),
.B2(n_1077),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1001),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1010),
.B(n_1087),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1056),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1006),
.A2(n_1008),
.B1(n_1071),
.B2(n_1022),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_1085),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1055),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_1003),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1043),
.B(n_1027),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_SL g1153 ( 
.A1(n_1092),
.A2(n_1009),
.B(n_1081),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1059),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1003),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1082),
.B(n_1060),
.Y(n_1156)
);

CKINVDCx11_ASAP7_75t_R g1157 ( 
.A(n_992),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1024),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1047),
.B(n_1063),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1020),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_990),
.B(n_1088),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1003),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1017),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1017),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1017),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1062),
.A2(n_1054),
.B(n_1073),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1078),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1062),
.A2(n_1066),
.B(n_1070),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1078),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1088),
.B(n_1033),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1030),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1052),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1069),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1061),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1065),
.A2(n_1064),
.B(n_1066),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_1067),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1068),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1013),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1034),
.B(n_1057),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1013),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1025),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1005),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1025),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1005),
.A2(n_1012),
.B1(n_1091),
.B2(n_805),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_996),
.A2(n_976),
.B1(n_977),
.B2(n_718),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_996),
.A2(n_284),
.B1(n_305),
.B2(n_304),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1097),
.B(n_1179),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1150),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1173),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1097),
.B(n_1179),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1100),
.B(n_1101),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1184),
.A2(n_1185),
.B(n_1103),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1100),
.B(n_1101),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_1153),
.A2(n_1166),
.B(n_1154),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1176),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1121),
.B(n_1130),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1119),
.A2(n_1156),
.B1(n_1103),
.B2(n_1112),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1111),
.Y(n_1198)
);

CKINVDCx6p67_ASAP7_75t_R g1199 ( 
.A(n_1096),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1115),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1115),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1174),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1123),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1176),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1174),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1142),
.B(n_1147),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1131),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1137),
.B(n_1135),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1104),
.B(n_1112),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1132),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1139),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1107),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1106),
.Y(n_1213)
);

AO21x2_ASAP7_75t_L g1214 ( 
.A1(n_1166),
.A2(n_1175),
.B(n_1146),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1128),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1141),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1129),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1144),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1168),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1109),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1117),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1142),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1147),
.B(n_1119),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1147),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1145),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1098),
.B(n_1178),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1145),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1136),
.B(n_1099),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1177),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1181),
.B(n_1183),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1108),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1172),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1159),
.B(n_1124),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1113),
.A2(n_1143),
.B(n_1185),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1105),
.Y(n_1235)
);

INVx4_ASAP7_75t_SL g1236 ( 
.A(n_1105),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1096),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1143),
.Y(n_1238)
);

AND2x4_ASAP7_75t_SL g1239 ( 
.A(n_1104),
.B(n_1112),
.Y(n_1239)
);

AOI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1125),
.A2(n_1118),
.B(n_1110),
.Y(n_1240)
);

INVxp67_ASAP7_75t_R g1241 ( 
.A(n_1170),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1180),
.B(n_1140),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1131),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1126),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1160),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1189),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1191),
.B(n_1122),
.Y(n_1247)
);

NOR2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1196),
.B(n_1094),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1189),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1191),
.B(n_1193),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1219),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1192),
.B(n_1116),
.C(n_1182),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1194),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1193),
.B(n_1170),
.Y(n_1254)
);

OAI211xp5_ASAP7_75t_L g1255 ( 
.A1(n_1192),
.A2(n_1186),
.B(n_1157),
.C(n_1152),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1187),
.B(n_1114),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1187),
.B(n_1190),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1190),
.B(n_1114),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1226),
.B(n_1138),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1223),
.B(n_1164),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1223),
.B(n_1165),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1206),
.B(n_1163),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1226),
.B(n_1167),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1204),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1225),
.B(n_1162),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1234),
.A2(n_1157),
.B1(n_1120),
.B2(n_1134),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1236),
.B(n_1224),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1227),
.B(n_1169),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1214),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1196),
.B(n_1148),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1203),
.B(n_1171),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1194),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1214),
.B(n_1161),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1214),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1214),
.B(n_1151),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1203),
.B(n_1155),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1222),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1234),
.A2(n_1120),
.B1(n_1134),
.B2(n_1095),
.Y(n_1279)
);

OAI221xp5_ASAP7_75t_L g1280 ( 
.A1(n_1271),
.A2(n_1252),
.B1(n_1208),
.B2(n_1255),
.C(n_1240),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1257),
.B(n_1250),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1257),
.B(n_1228),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1257),
.B(n_1228),
.Y(n_1283)
);

NAND4xp25_ASAP7_75t_L g1284 ( 
.A(n_1252),
.B(n_1212),
.C(n_1208),
.D(n_1240),
.Y(n_1284)
);

NAND4xp25_ASAP7_75t_L g1285 ( 
.A(n_1252),
.B(n_1229),
.C(n_1197),
.D(n_1220),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1271),
.A2(n_1234),
.B1(n_1238),
.B2(n_1233),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1246),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1250),
.B(n_1241),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1254),
.B(n_1241),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1270),
.B(n_1188),
.C(n_1229),
.Y(n_1290)
);

NOR3xp33_ASAP7_75t_SL g1291 ( 
.A(n_1255),
.B(n_1158),
.C(n_1133),
.Y(n_1291)
);

NAND4xp25_ASAP7_75t_L g1292 ( 
.A(n_1278),
.B(n_1221),
.C(n_1220),
.D(n_1195),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1246),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_L g1294 ( 
.A(n_1270),
.B(n_1213),
.C(n_1215),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1265),
.B(n_1204),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1254),
.B(n_1198),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_1270),
.B(n_1273),
.C(n_1253),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1253),
.B(n_1217),
.C(n_1222),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1248),
.B(n_1274),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1267),
.A2(n_1195),
.B(n_1233),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1267),
.A2(n_1234),
.B1(n_1238),
.B2(n_1235),
.Y(n_1301)
);

AOI221x1_ASAP7_75t_SL g1302 ( 
.A1(n_1272),
.A2(n_1221),
.B1(n_1211),
.B2(n_1218),
.C(n_1216),
.Y(n_1302)
);

NAND3xp33_ASAP7_75t_L g1303 ( 
.A(n_1273),
.B(n_1210),
.C(n_1211),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1272),
.B(n_1242),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1247),
.B(n_1242),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1275),
.B(n_1216),
.C(n_1218),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1247),
.B(n_1158),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1247),
.B(n_1149),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1260),
.B(n_1224),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1279),
.A2(n_1239),
.B(n_1209),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1277),
.B(n_1244),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1277),
.B(n_1230),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1266),
.A2(n_1230),
.B(n_1231),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1248),
.A2(n_1127),
.B1(n_1237),
.B2(n_1199),
.Y(n_1314)
);

AND4x1_ASAP7_75t_L g1315 ( 
.A(n_1276),
.B(n_1133),
.C(n_1237),
.D(n_1199),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1260),
.B(n_1194),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1266),
.B(n_1200),
.Y(n_1317)
);

AND2x2_ASAP7_75t_SL g1318 ( 
.A(n_1268),
.B(n_1239),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1275),
.A2(n_1231),
.B1(n_1201),
.B2(n_1232),
.C(n_1245),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1261),
.B(n_1194),
.Y(n_1320)
);

NAND4xp25_ASAP7_75t_L g1321 ( 
.A(n_1278),
.B(n_1204),
.C(n_1202),
.D(n_1205),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1269),
.B(n_1201),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1287),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1287),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1293),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1293),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1311),
.B(n_1263),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1304),
.B(n_1263),
.Y(n_1328)
);

INVxp33_ASAP7_75t_L g1329 ( 
.A(n_1308),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1305),
.B(n_1263),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1302),
.B(n_1246),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1299),
.B(n_1251),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1316),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1318),
.B(n_1265),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1309),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1303),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1281),
.B(n_1264),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1299),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1313),
.B(n_1319),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1313),
.B(n_1249),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1306),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1299),
.B(n_1258),
.Y(n_1346)
);

AND2x2_ASAP7_75t_SL g1347 ( 
.A(n_1318),
.B(n_1239),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1289),
.B(n_1248),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1317),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1312),
.B(n_1259),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1294),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1296),
.B(n_1259),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1322),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1338),
.B(n_1290),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1341),
.B(n_1292),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1331),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1331),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1323),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1323),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1325),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1324),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1342),
.B(n_1288),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1332),
.B(n_1340),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1338),
.B(n_1256),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_L g1365 ( 
.A(n_1345),
.B(n_1321),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1325),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1342),
.B(n_1289),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1326),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1345),
.B(n_1256),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1342),
.B(n_1307),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1344),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1347),
.B(n_1315),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1326),
.Y(n_1373)
);

NAND4xp25_ASAP7_75t_L g1374 ( 
.A(n_1341),
.B(n_1284),
.C(n_1280),
.D(n_1298),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1351),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1324),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1324),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1332),
.B(n_1315),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1344),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1351),
.B(n_1269),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1343),
.B(n_1295),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1337),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1349),
.B(n_1261),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1334),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1334),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1327),
.Y(n_1386)
);

OR2x6_ASAP7_75t_L g1387 ( 
.A(n_1336),
.B(n_1310),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1349),
.B(n_1261),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1346),
.B(n_1262),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1356),
.B(n_1339),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1378),
.B(n_1346),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1354),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1359),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1389),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1386),
.B(n_1327),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1364),
.B(n_1369),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1359),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1357),
.B(n_1339),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1378),
.B(n_1346),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1374),
.B(n_1329),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1360),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1355),
.B(n_1328),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1375),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1360),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1366),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1355),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1379),
.B(n_1371),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1378),
.B(n_1348),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1379),
.B(n_1384),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1372),
.B(n_1207),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1384),
.B(n_1339),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1366),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1368),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1370),
.B(n_1348),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1365),
.B(n_1347),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1380),
.B(n_1328),
.Y(n_1416)
);

OAI21xp33_ASAP7_75t_L g1417 ( 
.A1(n_1385),
.A2(n_1335),
.B(n_1340),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1387),
.A2(n_1300),
.B(n_1297),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1383),
.B(n_1388),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1385),
.B(n_1358),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_1363),
.B(n_1332),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1363),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1370),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1381),
.B(n_1207),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1368),
.B(n_1353),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1373),
.Y(n_1426)
);

NOR3x1_ASAP7_75t_L g1427 ( 
.A(n_1372),
.B(n_1314),
.C(n_1285),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1373),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1363),
.B(n_1332),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1376),
.Y(n_1430)
);

OAI33xp33_ASAP7_75t_L g1431 ( 
.A1(n_1376),
.A2(n_1335),
.A3(n_1353),
.B1(n_1352),
.B2(n_1350),
.B3(n_1330),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1415),
.B(n_1362),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1403),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1393),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1392),
.B(n_1207),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1400),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1406),
.B(n_1361),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1397),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1415),
.B(n_1362),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1401),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1390),
.B(n_1361),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1410),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1418),
.A2(n_1286),
.B1(n_1301),
.B2(n_1387),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1402),
.B(n_1382),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1390),
.B(n_1377),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1404),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1414),
.B(n_1367),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1410),
.Y(n_1448)
);

NAND3xp33_ASAP7_75t_L g1449 ( 
.A(n_1407),
.B(n_1409),
.C(n_1398),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1405),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1391),
.B(n_1367),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1399),
.B(n_1387),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1412),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1398),
.B(n_1377),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1421),
.B(n_1372),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1423),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1424),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1395),
.B(n_1382),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1422),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1413),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1422),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1408),
.B(n_1429),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1426),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1428),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1420),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1431),
.A2(n_1387),
.B1(n_1274),
.B2(n_1333),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1438),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1456),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1447),
.B(n_1394),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1438),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1433),
.B(n_1436),
.Y(n_1471)
);

AOI21xp33_ASAP7_75t_L g1472 ( 
.A1(n_1436),
.A2(n_1407),
.B(n_1409),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1452),
.A2(n_1411),
.B(n_1410),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1443),
.A2(n_1417),
.B1(n_1430),
.B2(n_1396),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1452),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1449),
.A2(n_1466),
.B(n_1437),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1447),
.B(n_1416),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1442),
.B(n_1347),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1446),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1442),
.Y(n_1481)
);

BUFx2_ASAP7_75t_SL g1482 ( 
.A(n_1442),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1464),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1464),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1464),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1448),
.A2(n_1427),
.B1(n_1420),
.B2(n_1425),
.C(n_1411),
.Y(n_1486)
);

AOI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1448),
.A2(n_1425),
.B(n_1419),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1434),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1437),
.B(n_1330),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1434),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1440),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1468),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1483),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1471),
.B(n_1449),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1478),
.B(n_1465),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1484),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1478),
.B(n_1465),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1485),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1481),
.B(n_1451),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1467),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1476),
.B(n_1451),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1482),
.B(n_1457),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1482),
.B(n_1462),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1469),
.B(n_1462),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_SL g1505 ( 
.A(n_1486),
.B(n_1439),
.C(n_1432),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1470),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1480),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1467),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1469),
.B(n_1432),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1489),
.B(n_1458),
.Y(n_1510)
);

AOI211xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1502),
.A2(n_1472),
.B(n_1487),
.C(n_1473),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1502),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1503),
.B(n_1474),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1494),
.A2(n_1475),
.B1(n_1479),
.B2(n_1477),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1494),
.B(n_1457),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1492),
.B(n_1473),
.C(n_1461),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1503),
.B(n_1448),
.Y(n_1517)
);

OAI211xp5_ASAP7_75t_L g1518 ( 
.A1(n_1505),
.A2(n_1491),
.B(n_1488),
.C(n_1490),
.Y(n_1518)
);

NOR3xp33_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1435),
.C(n_1479),
.Y(n_1519)
);

NAND4xp25_ASAP7_75t_SL g1520 ( 
.A(n_1509),
.B(n_1439),
.C(n_1461),
.D(n_1459),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1509),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1510),
.A2(n_1444),
.B1(n_1489),
.B2(n_1458),
.Y(n_1522)
);

AND3x1_ASAP7_75t_L g1523 ( 
.A(n_1511),
.B(n_1508),
.C(n_1500),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1515),
.B(n_1504),
.Y(n_1524)
);

NOR3xp33_ASAP7_75t_L g1525 ( 
.A(n_1512),
.B(n_1510),
.C(n_1497),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1521),
.B(n_1504),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1516),
.Y(n_1527)
);

NOR3x1_ASAP7_75t_L g1528 ( 
.A(n_1513),
.B(n_1501),
.C(n_1495),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1522),
.Y(n_1529)
);

NAND3xp33_ASAP7_75t_SL g1530 ( 
.A(n_1514),
.B(n_1507),
.C(n_1506),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1517),
.B(n_1493),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1520),
.B(n_1496),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1524),
.Y(n_1533)
);

AOI221x1_ASAP7_75t_L g1534 ( 
.A1(n_1530),
.A2(n_1519),
.B1(n_1498),
.B2(n_1461),
.C(n_1459),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1523),
.A2(n_1455),
.B1(n_1518),
.B2(n_1459),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1525),
.B(n_1149),
.C(n_1444),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1527),
.A2(n_1243),
.B1(n_1460),
.B2(n_1453),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1533),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1534),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1535),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1536),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1537),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1536),
.A2(n_1523),
.B1(n_1529),
.B2(n_1532),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1538),
.B(n_1526),
.Y(n_1544)
);

AOI211xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1539),
.A2(n_1531),
.B(n_1528),
.C(n_1453),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1541),
.B(n_1463),
.Y(n_1546)
);

NOR2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1540),
.B(n_1243),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1541),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1548),
.B(n_1543),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1547),
.Y(n_1550)
);

AND4x1_ASAP7_75t_L g1551 ( 
.A(n_1544),
.B(n_1542),
.C(n_1291),
.D(n_1102),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1549),
.B(n_1546),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1552),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1553),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1553),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1555),
.A2(n_1545),
.B(n_1554),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1555),
.A2(n_1550),
.B(n_1551),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1556),
.A2(n_1243),
.B1(n_1460),
.B2(n_1450),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1557),
.A2(n_1450),
.B(n_1440),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1559),
.B(n_1558),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1560),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_R g1562 ( 
.A1(n_1561),
.A2(n_1463),
.B1(n_1454),
.B2(n_1445),
.C(n_1441),
.Y(n_1562)
);

AOI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1562),
.A2(n_1441),
.B(n_1454),
.C(n_1445),
.Y(n_1563)
);


endmodule