module fake_netlist_6_1194_n_386 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_116, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_386);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_386;

wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_350;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_122;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_352;
wire n_374;
wire n_366;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_265;
wire n_260;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_277;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_364;
wire n_295;
wire n_385;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

BUFx3_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_30),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_18),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_48),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_38),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_51),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_23),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_31),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_27),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_57),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_6),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_39),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

INVxp33_ASAP7_75t_SL g151 ( 
.A(n_64),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_72),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_16),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_33),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_52),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_81),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_8),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_22),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_34),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_0),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_56),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_37),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_118),
.A2(n_130),
.B(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_0),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_58),
.B(n_115),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_126),
.B(n_54),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

OAI22x1_ASAP7_75t_R g191 ( 
.A1(n_127),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_135),
.A2(n_4),
.B(n_5),
.Y(n_192)
);

AND2x2_ASAP7_75t_R g193 ( 
.A(n_139),
.B(n_7),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_138),
.B(n_116),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_131),
.B(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_134),
.B(n_10),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_159),
.Y(n_201)
);

OR2x6_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_148),
.Y(n_202)
);

OR2x6_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_148),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_151),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_R g206 ( 
.A(n_192),
.B(n_119),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_164),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

OR2x6_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_193),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_184),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_161),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_121),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

AO221x1_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_189),
.B1(n_193),
.B2(n_126),
.C(n_157),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_137),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_124),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_132),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_220),
.B(n_141),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_203),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_144),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_147),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_150),
.Y(n_248)
);

NAND2x1_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_184),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_169),
.B1(n_170),
.B2(n_175),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_152),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_158),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_206),
.B(n_160),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_142),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_202),
.A2(n_163),
.B1(n_145),
.B2(n_146),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_162),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_166),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_165),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_228),
.B(n_172),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_183),
.B(n_156),
.Y(n_264)
);

CKINVDCx6p67_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_168),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_155),
.B(n_153),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_143),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_230),
.B(n_176),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_202),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_11),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_191),
.B1(n_13),
.B2(n_14),
.Y(n_275)
);

NAND2x1_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_12),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_19),
.B(n_20),
.Y(n_278)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_21),
.B(n_24),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_25),
.Y(n_280)
);

BUFx8_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

OR2x2_ASAP7_75t_SL g283 ( 
.A(n_258),
.B(n_251),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_32),
.B(n_35),
.C(n_40),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_241),
.B(n_41),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

INVx3_ASAP7_75t_SL g289 ( 
.A(n_265),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

BUFx8_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

AO31x2_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_250),
.A3(n_252),
.B(n_238),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_281),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_246),
.B1(n_234),
.B2(n_251),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_249),
.B(n_256),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_259),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_42),
.B(n_44),
.C(n_47),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_268),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_49),
.B(n_50),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_266),
.A2(n_53),
.B(n_59),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_60),
.B(n_62),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_67),
.B(n_68),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_71),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_73),
.C(n_75),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_SL g309 ( 
.A(n_284),
.B(n_79),
.C(n_80),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_308),
.B1(n_295),
.B2(n_290),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_281),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

NAND2x1p5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_282),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_271),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_283),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_302),
.B(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_291),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_316),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_297),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_299),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_322),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_320),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx5_ASAP7_75t_SL g336 ( 
.A(n_329),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_317),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_329),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_279),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_329),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_334),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_330),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_342),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_330),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_332),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_332),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_324),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_324),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_345),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_342),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_344),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_340),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_356),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_353),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_362),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

NAND4xp25_ASAP7_75t_L g367 ( 
.A(n_365),
.B(n_315),
.C(n_349),
.D(n_354),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_367),
.Y(n_369)
);

AOI211xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_364),
.B(n_363),
.C(n_306),
.Y(n_370)
);

O2A1O1Ixp5_ASAP7_75t_L g371 ( 
.A1(n_368),
.A2(n_359),
.B(n_360),
.C(n_355),
.Y(n_371)
);

NAND4xp25_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_352),
.C(n_350),
.D(n_358),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_R g373 ( 
.A1(n_371),
.A2(n_291),
.B1(n_285),
.B2(n_305),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_374),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_351),
.B1(n_373),
.B2(n_324),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_376),
.A2(n_351),
.B1(n_313),
.B2(n_276),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_378),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_377),
.Y(n_380)
);

AOI221xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_278),
.B1(n_280),
.B2(n_91),
.C(n_93),
.Y(n_381)
);

OAI221xp5_ASAP7_75t_L g382 ( 
.A1(n_379),
.A2(n_82),
.B1(n_88),
.B2(n_94),
.C(n_96),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_382),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_97),
.B(n_100),
.Y(n_384)
);

AO21x2_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_101),
.B(n_102),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_383),
.B1(n_105),
.B2(n_113),
.Y(n_386)
);


endmodule