module fake_jpeg_3864_n_310 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_40),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_23),
.B1(n_39),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_89),
.B1(n_90),
.B2(n_15),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_53),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_54),
.A2(n_63),
.B1(n_69),
.B2(n_72),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_67),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_62),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_23),
.B(n_7),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_15),
.B1(n_26),
.B2(n_20),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_65),
.B1(n_68),
.B2(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_29),
.B1(n_18),
.B2(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_18),
.B1(n_28),
.B2(n_19),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_78),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_37),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_13),
.B1(n_27),
.B2(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_84),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_25),
.B1(n_13),
.B2(n_14),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_91),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_39),
.A2(n_15),
.B1(n_17),
.B2(n_20),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_39),
.A2(n_15),
.B1(n_17),
.B2(n_20),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_96),
.Y(n_121)
);

INVxp67_ASAP7_75t_R g93 ( 
.A(n_36),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_97),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_20),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_99),
.A2(n_116),
.B1(n_118),
.B2(n_60),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_17),
.B1(n_12),
.B2(n_11),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_17),
.B1(n_10),
.B2(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_0),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_69),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_93),
.B(n_54),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_154),
.B(n_119),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_129),
.B(n_132),
.Y(n_193)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_131),
.Y(n_175)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_54),
.B1(n_97),
.B2(n_86),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_65),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_107),
.C(n_101),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_58),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_72),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_148),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_73),
.Y(n_147)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_59),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_63),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_83),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_86),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_51),
.B(n_90),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_75),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_98),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_7),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_89),
.B1(n_74),
.B2(n_60),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_123),
.B1(n_105),
.B2(n_104),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_108),
.B(n_74),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_159),
.B1(n_104),
.B2(n_122),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_98),
.B(n_82),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_167),
.C(n_177),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_101),
.C(n_115),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_107),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_195),
.B(n_130),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_107),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_49),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_180),
.C(n_181),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_115),
.C(n_49),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_49),
.C(n_114),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_105),
.B1(n_123),
.B2(n_114),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_122),
.C(n_119),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_187),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_132),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_145),
.B1(n_151),
.B2(n_138),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_191),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_201),
.B(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_167),
.C(n_181),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_207),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_144),
.B1(n_133),
.B2(n_142),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_223),
.B1(n_224),
.B2(n_188),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_192),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_210),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_139),
.B(n_137),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_180),
.B(n_184),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_162),
.A3(n_161),
.B1(n_134),
.B2(n_131),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_165),
.B(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_2),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

NAND4xp25_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_94),
.C(n_59),
.D(n_52),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_120),
.B1(n_146),
.B2(n_160),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_160),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_173),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_203),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_195),
.B(n_173),
.C(n_178),
.D(n_164),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_205),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_236),
.C(n_243),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_174),
.B1(n_168),
.B2(n_172),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_217),
.B(n_218),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_193),
.C(n_171),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_196),
.C(n_185),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_210),
.C(n_208),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g246 ( 
.A(n_211),
.B(n_198),
.C(n_185),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_252),
.C(n_259),
.Y(n_268)
);

AO221x1_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_221),
.B1(n_197),
.B2(n_213),
.C(n_179),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_207),
.C(n_206),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_204),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_228),
.B(n_231),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_215),
.B(n_201),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_245),
.B1(n_228),
.B2(n_232),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_226),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_203),
.C(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_223),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_276),
.B(n_270),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_246),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_267),
.B(n_234),
.C(n_229),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_256),
.B1(n_258),
.B2(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_243),
.C(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_247),
.C(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_237),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.C(n_285),
.Y(n_288)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_262),
.C(n_251),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_265),
.B(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_268),
.C(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_284),
.B(n_286),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_259),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_271),
.B1(n_264),
.B2(n_275),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_166),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_293),
.B(n_281),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_265),
.A3(n_268),
.B1(n_219),
.B2(n_237),
.C1(n_216),
.C2(n_239),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_294),
.C(n_277),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_292),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_238),
.B(n_176),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_238),
.A3(n_186),
.B1(n_179),
.B2(n_146),
.C1(n_94),
.C2(n_52),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_299),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_288),
.B(n_179),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_186),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_294),
.B(n_291),
.Y(n_304)
);

AOI221xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_2),
.C(n_3),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_298),
.B1(n_7),
.B2(n_4),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_2),
.B(n_3),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_3),
.Y(n_310)
);


endmodule