module fake_netlist_1_10377_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g10 ( .A(n_2), .B(n_4), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_15), .B(n_14), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_12), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_16), .B(n_13), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_18), .B(n_13), .Y(n_21) );
NAND3xp33_ASAP7_75t_L g22 ( .A(n_19), .B(n_10), .C(n_11), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_20), .B(n_17), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
OAI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_17), .B1(n_22), .B2(n_19), .C(n_21), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
NAND5xp2_ASAP7_75t_L g30 ( .A(n_28), .B(n_12), .C(n_1), .D(n_2), .E(n_3), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_27), .B(n_21), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_19), .Y(n_32) );
OAI22x1_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_0), .B1(n_4), .B2(n_5), .Y(n_33) );
OR2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_5), .Y(n_34) );
AOI22xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_19), .B1(n_7), .B2(n_8), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
NAND3xp33_ASAP7_75t_L g38 ( .A(n_37), .B(n_35), .C(n_34), .Y(n_38) );
endmodule