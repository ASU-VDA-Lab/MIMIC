module real_jpeg_23854_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_1),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_79),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_53),
.C(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_31),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_82),
.B1(n_161),
.B2(n_168),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_36),
.B1(n_92),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_8),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_74),
.Y(n_84)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_10),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_70),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_57),
.Y(n_118)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_86),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_19),
.B(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_75),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_20),
.A2(n_21),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_41),
.C(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_23),
.A2(n_37),
.B1(n_39),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_24),
.A2(n_31),
.B1(n_35),
.B2(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_32),
.Y(n_80)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_27),
.A2(n_30),
.A3(n_33),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_28),
.B(n_79),
.CON(n_78),
.SN(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_28),
.A2(n_45),
.B(n_90),
.C(n_93),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_44),
.C(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_32),
.A2(n_33),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_33),
.B(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_44),
.A2(n_45),
.B1(n_91),
.B2(n_92),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_55),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_58),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_50),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_53),
.B1(n_65),
.B2(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_52),
.B(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_60),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_71),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_73),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_63),
.A2(n_69),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_63),
.A2(n_131),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_63),
.A2(n_130),
.B1(n_131),
.B2(n_141),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_68),
.B(n_79),
.Y(n_166)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_77),
.B(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_79),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_82),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_82),
.A2(n_158),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_84),
.B(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_102),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_111),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_135),
.B(n_184),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_126),
.B(n_132),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.C(n_129),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_179),
.B(n_183),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_154),
.B(n_178),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_138),
.B(n_144),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_164),
.B(n_177),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_163),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_171),
.B(n_176),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);


endmodule