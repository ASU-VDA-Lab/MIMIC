module fake_jpeg_12305_n_63 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_20),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_22),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_9),
.B1(n_10),
.B2(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

OA22x2_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_16),
.B1(n_9),
.B2(n_17),
.Y(n_27)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_13),
.B1(n_21),
.B2(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_15),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_13),
.B(n_1),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_25),
.C(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_24),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_37),
.C(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_3),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_42),
.B1(n_38),
.B2(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_0),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_53),
.B1(n_6),
.B2(n_8),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_50),
.C(n_46),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_57),
.C(n_51),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_50),
.B(n_4),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_52),
.B(n_54),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_3),
.B1(n_8),
.B2(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_3),
.Y(n_63)
);


endmodule