module fake_netlist_1_256_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
BUFx6f_ASAP7_75t_SL g3 ( .A(n_2), .Y(n_3) );
AND3x2_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .C(n_1), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
NAND3xp33_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .C(n_1), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
NAND2x1p5_ASAP7_75t_L g8 ( .A(n_3), .B(n_2), .Y(n_8) );
AOI22xp33_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_3), .B1(n_4), .B2(n_2), .Y(n_9) );
BUFx3_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVxp67_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
NAND2x1p5_ASAP7_75t_L g12 ( .A(n_10), .B(n_7), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_10), .B1(n_9), .B2(n_6), .C(n_2), .Y(n_13) );
AOI22xp33_ASAP7_75t_SL g14 ( .A1(n_12), .A2(n_10), .B1(n_9), .B2(n_2), .Y(n_14) );
NAND5xp2_ASAP7_75t_L g15 ( .A(n_14), .B(n_0), .C(n_1), .D(n_12), .E(n_13), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_12), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_0), .B(n_1), .Y(n_17) );
OAI21xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_15), .B(n_1), .Y(n_18) );
endmodule