module fake_netlist_5_1925_n_2369 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_510, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_2369);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2369;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_1547;
wire n_1070;
wire n_777;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_1319;
wire n_561;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_514;
wire n_1079;
wire n_2093;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2340;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_703;
wire n_980;
wire n_1115;
wire n_698;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_2104;
wire n_518;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_517;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_542;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2268;

INVx2_ASAP7_75t_L g513 ( 
.A(n_509),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_174),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_411),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_80),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_52),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_317),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_79),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_448),
.Y(n_521)
);

BUFx5_ASAP7_75t_L g522 ( 
.A(n_187),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_20),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_58),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_63),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_484),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_227),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_43),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_198),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_405),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_452),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_427),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_213),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_507),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_453),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_390),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_126),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_59),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_261),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_72),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_0),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_419),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_60),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_89),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_508),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_363),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_80),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_353),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_267),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_414),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_159),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_42),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_144),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_247),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_395),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_466),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_29),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_302),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_83),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_93),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_374),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_219),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_462),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_235),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_51),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_92),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_481),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_277),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_114),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_173),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_92),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_147),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_371),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_391),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_491),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_244),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_447),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_511),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_354),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_495),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_373),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_232),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_489),
.Y(n_586)
);

CKINVDCx14_ASAP7_75t_R g587 ( 
.A(n_451),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_361),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_348),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_157),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_486),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_83),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_236),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_352),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_471),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_117),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_421),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_181),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_239),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_179),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_329),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_23),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_328),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_24),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_151),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_492),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_340),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_154),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_287),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_246),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_176),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_305),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_115),
.Y(n_616)
);

BUFx8_ASAP7_75t_SL g617 ( 
.A(n_380),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_244),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_347),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_344),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_185),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_315),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_388),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_193),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_4),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_498),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_196),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_216),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_300),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_496),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_109),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_253),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_502),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_409),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_134),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_246),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_412),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_155),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_325),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_510),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_68),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_49),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_286),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_330),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_406),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_269),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_506),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_166),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_234),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_402),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_332),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_39),
.Y(n_652)
);

CKINVDCx6p67_ASAP7_75t_R g653 ( 
.A(n_319),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_368),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_465),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_485),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_174),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_478),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_381),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_426),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_497),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_156),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_155),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_488),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_268),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_34),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_397),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_386),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_311),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_483),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_403),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_396),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_32),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_142),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_494),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_258),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_157),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_385),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_123),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_440),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_85),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_177),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_224),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_1),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_423),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_110),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_503),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_327),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_480),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_229),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_283),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_32),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_118),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_343),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_84),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_106),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_99),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_280),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_159),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_394),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_512),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_232),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_435),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_487),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_25),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_493),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_154),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_117),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_44),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_505),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_479),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_473),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_125),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_281),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_369),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_270),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_64),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_30),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_89),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_126),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_304),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_292),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_84),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_54),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_97),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_301),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_16),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_499),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_27),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_68),
.Y(n_731)
);

INVxp33_ASAP7_75t_L g732 ( 
.A(n_641),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_514),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_691),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_518),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_522),
.Y(n_736)
);

INVxp33_ASAP7_75t_SL g737 ( 
.A(n_637),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_590),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_522),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_522),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_522),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_522),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_522),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_514),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_522),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_573),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_664),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_515),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_573),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_515),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_628),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_628),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_537),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_706),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_558),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_664),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_715),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_706),
.Y(n_758)
);

INVxp33_ASAP7_75t_SL g759 ( 
.A(n_517),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_607),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_558),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_558),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_558),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_618),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_618),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_520),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_618),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_618),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_598),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_632),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_670),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_632),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_632),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_555),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_632),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_670),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_537),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_718),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_718),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_555),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_718),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_718),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_523),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_524),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_529),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_543),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_593),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_595),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_601),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_602),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_516),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_605),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_525),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_649),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_528),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_677),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_685),
.Y(n_798)
);

INVxp33_ASAP7_75t_L g799 ( 
.A(n_596),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_693),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_703),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_671),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_708),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_721),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_724),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_521),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_530),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_536),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_546),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_671),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_550),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_596),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_608),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_636),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_626),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_553),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_556),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_671),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_569),
.Y(n_820)
);

INVxp33_ASAP7_75t_SL g821 ( 
.A(n_538),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_664),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_636),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_608),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_533),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_574),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_580),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_581),
.Y(n_828)
);

CKINVDCx16_ASAP7_75t_R g829 ( 
.A(n_587),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_586),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_822),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_822),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_778),
.B(n_545),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_747),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_755),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_782),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_771),
.B(n_675),
.Y(n_837)
);

CKINVDCx6p67_ASAP7_75t_R g838 ( 
.A(n_769),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_762),
.Y(n_839)
);

AND2x4_ASAP7_75t_SL g840 ( 
.A(n_796),
.B(n_600),
.Y(n_840)
);

INVx6_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_822),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_747),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_755),
.Y(n_844)
);

AND2x6_ASAP7_75t_L g845 ( 
.A(n_822),
.B(n_664),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_791),
.B(n_513),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_822),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_776),
.B(n_587),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_818),
.B(n_513),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_763),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_761),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_747),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_761),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_733),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_737),
.A2(n_727),
.B1(n_629),
.B2(n_681),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_767),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_737),
.A2(n_541),
.B1(n_544),
.B2(n_540),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_764),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_775),
.B(n_588),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_802),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_816),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_756),
.Y(n_862)
);

OA21x2_ASAP7_75t_L g863 ( 
.A1(n_739),
.A2(n_643),
.B(n_588),
.Y(n_863)
);

INVx6_ASAP7_75t_L g864 ( 
.A(n_756),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_767),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_748),
.B(n_643),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_765),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_756),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_736),
.A2(n_680),
.B(n_591),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_732),
.A2(n_552),
.B1(n_554),
.B2(n_551),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_756),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_775),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_736),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_775),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_748),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_768),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_741),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_770),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_772),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_742),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_750),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_750),
.B(n_700),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_807),
.B(n_680),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_743),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_745),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_829),
.B(n_589),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_733),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_773),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_808),
.B(n_592),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_779),
.Y(n_891)
);

BUFx12f_ASAP7_75t_L g892 ( 
.A(n_744),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_781),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_809),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_810),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_760),
.A2(n_629),
.B1(n_681),
.B2(n_600),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_873),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_877),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_835),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_873),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_840),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_875),
.Y(n_902)
);

OAI21x1_ASAP7_75t_L g903 ( 
.A1(n_869),
.A2(n_817),
.B(n_812),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_877),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_873),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_833),
.B(n_744),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_835),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_878),
.Y(n_908)
);

INVx6_ASAP7_75t_L g909 ( 
.A(n_868),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_896),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_878),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_890),
.B(n_820),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_846),
.A2(n_738),
.B1(n_757),
.B2(n_732),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_885),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_844),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_885),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_843),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_833),
.B(n_826),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_833),
.B(n_827),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_875),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_886),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_886),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_881),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_883),
.B(n_774),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_883),
.B(n_774),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_881),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_844),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_860),
.B(n_759),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_881),
.Y(n_930)
);

OA21x2_ASAP7_75t_L g931 ( 
.A1(n_869),
.A2(n_830),
.B(n_828),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_839),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_882),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_850),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_863),
.A2(n_615),
.B(n_606),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_882),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_843),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_846),
.B(n_799),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_848),
.B(n_766),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_858),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_887),
.B(n_759),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_836),
.B(n_821),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_851),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_867),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_851),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_890),
.B(n_859),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_880),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_853),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_846),
.B(n_780),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_853),
.Y(n_950)
);

OA21x2_ASAP7_75t_L g951 ( 
.A1(n_866),
.A2(n_813),
.B(n_815),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_840),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_859),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_856),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_837),
.B(n_766),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_843),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_882),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_874),
.B(n_783),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_856),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_859),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_865),
.Y(n_961)
);

NOR2x1_ASAP7_75t_L g962 ( 
.A(n_868),
.B(n_542),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_865),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_894),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_895),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_889),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_889),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_862),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_890),
.B(n_884),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_843),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_862),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_874),
.B(n_783),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_874),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_862),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_884),
.B(n_813),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_884),
.B(n_780),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_849),
.B(n_799),
.Y(n_977)
);

AND2x6_ASAP7_75t_L g978 ( 
.A(n_832),
.B(n_622),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_874),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_863),
.B(n_815),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_842),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_832),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_834),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_863),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_941),
.B(n_821),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_905),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_905),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_946),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_938),
.B(n_727),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_832),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_938),
.B(n_949),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_980),
.A2(n_857),
.B1(n_640),
.B2(n_646),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_984),
.B(n_831),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_953),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_946),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_962),
.B(n_845),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_925),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_949),
.B(n_861),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_925),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_953),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_960),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_960),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_946),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_942),
.Y(n_1004)
);

AND2x2_ASAP7_75t_SL g1005 ( 
.A(n_910),
.B(n_855),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_909),
.Y(n_1006)
);

CKINVDCx11_ASAP7_75t_R g1007 ( 
.A(n_901),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_926),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_909),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_964),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_926),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_964),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_905),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_965),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_897),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_965),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_962),
.A2(n_568),
.B1(n_584),
.B2(n_557),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_975),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_897),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_902),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_975),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_984),
.B(n_831),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_980),
.B(n_831),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_955),
.B(n_760),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_975),
.Y(n_1025)
);

INVx6_ASAP7_75t_L g1026 ( 
.A(n_946),
.Y(n_1026)
);

INVx4_ASAP7_75t_SL g1027 ( 
.A(n_978),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_921),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_897),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_913),
.B(n_939),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_977),
.B(n_879),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_977),
.B(n_784),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_897),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_976),
.B(n_784),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_900),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_976),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_912),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_906),
.B(n_793),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_933),
.B(n_861),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_975),
.Y(n_1040)
);

AND3x2_ASAP7_75t_L g1041 ( 
.A(n_933),
.B(n_734),
.C(n_719),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_919),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_900),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_903),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_969),
.B(n_785),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_932),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_969),
.B(n_793),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_932),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_912),
.A2(n_644),
.B1(n_655),
.B2(n_650),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_934),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_958),
.B(n_854),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_912),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_910),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_929),
.B(n_870),
.C(n_735),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_934),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_931),
.Y(n_1056)
);

AND2x2_ASAP7_75t_SL g1057 ( 
.A(n_972),
.B(n_700),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_912),
.A2(n_661),
.B1(n_665),
.B2(n_658),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_920),
.B(n_936),
.Y(n_1059)
);

INVxp33_ASAP7_75t_L g1060 ( 
.A(n_940),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_940),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_900),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_957),
.B(n_854),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_931),
.B(n_672),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_944),
.Y(n_1065)
);

AND2x2_ASAP7_75t_SL g1066 ( 
.A(n_931),
.B(n_719),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_944),
.B(n_888),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_952),
.B(n_802),
.Y(n_1068)
);

BUFx8_ASAP7_75t_SL g1069 ( 
.A(n_947),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_947),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_973),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_973),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_979),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_951),
.B(n_811),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_903),
.B(n_888),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_924),
.B(n_879),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_909),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_924),
.B(n_879),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_931),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_967),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_967),
.B(n_838),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_898),
.B(n_892),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_927),
.B(n_879),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_927),
.B(n_893),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_951),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_930),
.A2(n_635),
.B1(n_728),
.B2(n_527),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_930),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_966),
.B(n_838),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_979),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_951),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_898),
.B(n_893),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_904),
.B(n_893),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_904),
.A2(n_699),
.B1(n_713),
.B2(n_690),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_908),
.B(n_893),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_908),
.B(n_786),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_900),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_966),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_911),
.B(n_892),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_899),
.Y(n_1099)
);

BUFx8_ASAP7_75t_SL g1100 ( 
.A(n_982),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_951),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_968),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_911),
.B(n_876),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_899),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_914),
.A2(n_728),
.B1(n_635),
.B2(n_687),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_907),
.Y(n_1106)
);

BUFx10_ASAP7_75t_L g1107 ( 
.A(n_914),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_917),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_917),
.B(n_597),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_922),
.B(n_876),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_922),
.B(n_811),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_923),
.B(n_787),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_923),
.B(n_819),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_978),
.A2(n_652),
.B1(n_594),
.B2(n_560),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_961),
.B(n_876),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_909),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_907),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_968),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_971),
.B(n_819),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_961),
.B(n_876),
.Y(n_1120)
);

NAND3x1_ASAP7_75t_L g1121 ( 
.A(n_971),
.B(n_789),
.C(n_788),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_983),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1104),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_985),
.B(n_825),
.C(n_749),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_997),
.B(n_692),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_997),
.B(n_746),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1031),
.B(n_974),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1031),
.B(n_974),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1032),
.B(n_777),
.C(n_753),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1018),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1011),
.B(n_915),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1011),
.B(n_716),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1104),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_999),
.B(n_751),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_L g1135 ( 
.A(n_989),
.B(n_998),
.C(n_1024),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_991),
.A2(n_978),
.B1(n_982),
.B2(n_928),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1006),
.A2(n_935),
.B(n_981),
.Y(n_1137)
);

NOR3xp33_ASAP7_75t_L g1138 ( 
.A(n_1039),
.B(n_754),
.C(n_752),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1021),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_1068),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1042),
.B(n_915),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_988),
.B(n_995),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1106),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1030),
.B(n_519),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1025),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1036),
.B(n_526),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1040),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1042),
.B(n_915),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1037),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1036),
.A2(n_978),
.B1(n_918),
.B2(n_956),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1008),
.B(n_1057),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1020),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1052),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_994),
.B(n_915),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1038),
.B(n_531),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1106),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1000),
.Y(n_1157)
);

BUFx8_ASAP7_75t_L g1158 ( 
.A(n_1034),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_988),
.B(n_532),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1001),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1002),
.B(n_918),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_995),
.B(n_918),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1045),
.B(n_790),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1004),
.B(n_753),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1054),
.B(n_814),
.C(n_777),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1047),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1028),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1087),
.Y(n_1168)
);

INVx8_ASAP7_75t_L g1169 ( 
.A(n_1075),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1003),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1003),
.B(n_1060),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1006),
.B(n_534),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1026),
.A2(n_978),
.B1(n_956),
.B2(n_918),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1026),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1010),
.B(n_956),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1012),
.B(n_956),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1108),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1004),
.B(n_814),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1014),
.B(n_1016),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1045),
.B(n_792),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1017),
.B(n_824),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1009),
.B(n_535),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1046),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1048),
.B(n_916),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1054),
.A2(n_978),
.B1(n_916),
.B2(n_943),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1066),
.A2(n_978),
.B1(n_928),
.B2(n_945),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1118),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1050),
.B(n_943),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1055),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1088),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1061),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1065),
.B(n_945),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1111),
.B(n_824),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1113),
.B(n_1067),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1070),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1023),
.B(n_948),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1009),
.B(n_539),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1095),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1023),
.B(n_948),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1099),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1026),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1097),
.B(n_950),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1100),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1077),
.B(n_548),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1077),
.B(n_1116),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1116),
.B(n_1107),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1117),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1095),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1112),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1112),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1107),
.B(n_1051),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1015),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1056),
.B(n_950),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1080),
.B(n_549),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1063),
.B(n_758),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1056),
.B(n_954),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1019),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1109),
.B(n_547),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1029),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1033),
.Y(n_1220)
);

O2A1O1Ixp5_ASAP7_75t_L g1221 ( 
.A1(n_1074),
.A2(n_1119),
.B(n_1076),
.C(n_1083),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1059),
.B(n_570),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_993),
.B(n_954),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1081),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1075),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_992),
.B(n_559),
.Y(n_1226)
);

AOI22x1_ASAP7_75t_R g1227 ( 
.A1(n_1053),
.A2(n_794),
.B1(n_797),
.B2(n_795),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_993),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1071),
.Y(n_1229)
);

INVx8_ASAP7_75t_L g1230 ( 
.A(n_1075),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1005),
.B(n_617),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1035),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1079),
.A2(n_963),
.B(n_959),
.C(n_798),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1022),
.B(n_959),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1022),
.B(n_963),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1043),
.Y(n_1236)
);

AND2x2_ASAP7_75t_SL g1237 ( 
.A(n_1114),
.B(n_617),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1062),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1096),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1102),
.B(n_983),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1082),
.B(n_561),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1079),
.B(n_983),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1041),
.B(n_1098),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1086),
.B(n_1041),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_990),
.A2(n_935),
.B(n_564),
.C(n_575),
.Y(n_1245)
);

NOR2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1069),
.B(n_653),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1027),
.B(n_800),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1072),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1007),
.Y(n_1249)
);

NAND2xp33_ASAP7_75t_L g1250 ( 
.A(n_1044),
.B(n_937),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1049),
.B(n_1058),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1101),
.B(n_983),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1076),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1101),
.B(n_983),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1071),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1073),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1078),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1089),
.B(n_983),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1090),
.B(n_937),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1090),
.B(n_937),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1027),
.B(n_801),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1122),
.B(n_562),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1122),
.B(n_576),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1086),
.B(n_563),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1105),
.B(n_1091),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1073),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1078),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1091),
.A2(n_1094),
.B1(n_1092),
.B2(n_1084),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1105),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1085),
.A2(n_804),
.B(n_805),
.C(n_803),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_L g1271 ( 
.A(n_1093),
.B(n_996),
.C(n_566),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_990),
.B(n_565),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1083),
.A2(n_579),
.B1(n_582),
.B2(n_578),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1084),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_986),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1092),
.B(n_583),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1094),
.B(n_937),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_987),
.B(n_1013),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1103),
.B(n_937),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1103),
.A2(n_609),
.B1(n_610),
.B2(n_604),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_SL g1281 ( 
.A(n_1044),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1110),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1110),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1115),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1115),
.B(n_937),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1120),
.B(n_970),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1027),
.B(n_612),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1121),
.A2(n_620),
.B1(n_623),
.B2(n_619),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1064),
.B(n_806),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1064),
.A2(n_621),
.B1(n_638),
.B2(n_572),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1120),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1044),
.B(n_630),
.Y(n_1292)
);

AO221x1_ASAP7_75t_L g1293 ( 
.A1(n_1105),
.A2(n_970),
.B1(n_871),
.B2(n_852),
.C(n_834),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1031),
.B(n_970),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1031),
.B(n_970),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1037),
.B(n_970),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1068),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_985),
.B(n_567),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_985),
.B(n_577),
.C(n_571),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_L g1300 ( 
.A(n_1030),
.B(n_970),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_997),
.B(n_633),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1031),
.B(n_634),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1018),
.Y(n_1303)
);

AOI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1105),
.A2(n_611),
.B1(n_613),
.B2(n_599),
.C(n_585),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1031),
.B(n_639),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1104),
.Y(n_1306)
);

AND2x6_ASAP7_75t_L g1307 ( 
.A(n_1090),
.B(n_823),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_985),
.B(n_614),
.C(n_603),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1031),
.B(n_645),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1030),
.A2(n_657),
.B1(n_684),
.B2(n_627),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_997),
.B(n_647),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1053),
.A2(n_662),
.B1(n_694),
.B2(n_631),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_985),
.B(n_624),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1031),
.B(n_651),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1068),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_991),
.A2(n_823),
.B(n_656),
.C(n_659),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_985),
.B(n_642),
.C(n_625),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1018),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1031),
.B(n_654),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1031),
.B(n_660),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1104),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_991),
.A2(n_668),
.B(n_669),
.C(n_667),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_985),
.B(n_648),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1169),
.B(n_868),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1228),
.B(n_1298),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1284),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1313),
.A2(n_678),
.B1(n_686),
.B2(n_676),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1152),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1291),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1184),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1174),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1130),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1149),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1323),
.A2(n_689),
.B1(n_695),
.B2(n_688),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1157),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1272),
.B(n_1253),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1160),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1225),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1257),
.B(n_1267),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1193),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1274),
.B(n_701),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1174),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1194),
.B(n_663),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1167),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1222),
.A2(n_704),
.B(n_705),
.C(n_702),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1282),
.B(n_707),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1149),
.B(n_834),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1135),
.A2(n_712),
.B1(n_717),
.B2(n_711),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1187),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1283),
.B(n_722),
.Y(n_1350)
);

NAND2xp33_ASAP7_75t_SL g1351 ( 
.A(n_1281),
.B(n_723),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1225),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1183),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1189),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1190),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1191),
.Y(n_1356)
);

NAND2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1149),
.B(n_834),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1166),
.A2(n_729),
.B1(n_891),
.B2(n_876),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1179),
.B(n_666),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1195),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1134),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1158),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1139),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1158),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1145),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1153),
.B(n_673),
.Y(n_1366)
);

AND2x2_ASAP7_75t_SL g1367 ( 
.A(n_1181),
.B(n_0),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1265),
.B(n_674),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1177),
.B(n_679),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1153),
.B(n_852),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1153),
.B(n_852),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1249),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1131),
.B(n_682),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1251),
.A2(n_891),
.B1(n_696),
.B2(n_697),
.Y(n_1374)
);

NOR2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1129),
.B(n_683),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1125),
.B(n_1132),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1225),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1178),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1147),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1303),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1318),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1168),
.B(n_698),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1165),
.A2(n_891),
.B1(n_710),
.B2(n_714),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1163),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1227),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1188),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1275),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1192),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1169),
.B(n_891),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1202),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1123),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1302),
.B(n_709),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1305),
.B(n_725),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1164),
.B(n_726),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1200),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1133),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1143),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1201),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1163),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1156),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1203),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1180),
.Y(n_1402)
);

NOR2x1p5_ASAP7_75t_L g1403 ( 
.A(n_1198),
.B(n_730),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1306),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1180),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1169),
.B(n_891),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1309),
.B(n_731),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1140),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1314),
.B(n_845),
.Y(n_1409)
);

BUFx4f_ASAP7_75t_L g1410 ( 
.A(n_1230),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1297),
.B(n_1),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1201),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1207),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1218),
.B(n_2),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1208),
.B(n_256),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1127),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1128),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1321),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1255),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1315),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1319),
.B(n_845),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1256),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1320),
.B(n_845),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1201),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1209),
.B(n_257),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1175),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1176),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1215),
.B(n_845),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1248),
.B(n_852),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1170),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1224),
.B(n_2),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1269),
.A2(n_872),
.B1(n_864),
.B2(n_841),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1266),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1220),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1126),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1236),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1229),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1229),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1141),
.B(n_845),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1210),
.B(n_259),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1230),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1211),
.B(n_1231),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1212),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1281),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1217),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1151),
.A2(n_864),
.B1(n_841),
.B2(n_872),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1219),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1230),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1232),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1238),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1248),
.B(n_871),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1248),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1239),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1264),
.A2(n_864),
.B1(n_841),
.B2(n_871),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1148),
.B(n_3),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1247),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1278),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1196),
.B(n_3),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1244),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1243),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1154),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1243),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_SL g1463 ( 
.A(n_1237),
.Y(n_1463)
);

NOR3xp33_ASAP7_75t_SL g1464 ( 
.A(n_1312),
.B(n_4),
.C(n_5),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1247),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1161),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1213),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1171),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1296),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1299),
.B(n_871),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1144),
.A2(n_864),
.B1(n_841),
.B2(n_872),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1308),
.A2(n_872),
.B1(n_981),
.B2(n_847),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1261),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1241),
.A2(n_872),
.B(n_7),
.C(n_5),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1270),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1199),
.B(n_6),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1294),
.B(n_6),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1261),
.B(n_260),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1295),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1268),
.B(n_7),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1252),
.B(n_8),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1240),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1317),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1216),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1258),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1242),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1246),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1226),
.A2(n_981),
.B1(n_847),
.B2(n_842),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1254),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1142),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1142),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1310),
.B(n_8),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1223),
.B(n_9),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1289),
.Y(n_1494)
);

AND2x6_ASAP7_75t_SL g1495 ( 
.A(n_1289),
.B(n_9),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1304),
.B(n_10),
.C(n_11),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1307),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1277),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1279),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1301),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1285),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1290),
.A2(n_981),
.B1(n_847),
.B2(n_842),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1206),
.B(n_262),
.Y(n_1503)
);

NAND2xp33_ASAP7_75t_L g1504 ( 
.A(n_1307),
.B(n_1205),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1280),
.B(n_1155),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1289),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1311),
.B(n_263),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1286),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1271),
.A2(n_847),
.B1(n_842),
.B2(n_12),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1293),
.A2(n_847),
.B1(n_842),
.B2(n_12),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1234),
.B(n_10),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1235),
.B(n_11),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1288),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1146),
.B(n_13),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1288),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1307),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1307),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1214),
.B(n_13),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1259),
.B(n_14),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1280),
.B(n_264),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1150),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1162),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1260),
.B(n_14),
.Y(n_1523)
);

XOR2xp5_ASAP7_75t_L g1524 ( 
.A(n_1159),
.B(n_265),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1162),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1273),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1173),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1124),
.B(n_1138),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1292),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1221),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1185),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1276),
.B(n_15),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1435),
.B(n_1322),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1325),
.B(n_1316),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1416),
.B(n_1300),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_SL g1536 ( 
.A(n_1513),
.B(n_1172),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1367),
.B(n_1136),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1526),
.B(n_1186),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1452),
.B(n_1182),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1336),
.B(n_1197),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1416),
.B(n_1204),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1378),
.B(n_1262),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1361),
.B(n_1263),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1376),
.B(n_1233),
.Y(n_1544)
);

NAND2xp33_ASAP7_75t_SL g1545 ( 
.A(n_1452),
.B(n_1441),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1442),
.B(n_1245),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1459),
.B(n_1287),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1515),
.B(n_1340),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1528),
.B(n_1137),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1408),
.B(n_1250),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1394),
.B(n_17),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1452),
.B(n_18),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_SL g1553 ( 
.A(n_1441),
.B(n_18),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1402),
.B(n_19),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1405),
.B(n_19),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1500),
.B(n_20),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1349),
.B(n_21),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1483),
.B(n_21),
.Y(n_1558)
);

NAND2xp33_ASAP7_75t_SL g1559 ( 
.A(n_1441),
.B(n_22),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1507),
.B(n_22),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1507),
.B(n_23),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1462),
.B(n_24),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1417),
.B(n_25),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1417),
.B(n_26),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1384),
.B(n_26),
.Y(n_1565)
);

NAND2xp33_ASAP7_75t_SL g1566 ( 
.A(n_1448),
.B(n_27),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1399),
.B(n_28),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1415),
.B(n_28),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1415),
.B(n_29),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1425),
.B(n_30),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1425),
.B(n_31),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1440),
.B(n_31),
.Y(n_1572)
);

NAND2xp33_ASAP7_75t_SL g1573 ( 
.A(n_1448),
.B(n_33),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1440),
.B(n_33),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1355),
.B(n_34),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1420),
.B(n_35),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1343),
.B(n_35),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1414),
.B(n_36),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_SL g1579 ( 
.A(n_1448),
.B(n_36),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1344),
.B(n_37),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1468),
.B(n_37),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1339),
.B(n_38),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1328),
.B(n_38),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1463),
.B(n_39),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1390),
.B(n_40),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1529),
.B(n_1333),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_SL g1587 ( 
.A(n_1463),
.B(n_40),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1333),
.B(n_41),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1332),
.B(n_41),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1444),
.B(n_42),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1365),
.B(n_43),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_SL g1592 ( 
.A(n_1444),
.B(n_44),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1473),
.B(n_266),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1392),
.B(n_45),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1393),
.B(n_45),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1407),
.B(n_46),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1388),
.B(n_46),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1326),
.B(n_47),
.Y(n_1598)
);

NAND2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1531),
.B(n_47),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1326),
.B(n_48),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_SL g1601 ( 
.A(n_1338),
.B(n_48),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1338),
.B(n_49),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1465),
.B(n_271),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1329),
.B(n_50),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1329),
.B(n_50),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_SL g1606 ( 
.A(n_1338),
.B(n_51),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1359),
.B(n_52),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1385),
.B(n_53),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1489),
.B(n_53),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1514),
.B(n_54),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1494),
.B(n_1506),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1352),
.B(n_55),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1506),
.B(n_55),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1520),
.B(n_56),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1330),
.B(n_56),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1330),
.B(n_57),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1386),
.B(n_1335),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1352),
.B(n_57),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1352),
.B(n_58),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1386),
.B(n_59),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1337),
.B(n_60),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1353),
.B(n_61),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1354),
.B(n_61),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1356),
.B(n_62),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1360),
.B(n_62),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1518),
.B(n_63),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1505),
.B(n_64),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1492),
.B(n_65),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1341),
.B(n_65),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1410),
.B(n_66),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1410),
.B(n_66),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1456),
.B(n_67),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1456),
.B(n_1424),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_SL g1634 ( 
.A(n_1377),
.B(n_67),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1456),
.B(n_69),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1424),
.B(n_69),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1424),
.B(n_70),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1346),
.B(n_70),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1350),
.B(n_71),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1467),
.B(n_71),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1497),
.B(n_72),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1497),
.B(n_73),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1497),
.B(n_73),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1363),
.B(n_1379),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1373),
.B(n_74),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1380),
.B(n_74),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1381),
.B(n_75),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1368),
.B(n_75),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1331),
.B(n_76),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1467),
.B(n_76),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1331),
.B(n_77),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1342),
.B(n_77),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1342),
.B(n_78),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1532),
.B(n_78),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1348),
.B(n_79),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1398),
.B(n_272),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1375),
.B(n_81),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1457),
.B(n_1377),
.Y(n_1658)
);

NAND2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1377),
.B(n_81),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1327),
.B(n_82),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1411),
.B(n_1431),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1478),
.B(n_82),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1478),
.B(n_85),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1395),
.B(n_86),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1413),
.B(n_86),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1490),
.B(n_1491),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1479),
.B(n_87),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1403),
.B(n_87),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1484),
.B(n_88),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1369),
.B(n_1382),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1464),
.B(n_88),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1516),
.B(n_90),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1516),
.B(n_1434),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1486),
.B(n_90),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1516),
.B(n_91),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1436),
.B(n_91),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1437),
.B(n_93),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1437),
.B(n_94),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1438),
.B(n_94),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1438),
.B(n_95),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1391),
.B(n_95),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1499),
.B(n_96),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1396),
.B(n_96),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1397),
.B(n_97),
.Y(n_1684)
);

NAND2xp33_ASAP7_75t_SL g1685 ( 
.A(n_1487),
.B(n_98),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1400),
.B(n_98),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1404),
.B(n_99),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1419),
.B(n_100),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1501),
.B(n_100),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1422),
.B(n_101),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1433),
.B(n_101),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1387),
.B(n_102),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1480),
.B(n_102),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1398),
.B(n_103),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1412),
.B(n_103),
.Y(n_1695)
);

NAND2xp33_ASAP7_75t_SL g1696 ( 
.A(n_1364),
.B(n_104),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_SL g1697 ( 
.A(n_1366),
.B(n_104),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1412),
.B(n_273),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1475),
.B(n_105),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1508),
.B(n_105),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1334),
.B(n_106),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1418),
.B(n_1447),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1383),
.B(n_1443),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1445),
.B(n_107),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1498),
.B(n_107),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1449),
.B(n_108),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1450),
.B(n_1453),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1458),
.B(n_108),
.Y(n_1708)
);

NAND2xp33_ASAP7_75t_SL g1709 ( 
.A(n_1372),
.B(n_109),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1426),
.B(n_110),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1430),
.B(n_111),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1427),
.B(n_111),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1476),
.B(n_112),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_SL g1714 ( 
.A(n_1401),
.B(n_112),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1461),
.B(n_113),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1466),
.B(n_113),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1345),
.B(n_114),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1469),
.B(n_115),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1521),
.B(n_116),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1324),
.B(n_274),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1493),
.B(n_116),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1482),
.B(n_118),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1511),
.B(n_119),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1512),
.B(n_119),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1455),
.B(n_120),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_L g1726 ( 
.A(n_1655),
.B(n_1661),
.C(n_1628),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1714),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1585),
.B(n_1524),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1541),
.B(n_1496),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1644),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1670),
.B(n_1481),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1656),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1707),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1599),
.A2(n_1660),
.B1(n_1701),
.B2(n_1693),
.Y(n_1734)
);

NOR2xp67_ASAP7_75t_L g1735 ( 
.A(n_1540),
.B(n_1477),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1537),
.B(n_1374),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1626),
.A2(n_1474),
.B1(n_1527),
.B2(n_1460),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1593),
.B(n_1324),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1645),
.B(n_1519),
.Y(n_1739)
);

NAND2x1p5_ASAP7_75t_L g1740 ( 
.A(n_1586),
.B(n_1362),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1702),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1610),
.A2(n_1527),
.B1(n_1509),
.B2(n_1351),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1538),
.B(n_1523),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1548),
.B(n_1485),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1711),
.B(n_1347),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1550),
.A2(n_1535),
.B1(n_1543),
.B2(n_1547),
.Y(n_1746)
);

BUFx12f_ASAP7_75t_L g1747 ( 
.A(n_1648),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_R g1748 ( 
.A(n_1536),
.B(n_1495),
.Y(n_1748)
);

NAND2x1p5_ASAP7_75t_L g1749 ( 
.A(n_1593),
.B(n_1503),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1560),
.B(n_1470),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1640),
.Y(n_1751)
);

INVx4_ASAP7_75t_L g1752 ( 
.A(n_1656),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1650),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1617),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1667),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1682),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1544),
.B(n_1522),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1597),
.A2(n_1712),
.B1(n_1710),
.B2(n_1700),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1657),
.Y(n_1759)
);

AOI22x1_ASAP7_75t_L g1760 ( 
.A1(n_1720),
.A2(n_1530),
.B1(n_1525),
.B2(n_1517),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1654),
.B(n_1357),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1561),
.A2(n_1510),
.B1(n_1389),
.B2(n_1406),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1719),
.A2(n_1428),
.B1(n_1358),
.B2(n_1504),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1611),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1593),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1705),
.B(n_1429),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1689),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1563),
.B(n_1370),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1609),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1546),
.A2(n_1421),
.B(n_1409),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1674),
.B(n_1451),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1656),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1568),
.B(n_1432),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1564),
.B(n_1371),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1584),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1569),
.B(n_1389),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1698),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1722),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1662),
.B(n_1406),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1658),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1720),
.B(n_1446),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1627),
.B(n_1454),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1698),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1572),
.B(n_1471),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1666),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1574),
.B(n_1423),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1582),
.B(n_1615),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1663),
.B(n_1439),
.Y(n_1789)
);

BUFx12f_ASAP7_75t_L g1790 ( 
.A(n_1720),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1671),
.A2(n_1558),
.B1(n_1699),
.B2(n_1551),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1673),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1633),
.B(n_1472),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1616),
.B(n_120),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1708),
.B(n_121),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1587),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1713),
.B(n_121),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1698),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1703),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1685),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1577),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1669),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1697),
.A2(n_1502),
.B1(n_1488),
.B2(n_124),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1721),
.B(n_122),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1603),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1603),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1614),
.B(n_122),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1603),
.Y(n_1808)
);

CKINVDCx8_ASAP7_75t_R g1809 ( 
.A(n_1545),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1620),
.B(n_123),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1715),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1578),
.B(n_124),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1549),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1716),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1598),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1723),
.B(n_125),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1542),
.B(n_275),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1696),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1533),
.B(n_1613),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1629),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1668),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1600),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1604),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1724),
.B(n_130),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1539),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1534),
.A2(n_278),
.B(n_276),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1725),
.B(n_131),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1562),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1605),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1709),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1641),
.B(n_279),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1590),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1608),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1607),
.B(n_132),
.Y(n_1834)
);

AND3x1_ASAP7_75t_SL g1835 ( 
.A(n_1592),
.B(n_133),
.C(n_134),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1717),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1601),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1681),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1683),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1602),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1684),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1594),
.A2(n_1595),
.B1(n_1596),
.B2(n_1638),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1639),
.A2(n_284),
.B(n_282),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1581),
.B(n_135),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1621),
.B(n_1622),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1718),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1623),
.B(n_136),
.Y(n_1847)
);

O2A1O1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1556),
.A2(n_1631),
.B(n_1630),
.C(n_1580),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1686),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1687),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1624),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1625),
.B(n_1646),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1688),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1647),
.B(n_138),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1690),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1691),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1676),
.B(n_139),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1642),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_1858)
);

NAND2x1_ASAP7_75t_L g1859 ( 
.A(n_1606),
.B(n_285),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1692),
.Y(n_1860)
);

BUFx10_ASAP7_75t_L g1861 ( 
.A(n_1583),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1664),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1589),
.B(n_140),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1694),
.Y(n_1864)
);

AND3x1_ASAP7_75t_SL g1865 ( 
.A(n_1557),
.B(n_141),
.C(n_143),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1695),
.B(n_288),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1591),
.B(n_143),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1665),
.A2(n_290),
.B(n_289),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1704),
.B(n_144),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1706),
.Y(n_1870)
);

INVx5_ASAP7_75t_L g1871 ( 
.A(n_1612),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1677),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1680),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1643),
.A2(n_1554),
.B1(n_1555),
.B2(n_1672),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1678),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1632),
.B(n_145),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1635),
.B(n_145),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1636),
.B(n_146),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1679),
.Y(n_1879)
);

AND3x1_ASAP7_75t_SL g1880 ( 
.A(n_1576),
.B(n_146),
.C(n_147),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1565),
.B(n_148),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1553),
.B(n_1559),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1567),
.B(n_148),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1649),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1618),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1651),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1637),
.B(n_149),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1566),
.B(n_150),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1552),
.B(n_152),
.Y(n_1889)
);

INVx5_ASAP7_75t_L g1890 ( 
.A(n_1619),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1751),
.B(n_1652),
.Y(n_1891)
);

BUFx12f_ASAP7_75t_L g1892 ( 
.A(n_1759),
.Y(n_1892)
);

AOI22x1_ASAP7_75t_L g1893 ( 
.A1(n_1826),
.A2(n_1843),
.B1(n_1868),
.B2(n_1825),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1813),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1799),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1739),
.A2(n_1653),
.B(n_1588),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1780),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1790),
.Y(n_1898)
);

OAI21x1_ASAP7_75t_L g1899 ( 
.A1(n_1770),
.A2(n_1675),
.B(n_1575),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1770),
.A2(n_1659),
.B(n_1634),
.Y(n_1900)
);

OA21x2_ASAP7_75t_L g1901 ( 
.A1(n_1757),
.A2(n_1579),
.B(n_1573),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1726),
.A2(n_1758),
.B1(n_1832),
.B2(n_1734),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1747),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1733),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1741),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1730),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1753),
.B(n_152),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1754),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1760),
.A2(n_293),
.B(n_291),
.Y(n_1909)
);

BUFx12f_ASAP7_75t_L g1910 ( 
.A(n_1861),
.Y(n_1910)
);

INVx3_ASAP7_75t_SL g1911 ( 
.A(n_1727),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1757),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1786),
.Y(n_1913)
);

BUFx5_ASAP7_75t_L g1914 ( 
.A(n_1792),
.Y(n_1914)
);

CKINVDCx6p67_ASAP7_75t_R g1915 ( 
.A(n_1861),
.Y(n_1915)
);

INVx5_ASAP7_75t_L g1916 ( 
.A(n_1825),
.Y(n_1916)
);

AO21x2_ASAP7_75t_L g1917 ( 
.A1(n_1735),
.A2(n_153),
.B(n_156),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1735),
.A2(n_153),
.B(n_158),
.Y(n_1918)
);

OR2x6_ASAP7_75t_L g1919 ( 
.A(n_1765),
.B(n_294),
.Y(n_1919)
);

AOI22x1_ASAP7_75t_L g1920 ( 
.A1(n_1826),
.A2(n_161),
.B1(n_158),
.B2(n_160),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1765),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1744),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1740),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1764),
.Y(n_1924)
);

AOI22x1_ASAP7_75t_L g1925 ( 
.A1(n_1843),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1793),
.A2(n_1731),
.B(n_1763),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1809),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1738),
.Y(n_1928)
);

OAI21x1_ASAP7_75t_L g1929 ( 
.A1(n_1763),
.A2(n_296),
.B(n_295),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1745),
.Y(n_1930)
);

BUFx8_ASAP7_75t_L g1931 ( 
.A(n_1728),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1743),
.A2(n_162),
.B(n_163),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1738),
.Y(n_1933)
);

AO21x2_ASAP7_75t_L g1934 ( 
.A1(n_1729),
.A2(n_163),
.B(n_164),
.Y(n_1934)
);

OR3x4_ASAP7_75t_SL g1935 ( 
.A(n_1748),
.B(n_164),
.C(n_165),
.Y(n_1935)
);

NAND2x1p5_ASAP7_75t_L g1936 ( 
.A(n_1752),
.B(n_297),
.Y(n_1936)
);

BUFx2_ASAP7_75t_R g1937 ( 
.A(n_1800),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1765),
.B(n_298),
.Y(n_1938)
);

INVx8_ASAP7_75t_L g1939 ( 
.A(n_1846),
.Y(n_1939)
);

OAI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1732),
.A2(n_303),
.B(n_299),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1808),
.Y(n_1941)
);

INVxp67_ASAP7_75t_SL g1942 ( 
.A(n_1732),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1808),
.Y(n_1943)
);

NAND2x1p5_ASAP7_75t_L g1944 ( 
.A(n_1752),
.B(n_306),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1772),
.B(n_307),
.Y(n_1945)
);

INVx4_ASAP7_75t_L g1946 ( 
.A(n_1871),
.Y(n_1946)
);

INVx4_ASAP7_75t_L g1947 ( 
.A(n_1871),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1749),
.A2(n_309),
.B(n_308),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1755),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_1833),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1736),
.B(n_310),
.Y(n_1951)
);

INVx5_ASAP7_75t_L g1952 ( 
.A(n_1871),
.Y(n_1952)
);

BUFx12f_ASAP7_75t_L g1953 ( 
.A(n_1775),
.Y(n_1953)
);

OAI21x1_ASAP7_75t_L g1954 ( 
.A1(n_1746),
.A2(n_1806),
.B(n_1805),
.Y(n_1954)
);

NAND2x1p5_ASAP7_75t_L g1955 ( 
.A(n_1890),
.B(n_312),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1808),
.Y(n_1956)
);

CKINVDCx14_ASAP7_75t_R g1957 ( 
.A(n_1818),
.Y(n_1957)
);

INVx4_ASAP7_75t_L g1958 ( 
.A(n_1890),
.Y(n_1958)
);

INVx6_ASAP7_75t_L g1959 ( 
.A(n_1846),
.Y(n_1959)
);

BUFx12f_ASAP7_75t_L g1960 ( 
.A(n_1796),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1777),
.B(n_313),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1769),
.B(n_165),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1864),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1756),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1830),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1767),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1784),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1773),
.A2(n_1787),
.B(n_1762),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1846),
.Y(n_1969)
);

INVx1_ASAP7_75t_SL g1970 ( 
.A(n_1761),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1819),
.Y(n_1971)
);

INVx6_ASAP7_75t_SL g1972 ( 
.A(n_1819),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1815),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1798),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1801),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1778),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1781),
.Y(n_1977)
);

NAND2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1890),
.B(n_314),
.Y(n_1978)
);

AOI22x1_ASAP7_75t_L g1979 ( 
.A1(n_1868),
.A2(n_1831),
.B1(n_1782),
.B2(n_1829),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1737),
.A2(n_166),
.B(n_167),
.Y(n_1980)
);

AO21x2_ASAP7_75t_L g1981 ( 
.A1(n_1783),
.A2(n_167),
.B(n_168),
.Y(n_1981)
);

BUFx5_ASAP7_75t_L g1982 ( 
.A(n_1822),
.Y(n_1982)
);

CKINVDCx11_ASAP7_75t_R g1983 ( 
.A(n_1866),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1837),
.B(n_316),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1828),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1758),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_1986)
);

CKINVDCx14_ASAP7_75t_R g1987 ( 
.A(n_1812),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1823),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1776),
.Y(n_1989)
);

OAI21x1_ASAP7_75t_L g1990 ( 
.A1(n_1789),
.A2(n_320),
.B(n_318),
.Y(n_1990)
);

NAND2x1p5_ASAP7_75t_L g1991 ( 
.A(n_1837),
.B(n_321),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1802),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1788),
.B(n_1750),
.Y(n_1993)
);

BUFx12f_ASAP7_75t_L g1994 ( 
.A(n_1866),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1811),
.Y(n_1995)
);

BUFx2_ASAP7_75t_SL g1996 ( 
.A(n_1840),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1768),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1906),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1913),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_SL g2000 ( 
.A1(n_1980),
.A2(n_1832),
.B1(n_1821),
.B2(n_1842),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1893),
.A2(n_1882),
.B1(n_1840),
.B2(n_1737),
.Y(n_2001)
);

INVx8_ASAP7_75t_L g2002 ( 
.A(n_1939),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1893),
.A2(n_1888),
.B1(n_1836),
.B2(n_1820),
.Y(n_2003)
);

BUFx8_ASAP7_75t_L g2004 ( 
.A(n_1927),
.Y(n_2004)
);

CKINVDCx20_ASAP7_75t_R g2005 ( 
.A(n_1950),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1925),
.A2(n_1920),
.B1(n_1902),
.B2(n_1932),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_SL g2007 ( 
.A1(n_1920),
.A2(n_1842),
.B1(n_1874),
.B2(n_1858),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1913),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1902),
.A2(n_1791),
.B1(n_1874),
.B2(n_1779),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1925),
.A2(n_1817),
.B1(n_1858),
.B2(n_1885),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1905),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1895),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1985),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1994),
.A2(n_1791),
.B1(n_1742),
.B2(n_1852),
.Y(n_2014)
);

BUFx8_ASAP7_75t_L g2015 ( 
.A(n_1927),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1979),
.A2(n_1807),
.B1(n_1814),
.B2(n_1879),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1895),
.Y(n_2017)
);

BUFx8_ASAP7_75t_SL g2018 ( 
.A(n_1927),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1992),
.Y(n_2019)
);

OAI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1918),
.A2(n_1851),
.B1(n_1742),
.B2(n_1803),
.Y(n_2020)
);

INVx6_ASAP7_75t_L g2021 ( 
.A(n_1892),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1973),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1973),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1988),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1970),
.B(n_1816),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1988),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_1924),
.Y(n_2027)
);

BUFx12f_ASAP7_75t_L g2028 ( 
.A(n_1910),
.Y(n_2028)
);

BUFx2_ASAP7_75t_SL g2029 ( 
.A(n_1952),
.Y(n_2029)
);

BUFx10_ASAP7_75t_L g2030 ( 
.A(n_1984),
.Y(n_2030)
);

BUFx2_ASAP7_75t_SL g2031 ( 
.A(n_1952),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1972),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1922),
.B(n_1870),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1979),
.A2(n_1872),
.B1(n_1875),
.B2(n_1873),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1968),
.A2(n_1884),
.B1(n_1886),
.B2(n_1862),
.Y(n_2035)
);

CKINVDCx11_ASAP7_75t_R g2036 ( 
.A(n_1911),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1952),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1995),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_1959),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1949),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1949),
.B(n_1838),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1989),
.B(n_1824),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1964),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_SL g2044 ( 
.A1(n_1987),
.A2(n_1762),
.B1(n_1810),
.B2(n_1794),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_1963),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1964),
.B(n_1839),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1995),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1986),
.A2(n_1849),
.B1(n_1853),
.B2(n_1850),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1993),
.A2(n_1851),
.B1(n_1834),
.B2(n_1797),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_1977),
.B(n_1766),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1897),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1908),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1965),
.B(n_1844),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1953),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_1912),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_1957),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1999),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2045),
.B(n_1926),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2008),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_2002),
.Y(n_2060)
);

AOI21x1_ASAP7_75t_L g2061 ( 
.A1(n_2032),
.A2(n_1912),
.B(n_2049),
.Y(n_2061)
);

AND2x4_ASAP7_75t_L g2062 ( 
.A(n_2051),
.B(n_1997),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2012),
.Y(n_2063)
);

OR2x6_ASAP7_75t_L g2064 ( 
.A(n_2029),
.B(n_1996),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2045),
.B(n_1976),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_2055),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_2020),
.A2(n_1916),
.B(n_1901),
.Y(n_2067)
);

OAI221xp5_ASAP7_75t_L g2068 ( 
.A1(n_2000),
.A2(n_1896),
.B1(n_1848),
.B2(n_1804),
.C(n_1795),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2013),
.B(n_1930),
.Y(n_2069)
);

OA21x2_ASAP7_75t_L g2070 ( 
.A1(n_2006),
.A2(n_1954),
.B(n_1909),
.Y(n_2070)
);

AOI21xp33_ASAP7_75t_L g2071 ( 
.A1(n_2007),
.A2(n_1981),
.B(n_1934),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2017),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2013),
.B(n_1975),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2027),
.B(n_1971),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2022),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2040),
.Y(n_2076)
);

A2O1A1Ixp33_ASAP7_75t_L g2077 ( 
.A1(n_2009),
.A2(n_1900),
.B(n_1984),
.C(n_1929),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2010),
.A2(n_1983),
.B1(n_1827),
.B2(n_1981),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_2036),
.Y(n_2079)
);

OA21x2_ASAP7_75t_L g2080 ( 
.A1(n_2023),
.A2(n_1990),
.B(n_1899),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2024),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_2055),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_2026),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2001),
.A2(n_1847),
.B(n_1881),
.Y(n_2084)
);

NAND2x1p5_ASAP7_75t_L g2085 ( 
.A(n_2037),
.B(n_1916),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2043),
.Y(n_2086)
);

BUFx12f_ASAP7_75t_L g2087 ( 
.A(n_2004),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2003),
.A2(n_1916),
.B(n_1901),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_2049),
.A2(n_1919),
.B(n_1946),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2050),
.B(n_1966),
.Y(n_2090)
);

AO31x2_ASAP7_75t_L g2091 ( 
.A1(n_2037),
.A2(n_2047),
.A3(n_2038),
.B(n_2052),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_2034),
.A2(n_1919),
.B(n_1946),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2041),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1998),
.Y(n_2094)
);

AOI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_2033),
.A2(n_1958),
.B(n_1947),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_2068),
.A2(n_2044),
.B1(n_2014),
.B2(n_1917),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2091),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_2078),
.A2(n_1917),
.B1(n_1934),
.B2(n_2048),
.Y(n_2098)
);

AOI322xp5_ASAP7_75t_L g2099 ( 
.A1(n_2078),
.A2(n_1935),
.A3(n_2053),
.B1(n_1854),
.B2(n_1857),
.C1(n_1887),
.C2(n_1878),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_2067),
.A2(n_2016),
.B(n_1877),
.C(n_1876),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_2064),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2084),
.A2(n_1863),
.B1(n_1889),
.B2(n_1883),
.Y(n_2102)
);

AOI221xp5_ASAP7_75t_SL g2103 ( 
.A1(n_2088),
.A2(n_2046),
.B1(n_2041),
.B2(n_2035),
.C(n_2025),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2093),
.B(n_2042),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2093),
.B(n_2011),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_2079),
.Y(n_2106)
);

INVx5_ASAP7_75t_SL g2107 ( 
.A(n_2079),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2083),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2083),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2058),
.B(n_2019),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2057),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_2064),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2066),
.B(n_2082),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_SL g2114 ( 
.A1(n_2089),
.A2(n_1971),
.B1(n_2030),
.B2(n_1958),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2059),
.Y(n_2115)
);

OAI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_2071),
.A2(n_2033),
.B1(n_1907),
.B2(n_1962),
.C(n_1923),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2063),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_SL g2118 ( 
.A1(n_2092),
.A2(n_1971),
.B1(n_2030),
.B2(n_1947),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2077),
.A2(n_1972),
.B1(n_1915),
.B2(n_1991),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2110),
.B(n_2066),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2101),
.B(n_2112),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2108),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2109),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2097),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2104),
.B(n_2073),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2104),
.B(n_2069),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_2106),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2105),
.B(n_2062),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2121),
.B(n_2105),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2124),
.Y(n_2130)
);

INVx6_ASAP7_75t_L g2131 ( 
.A(n_2127),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_2127),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2122),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2123),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_2131),
.B(n_2079),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2129),
.B(n_2121),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2133),
.B(n_2120),
.Y(n_2137)
);

INVx5_ASAP7_75t_L g2138 ( 
.A(n_2132),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2132),
.B(n_2128),
.Y(n_2139)
);

BUFx3_ASAP7_75t_L g2140 ( 
.A(n_2131),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_SL g2141 ( 
.A1(n_2132),
.A2(n_2079),
.B(n_2106),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2134),
.B(n_2125),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_2131),
.B(n_2107),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_2132),
.A2(n_2119),
.B1(n_2096),
.B2(n_2098),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2136),
.B(n_2107),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2137),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2139),
.B(n_2107),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2142),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2138),
.Y(n_2149)
);

OAI211xp5_ASAP7_75t_L g2150 ( 
.A1(n_2144),
.A2(n_2099),
.B(n_2096),
.C(n_2098),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_2138),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2135),
.B(n_2127),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_2138),
.B(n_2143),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2140),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2141),
.B(n_2125),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_2151),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2146),
.B(n_2130),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_2151),
.Y(n_2158)
);

XNOR2xp5_ASAP7_75t_L g2159 ( 
.A(n_2145),
.B(n_2056),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2148),
.Y(n_2160)
);

NAND4xp75_ASAP7_75t_L g2161 ( 
.A(n_2153),
.B(n_2103),
.C(n_2095),
.D(n_1951),
.Y(n_2161)
);

NOR3xp33_ASAP7_75t_SL g2162 ( 
.A(n_2153),
.B(n_2054),
.C(n_2116),
.Y(n_2162)
);

XNOR2xp5_ASAP7_75t_L g2163 ( 
.A(n_2147),
.B(n_2118),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2159),
.B(n_2154),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2158),
.B(n_2154),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2156),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2160),
.B(n_2149),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2164),
.A2(n_2150),
.B(n_2149),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2166),
.B(n_2157),
.Y(n_2169)
);

AOI211xp5_ASAP7_75t_L g2170 ( 
.A1(n_2165),
.A2(n_2157),
.B(n_2155),
.C(n_2163),
.Y(n_2170)
);

OAI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_2167),
.A2(n_2161),
.B(n_2162),
.Y(n_2171)
);

OAI21xp5_ASAP7_75t_SL g2172 ( 
.A1(n_2171),
.A2(n_2152),
.B(n_2114),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2168),
.B(n_2127),
.Y(n_2173)
);

A2O1A1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_2170),
.A2(n_2100),
.B(n_2102),
.C(n_1903),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2169),
.B(n_2126),
.Y(n_2175)
);

INVx1_ASAP7_75t_SL g2176 ( 
.A(n_2169),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2173),
.B(n_2005),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2176),
.B(n_2126),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_2175),
.Y(n_2179)
);

AND2x2_ASAP7_75t_SL g2180 ( 
.A(n_2172),
.B(n_2018),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2174),
.Y(n_2181)
);

AOI221xp5_ASAP7_75t_L g2182 ( 
.A1(n_2176),
.A2(n_2100),
.B1(n_2102),
.B2(n_2130),
.C(n_2077),
.Y(n_2182)
);

OAI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2173),
.A2(n_2021),
.B1(n_2087),
.B2(n_2028),
.Y(n_2183)
);

INVx2_ASAP7_75t_SL g2184 ( 
.A(n_2175),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2173),
.A2(n_2015),
.B1(n_2004),
.B2(n_2021),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_2173),
.B(n_1960),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2178),
.B(n_1931),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2183),
.B(n_1931),
.Y(n_2188)
);

NOR2x1_ASAP7_75t_L g2189 ( 
.A(n_2177),
.B(n_1898),
.Y(n_2189)
);

OAI221xp5_ASAP7_75t_SL g2190 ( 
.A1(n_2181),
.A2(n_2179),
.B1(n_2184),
.B2(n_2185),
.C(n_2182),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2180),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2186),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2183),
.A2(n_1869),
.B(n_1867),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_2183),
.A2(n_1845),
.B(n_1891),
.Y(n_2194)
);

NOR3xp33_ASAP7_75t_L g2195 ( 
.A(n_2183),
.B(n_2060),
.C(n_1771),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_2183),
.B(n_2015),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2178),
.B(n_2111),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_SL g2198 ( 
.A(n_2177),
.B(n_1937),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2179),
.B(n_2113),
.Y(n_2199)
);

OAI32xp33_ASAP7_75t_L g2200 ( 
.A1(n_2187),
.A2(n_2124),
.A3(n_2060),
.B1(n_1978),
.B2(n_1955),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2190),
.A2(n_2064),
.B1(n_2039),
.B2(n_1959),
.Y(n_2201)
);

AOI322xp5_ASAP7_75t_L g2202 ( 
.A1(n_2189),
.A2(n_2097),
.A3(n_2082),
.B1(n_2062),
.B2(n_2128),
.C1(n_2074),
.C2(n_1835),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2199),
.Y(n_2203)
);

OAI21xp33_ASAP7_75t_SL g2204 ( 
.A1(n_2196),
.A2(n_2117),
.B(n_2115),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_2188),
.A2(n_2061),
.B(n_1948),
.Y(n_2205)
);

AOI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2198),
.A2(n_2002),
.B1(n_1865),
.B2(n_1939),
.Y(n_2206)
);

AOI211xp5_ASAP7_75t_L g2207 ( 
.A1(n_2191),
.A2(n_1938),
.B(n_171),
.C(n_169),
.Y(n_2207)
);

O2A1O1Ixp33_ASAP7_75t_SL g2208 ( 
.A1(n_2192),
.A2(n_1859),
.B(n_2065),
.C(n_1880),
.Y(n_2208)
);

NAND2xp33_ASAP7_75t_R g2209 ( 
.A(n_2193),
.B(n_170),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_2195),
.B(n_1969),
.Y(n_2210)
);

OAI221xp5_ASAP7_75t_L g2211 ( 
.A1(n_2197),
.A2(n_2085),
.B1(n_2031),
.B2(n_1936),
.C(n_1944),
.Y(n_2211)
);

AOI322xp5_ASAP7_75t_L g2212 ( 
.A1(n_2194),
.A2(n_2002),
.A3(n_1803),
.B1(n_2090),
.B2(n_1938),
.C1(n_1969),
.C2(n_1945),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2203),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_SL g2214 ( 
.A1(n_2201),
.A2(n_1969),
.B1(n_2085),
.B2(n_1855),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2207),
.Y(n_2215)
);

O2A1O1Ixp33_ASAP7_75t_L g2216 ( 
.A1(n_2210),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2216)
);

OAI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_2204),
.A2(n_1860),
.B1(n_1785),
.B2(n_1841),
.C(n_1856),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_2205),
.A2(n_1982),
.B1(n_1943),
.B2(n_1914),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2208),
.Y(n_2219)
);

O2A1O1Ixp33_ASAP7_75t_SL g2220 ( 
.A1(n_2202),
.A2(n_176),
.B(n_172),
.C(n_175),
.Y(n_2220)
);

A2O1A1Ixp33_ASAP7_75t_SL g2221 ( 
.A1(n_2209),
.A2(n_178),
.B(n_175),
.C(n_177),
.Y(n_2221)
);

AOI22x1_ASAP7_75t_L g2222 ( 
.A1(n_2200),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2206),
.Y(n_2223)
);

OAI22xp33_ASAP7_75t_L g2224 ( 
.A1(n_2211),
.A2(n_2046),
.B1(n_1928),
.B2(n_1933),
.Y(n_2224)
);

AOI211xp5_ASAP7_75t_L g2225 ( 
.A1(n_2213),
.A2(n_2212),
.B(n_182),
.C(n_180),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_L g2226 ( 
.A1(n_2220),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_2226)
);

OAI222xp33_ASAP7_75t_L g2227 ( 
.A1(n_2222),
.A2(n_1945),
.B1(n_1961),
.B2(n_1933),
.C1(n_1928),
.C2(n_2094),
.Y(n_2227)
);

AOI211xp5_ASAP7_75t_L g2228 ( 
.A1(n_2216),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2215),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_2214),
.B(n_2219),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2223),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_R g2232 ( 
.A(n_2221),
.B(n_186),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2224),
.A2(n_1961),
.B1(n_1774),
.B2(n_1982),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2218),
.A2(n_186),
.B(n_187),
.Y(n_2234)
);

NAND5xp2_ASAP7_75t_L g2235 ( 
.A(n_2217),
.B(n_190),
.C(n_188),
.D(n_189),
.E(n_191),
.Y(n_2235)
);

AOI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2220),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_2236)
);

AOI21xp33_ASAP7_75t_SL g2237 ( 
.A1(n_2213),
.A2(n_192),
.B(n_193),
.Y(n_2237)
);

AOI222xp33_ASAP7_75t_L g2238 ( 
.A1(n_2213),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.C1(n_196),
.C2(n_197),
.Y(n_2238)
);

OAI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2213),
.A2(n_1904),
.B1(n_1921),
.B2(n_1908),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2213),
.B(n_194),
.Y(n_2240)
);

AOI221xp5_ASAP7_75t_L g2241 ( 
.A1(n_2231),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.C(n_199),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2229),
.A2(n_1982),
.B1(n_1921),
.B2(n_1940),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2240),
.Y(n_2243)
);

AOI222xp33_ASAP7_75t_L g2244 ( 
.A1(n_2230),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.C1(n_202),
.C2(n_203),
.Y(n_2244)
);

AOI211xp5_ASAP7_75t_L g2245 ( 
.A1(n_2226),
.A2(n_202),
.B(n_200),
.C(n_201),
.Y(n_2245)
);

NOR4xp25_ASAP7_75t_SL g2246 ( 
.A(n_2236),
.B(n_205),
.C(n_203),
.D(n_204),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2233),
.Y(n_2247)
);

OAI211xp5_ASAP7_75t_L g2248 ( 
.A1(n_2232),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_2248)
);

NAND4xp75_ASAP7_75t_L g2249 ( 
.A(n_2234),
.B(n_208),
.C(n_206),
.D(n_207),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2237),
.Y(n_2250)
);

AOI222xp33_ASAP7_75t_L g2251 ( 
.A1(n_2227),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.C1(n_210),
.C2(n_211),
.Y(n_2251)
);

O2A1O1Ixp33_ASAP7_75t_L g2252 ( 
.A1(n_2228),
.A2(n_2225),
.B(n_2235),
.C(n_2238),
.Y(n_2252)
);

O2A1O1Ixp33_ASAP7_75t_L g2253 ( 
.A1(n_2239),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_2253)
);

A2O1A1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_2237),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_2254)
);

NAND2x1p5_ASAP7_75t_SL g2255 ( 
.A(n_2230),
.B(n_212),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2226),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.C(n_217),
.Y(n_2256)
);

INVx2_ASAP7_75t_SL g2257 ( 
.A(n_2240),
.Y(n_2257)
);

NAND3xp33_ASAP7_75t_L g2258 ( 
.A(n_2226),
.B(n_215),
.C(n_217),
.Y(n_2258)
);

OAI21xp5_ASAP7_75t_SL g2259 ( 
.A1(n_2227),
.A2(n_218),
.B(n_219),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2231),
.B(n_218),
.Y(n_2260)
);

NAND4xp25_ASAP7_75t_L g2261 ( 
.A(n_2225),
.B(n_222),
.C(n_220),
.D(n_221),
.Y(n_2261)
);

OAI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2231),
.A2(n_2075),
.B1(n_2081),
.B2(n_2072),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2231),
.A2(n_1982),
.B1(n_1956),
.B2(n_1941),
.Y(n_2263)
);

AOI221xp5_ASAP7_75t_L g2264 ( 
.A1(n_2231),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.C(n_223),
.Y(n_2264)
);

AO22x2_ASAP7_75t_L g2265 ( 
.A1(n_2231),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2265)
);

AOI221xp5_ASAP7_75t_L g2266 ( 
.A1(n_2252),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.C(n_228),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2260),
.Y(n_2267)
);

AO211x2_ASAP7_75t_L g2268 ( 
.A1(n_2261),
.A2(n_229),
.B(n_226),
.C(n_228),
.Y(n_2268)
);

AOI221xp5_ASAP7_75t_L g2269 ( 
.A1(n_2250),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.C(n_234),
.Y(n_2269)
);

OAI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2258),
.A2(n_230),
.B(n_231),
.Y(n_2270)
);

AOI221xp5_ASAP7_75t_L g2271 ( 
.A1(n_2253),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.C(n_237),
.Y(n_2271)
);

NOR2x1_ASAP7_75t_L g2272 ( 
.A(n_2248),
.B(n_237),
.Y(n_2272)
);

NOR3xp33_ASAP7_75t_L g2273 ( 
.A(n_2257),
.B(n_238),
.C(n_239),
.Y(n_2273)
);

O2A1O1Ixp33_ASAP7_75t_L g2274 ( 
.A1(n_2254),
.A2(n_241),
.B(n_238),
.C(n_240),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2265),
.Y(n_2275)
);

A2O1A1Ixp33_ASAP7_75t_L g2276 ( 
.A1(n_2259),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2243),
.B(n_242),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2244),
.B(n_243),
.Y(n_2278)
);

OAI322xp33_ASAP7_75t_L g2279 ( 
.A1(n_2247),
.A2(n_243),
.A3(n_245),
.B1(n_247),
.B2(n_248),
.C1(n_249),
.C2(n_250),
.Y(n_2279)
);

AOI221xp5_ASAP7_75t_L g2280 ( 
.A1(n_2256),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.C(n_250),
.Y(n_2280)
);

NOR2x1_ASAP7_75t_L g2281 ( 
.A(n_2249),
.B(n_251),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2265),
.Y(n_2282)
);

NAND3xp33_ASAP7_75t_SL g2283 ( 
.A(n_2246),
.B(n_2245),
.C(n_2251),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2241),
.B(n_1982),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2282),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2267),
.B(n_2263),
.Y(n_2286)
);

NAND4xp25_ASAP7_75t_L g2287 ( 
.A(n_2276),
.B(n_2264),
.C(n_2255),
.D(n_2242),
.Y(n_2287)
);

NAND4xp75_ASAP7_75t_L g2288 ( 
.A(n_2272),
.B(n_2262),
.C(n_252),
.D(n_253),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_R g2289 ( 
.A(n_2283),
.B(n_251),
.Y(n_2289)
);

NOR3xp33_ASAP7_75t_L g2290 ( 
.A(n_2278),
.B(n_252),
.C(n_254),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2277),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2281),
.B(n_254),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2275),
.A2(n_1956),
.B1(n_1941),
.B2(n_1894),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2273),
.B(n_255),
.Y(n_2294)
);

NAND5xp2_ASAP7_75t_L g2295 ( 
.A(n_2270),
.B(n_255),
.C(n_322),
.D(n_323),
.E(n_324),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2268),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2279),
.B(n_326),
.Y(n_2297)
);

NAND2x1p5_ASAP7_75t_L g2298 ( 
.A(n_2284),
.B(n_1974),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2274),
.B(n_2091),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2280),
.A2(n_1894),
.B1(n_2070),
.B2(n_2076),
.Y(n_2300)
);

A2O1A1Ixp33_ASAP7_75t_L g2301 ( 
.A1(n_2271),
.A2(n_2086),
.B(n_2076),
.C(n_1942),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2266),
.Y(n_2302)
);

AOI32xp33_ASAP7_75t_L g2303 ( 
.A1(n_2269),
.A2(n_2086),
.A3(n_1967),
.B1(n_334),
.B2(n_335),
.Y(n_2303)
);

BUFx2_ASAP7_75t_L g2304 ( 
.A(n_2282),
.Y(n_2304)
);

OAI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2304),
.A2(n_2070),
.B1(n_2080),
.B2(n_1967),
.Y(n_2305)
);

NOR2x1_ASAP7_75t_L g2306 ( 
.A(n_2292),
.B(n_331),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2285),
.B(n_2296),
.Y(n_2307)
);

OA22x2_ASAP7_75t_L g2308 ( 
.A1(n_2291),
.A2(n_333),
.B1(n_336),
.B2(n_337),
.Y(n_2308)
);

NAND5xp2_ASAP7_75t_L g2309 ( 
.A(n_2297),
.B(n_338),
.C(n_339),
.D(n_341),
.E(n_342),
.Y(n_2309)
);

OR3x1_ASAP7_75t_L g2310 ( 
.A(n_2295),
.B(n_345),
.C(n_346),
.Y(n_2310)
);

NAND3xp33_ASAP7_75t_SL g2311 ( 
.A(n_2289),
.B(n_349),
.C(n_350),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2288),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_2286),
.Y(n_2313)
);

NOR3xp33_ASAP7_75t_SL g2314 ( 
.A(n_2302),
.B(n_351),
.C(n_355),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2294),
.B(n_2091),
.Y(n_2315)
);

OAI211xp5_ASAP7_75t_SL g2316 ( 
.A1(n_2290),
.A2(n_2303),
.B(n_2301),
.C(n_2287),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2299),
.A2(n_2298),
.B1(n_2293),
.B2(n_2300),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2295),
.B(n_2091),
.Y(n_2318)
);

OR2x2_ASAP7_75t_L g2319 ( 
.A(n_2295),
.B(n_356),
.Y(n_2319)
);

NAND4xp25_ASAP7_75t_L g2320 ( 
.A(n_2297),
.B(n_357),
.C(n_358),
.D(n_360),
.Y(n_2320)
);

AOI21xp33_ASAP7_75t_L g2321 ( 
.A1(n_2307),
.A2(n_2313),
.B(n_2312),
.Y(n_2321)
);

NOR2xp67_ASAP7_75t_L g2322 ( 
.A(n_2309),
.B(n_362),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2319),
.B(n_364),
.Y(n_2323)
);

INVx1_ASAP7_75t_SL g2324 ( 
.A(n_2306),
.Y(n_2324)
);

NAND5xp2_ASAP7_75t_L g2325 ( 
.A(n_2317),
.B(n_365),
.C(n_366),
.D(n_367),
.E(n_370),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2314),
.B(n_2080),
.Y(n_2326)
);

OAI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2320),
.A2(n_2316),
.B1(n_2318),
.B2(n_2315),
.C(n_2311),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2310),
.A2(n_2070),
.B1(n_2080),
.B2(n_376),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2308),
.Y(n_2329)
);

INVx1_ASAP7_75t_SL g2330 ( 
.A(n_2305),
.Y(n_2330)
);

OR4x2_ASAP7_75t_L g2331 ( 
.A(n_2309),
.B(n_372),
.C(n_375),
.D(n_377),
.Y(n_2331)
);

NOR2x1_ASAP7_75t_L g2332 ( 
.A(n_2306),
.B(n_378),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2319),
.Y(n_2333)
);

AOI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2313),
.A2(n_1914),
.B1(n_382),
.B2(n_383),
.Y(n_2334)
);

XNOR2xp5_ASAP7_75t_L g2335 ( 
.A(n_2310),
.B(n_379),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2307),
.B(n_384),
.Y(n_2336)
);

OAI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2336),
.A2(n_387),
.B1(n_389),
.B2(n_392),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2322),
.A2(n_1914),
.B1(n_398),
.B2(n_399),
.Y(n_2338)
);

AO22x2_ASAP7_75t_L g2339 ( 
.A1(n_2324),
.A2(n_393),
.B1(n_400),
.B2(n_401),
.Y(n_2339)
);

AOI31xp33_ASAP7_75t_L g2340 ( 
.A1(n_2335),
.A2(n_404),
.A3(n_407),
.B(n_408),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2323),
.A2(n_410),
.B1(n_413),
.B2(n_415),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2332),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2331),
.Y(n_2343)
);

AO22x2_ASAP7_75t_L g2344 ( 
.A1(n_2329),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_2344)
);

OAI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2327),
.A2(n_420),
.B1(n_422),
.B2(n_424),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2333),
.A2(n_425),
.B1(n_428),
.B2(n_429),
.Y(n_2346)
);

OAI31xp33_ASAP7_75t_SL g2347 ( 
.A1(n_2342),
.A2(n_2321),
.A3(n_2330),
.B(n_2328),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2344),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2343),
.A2(n_2326),
.B1(n_2334),
.B2(n_2325),
.Y(n_2349)
);

OAI22xp5_ASAP7_75t_SL g2350 ( 
.A1(n_2338),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_2350)
);

AOI22x1_ASAP7_75t_L g2351 ( 
.A1(n_2339),
.A2(n_433),
.B1(n_434),
.B2(n_436),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2340),
.B(n_438),
.Y(n_2352)
);

AOI31xp33_ASAP7_75t_L g2353 ( 
.A1(n_2345),
.A2(n_439),
.A3(n_441),
.B(n_442),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_2351),
.A2(n_2348),
.B1(n_2350),
.B2(n_2352),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2347),
.A2(n_2341),
.B(n_2346),
.C(n_2337),
.Y(n_2355)
);

NOR4xp25_ASAP7_75t_L g2356 ( 
.A(n_2353),
.B(n_2349),
.C(n_444),
.D(n_446),
.Y(n_2356)
);

OR5x1_ASAP7_75t_L g2357 ( 
.A(n_2347),
.B(n_443),
.C(n_449),
.D(n_450),
.E(n_454),
.Y(n_2357)
);

AOI31xp33_ASAP7_75t_L g2358 ( 
.A1(n_2354),
.A2(n_455),
.A3(n_456),
.B(n_457),
.Y(n_2358)
);

AOI22xp33_ASAP7_75t_L g2359 ( 
.A1(n_2357),
.A2(n_1914),
.B1(n_459),
.B2(n_460),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2356),
.A2(n_2355),
.B1(n_1914),
.B2(n_463),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2360),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2358),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_SL g2363 ( 
.A1(n_2362),
.A2(n_2359),
.B(n_461),
.Y(n_2363)
);

NAND3xp33_ASAP7_75t_L g2364 ( 
.A(n_2363),
.B(n_2361),
.C(n_464),
.Y(n_2364)
);

XNOR2xp5_ASAP7_75t_L g2365 ( 
.A(n_2364),
.B(n_458),
.Y(n_2365)
);

OA21x2_ASAP7_75t_L g2366 ( 
.A1(n_2365),
.A2(n_467),
.B(n_468),
.Y(n_2366)
);

OR2x6_ASAP7_75t_L g2367 ( 
.A(n_2365),
.B(n_469),
.Y(n_2367)
);

AOI221xp5_ASAP7_75t_L g2368 ( 
.A1(n_2367),
.A2(n_470),
.B1(n_472),
.B2(n_474),
.C(n_475),
.Y(n_2368)
);

AOI211xp5_ASAP7_75t_L g2369 ( 
.A1(n_2368),
.A2(n_2366),
.B(n_476),
.C(n_477),
.Y(n_2369)
);


endmodule