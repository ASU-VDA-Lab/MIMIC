module fake_jpeg_2676_n_192 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_80),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_53),
.B1(n_46),
.B2(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_70),
.B1(n_65),
.B2(n_63),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_45),
.C(n_53),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_62),
.Y(n_93)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_92),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_68),
.B(n_71),
.C(n_57),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_36),
.B(n_31),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_65),
.B1(n_70),
.B2(n_63),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_77),
.B(n_59),
.C(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_96),
.B1(n_74),
.B2(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_44),
.B1(n_51),
.B2(n_60),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_74),
.B1(n_52),
.B2(n_55),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_49),
.B1(n_47),
.B2(n_61),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_77),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_121),
.B(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_88),
.B1(n_87),
.B2(n_4),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_131),
.B1(n_135),
.B2(n_15),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_88),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_11),
.C(n_13),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_26),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_5),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_6),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_110),
.B(n_10),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_153),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_24),
.B(n_23),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_17),
.C(n_18),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_158),
.B1(n_131),
.B2(n_135),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_8),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_159),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_22),
.B(n_12),
.C(n_13),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_152),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_141),
.B1(n_132),
.B2(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_130),
.B1(n_137),
.B2(n_127),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_16),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_16),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_163),
.B1(n_169),
.B2(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_21),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_18),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_150),
.B1(n_142),
.B2(n_144),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_153),
.C(n_149),
.Y(n_171)
);

XOR2x1_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_162),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_154),
.B(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_175),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_156),
.B1(n_164),
.B2(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_181),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_151),
.B1(n_159),
.B2(n_167),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_172),
.C(n_177),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_180),
.B(n_162),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_184),
.B(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_176),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_177),
.C(n_19),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_19),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_20),
.Y(n_192)
);


endmodule