module real_jpeg_27024_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_0),
.A2(n_105),
.B(n_118),
.Y(n_117)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_0),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_76),
.B1(n_77),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_1),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_85),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_85),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_1),
.A2(n_25),
.B1(n_28),
.B2(n_85),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_3),
.B(n_63),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_3),
.A2(n_63),
.B(n_131),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_11),
.B(n_25),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_42),
.B1(n_49),
.B2(n_184),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_5),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_71),
.Y(n_176)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_56),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_105)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_73),
.Y(n_168)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_106),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_35),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_24),
.A2(n_37),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_24),
.A2(n_37),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_24),
.A2(n_37),
.B1(n_138),
.B2(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_24),
.B(n_78),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_27),
.A2(n_32),
.B(n_78),
.C(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_28),
.B(n_188),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_31),
.A2(n_64),
.A3(n_68),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_32),
.B(n_69),
.Y(n_132)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_54),
.B(n_57),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_37),
.A2(n_139),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_47),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_42),
.B(n_50),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_42),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_42),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_42),
.A2(n_171),
.B1(n_176),
.B2(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_43),
.B(n_78),
.Y(n_188)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_48),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.C(n_74),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_55),
.B(n_58),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_61),
.A2(n_67),
.B1(n_70),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_67),
.B1(n_114),
.B2(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_64),
.B1(n_80),
.B2(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_80),
.Y(n_102)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_75),
.B1(n_82),
.B2(n_102),
.Y(n_101)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.CON(n_75),
.SN(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_80),
.Y(n_82)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_93),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_100),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_103),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_107),
.A2(n_108),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.C(n_116),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_199),
.B(n_205),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_150),
.B(n_198),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_140),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_124),
.B(n_140),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.C(n_136),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_125),
.A2(n_126),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_170),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_141),
.B(n_147),
.C(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_192),
.B(n_197),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_172),
.B(n_191),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_160),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_180),
.B(n_190),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_178),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B(n_189),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);


endmodule