module real_jpeg_15266_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_0),
.B(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_0),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_0),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_0),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_0),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_0),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_0),
.B(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_2),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_2),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_3),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_3),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_3),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_4),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_66),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_5),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_5),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_6),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_6),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_6),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_8),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_8),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_8),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_8),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_8),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_8),
.B(n_227),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_8),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_8),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_78),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_9),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_9),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_9),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_9),
.B(n_295),
.Y(n_424)
);

BUFx2_ASAP7_75t_R g444 ( 
.A(n_9),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_10),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_10),
.B(n_210),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_10),
.B(n_66),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_10),
.B(n_246),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_10),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_10),
.B(n_397),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_11),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_12),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_12),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_12),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_12),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_15),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_12),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_13),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_13),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_13),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_13),
.B(n_238),
.Y(n_237)
);

AND2x4_ASAP7_75t_SL g249 ( 
.A(n_13),
.B(n_246),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_13),
.B(n_286),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_14),
.Y(n_240)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_14),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_15),
.B(n_125),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_15),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_15),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_15),
.B(n_66),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_15),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_15),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_15),
.B(n_430),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_215),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_213),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_173),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_21),
.B(n_173),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_95),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.C(n_85),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_24),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_46),
.C(n_52),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_25),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_26),
.B(n_235),
.C(n_237),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_26),
.A2(n_27),
.B1(n_237),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_27),
.B(n_33),
.C(n_40),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_33),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_38),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_39),
.A2(n_40),
.B1(n_51),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_47),
.C(n_51),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_43),
.Y(n_287)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_44),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_101),
.C(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_46),
.B(n_52),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_47),
.B(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_51),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_53),
.B(n_58),
.C(n_63),
.Y(n_168)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_61),
.Y(n_236)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_67),
.B(n_86),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_77),
.C(n_80),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_68),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.C(n_73),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_69),
.B(n_73),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_70),
.B(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_71),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2x1_ASAP7_75t_SL g212 ( 
.A(n_77),
.B(n_81),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_88),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_94),
.C(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_84),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_88),
.B(n_196),
.C(n_200),
.Y(n_195)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_139),
.B1(n_171),
.B2(n_172),
.Y(n_95)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

XNOR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_113),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_123),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_134),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_134),
.Y(n_170)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_142),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_157),
.B1(n_158),
.B2(n_164),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_155),
.Y(n_352)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_156),
.Y(n_334)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_174),
.B(n_176),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_178),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_194),
.C(n_211),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_179),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_192),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_180),
.B(n_183),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_184),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_187),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_188),
.B(n_351),
.C(n_353),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_188),
.A2(n_189),
.B1(n_351),
.B2(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_190),
.Y(n_380)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_194),
.B(n_211),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_203),
.C(n_208),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_195),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_199),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_202),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_209),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_208),
.A2(n_209),
.B1(n_324),
.B2(n_325),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_209),
.B(n_318),
.C(n_324),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AO21x2_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_312),
.B(n_479),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_306),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_262),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_219),
.B(n_262),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_255),
.Y(n_219)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_241),
.C(n_252),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_234),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_223),
.B(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_225),
.A2(n_226),
.B1(n_234),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_226),
.A2(n_331),
.B(n_335),
.Y(n_330)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_234),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_240),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_241),
.A2(n_252),
.B1(n_253),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.C(n_250),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_242),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_243),
.A2(n_245),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_243),
.B(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_244),
.B(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_245),
.Y(n_343)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_247),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_310),
.C(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.C(n_271),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

XOR2x2_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_272),
.B(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_299),
.C(n_303),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_273),
.B(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.C(n_288),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g356 ( 
.A(n_275),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_278),
.B(n_288),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_285),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_289),
.A2(n_293),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_293),
.B(n_421),
.C(n_423),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_293),
.A2(n_348),
.B1(n_423),
.B2(n_424),
.Y(n_434)
);

XOR2x1_ASAP7_75t_L g345 ( 
.A(n_294),
.B(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_303),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_306),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_307),
.B(n_309),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_475),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_366),
.C(n_371),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_358),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_315),
.B(n_358),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_344),
.C(n_356),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_316),
.B(n_473),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_329),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_330),
.C(n_340),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_318),
.B(n_465),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_SL g410 ( 
.A(n_319),
.B(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_319),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_319),
.A2(n_428),
.B1(n_429),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_340),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_342),
.B(n_378),
.C(n_381),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_344),
.B(n_356),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.C(n_354),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_345),
.B(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_350),
.B(n_355),
.Y(n_460)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

XOR2x2_ASAP7_75t_SL g404 ( 
.A(n_353),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_364),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_361),
.C(n_364),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_367),
.Y(n_477)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_470),
.B(n_474),
.Y(n_371)
);

AOI21x1_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_456),
.B(n_469),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_415),
.B(n_455),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_401),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_401),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_385),
.C(n_392),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_385),
.A2(n_386),
.B1(n_392),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_387),
.B(n_391),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

AO22x1_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_396),
.B1(n_399),
.B2(n_400),
.Y(n_392)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_393),
.Y(n_399)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_396),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_399),
.Y(n_408)
);

INVx5_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_407),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_403),
.B(n_404),
.C(n_407),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_410),
.C(n_411),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_425),
.B(n_454),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_420),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_420),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_421),
.A2(n_422),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_435),
.B(n_453),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_432),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_429),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_447),
.B(n_452),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_445),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_445),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_444),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_444),
.B(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_468),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_468),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_461),
.B2(n_462),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_463),
.C(n_467),
.Y(n_471)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_466),
.B2(n_467),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_471),
.B(n_472),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.C(n_478),
.Y(n_475)
);


endmodule