module fake_netlist_6_3470_n_1022 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1022);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1022;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_953;
wire n_448;
wire n_844;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_111),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_69),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_23),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_77),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_63),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_94),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_75),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_82),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_74),
.Y(n_229)
);

BUFx4f_ASAP7_75t_SL g230 ( 
.A(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_154),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_62),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_141),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_43),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_159),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_58),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_44),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_37),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_70),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_29),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_26),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_145),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_88),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_4),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_25),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_72),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_119),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_174),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_113),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_76),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_120),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_123),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_0),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_18),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_10),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_68),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_56),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_33),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_202),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_195),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_197),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_103),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_117),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_90),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_64),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_99),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_104),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_47),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_155),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_146),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_126),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_194),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_45),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_199),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_173),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_84),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_98),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_67),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_177),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_108),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_196),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_110),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_60),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_100),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_151),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_171),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_116),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_131),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_97),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_105),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_13),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_29),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_26),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_42),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_132),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_R g315 ( 
.A(n_232),
.B(n_38),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_247),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_230),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_265),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_227),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_232),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_252),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_254),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_243),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_243),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_218),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_250),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_264),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_250),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_219),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_223),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_268),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_268),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_307),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_0),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_270),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_275),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_308),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_282),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_222),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_217),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_228),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_234),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_226),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_221),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_225),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_298),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_231),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_252),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_233),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_244),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_305),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_248),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_335),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_340),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_341),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_277),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_323),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_292),
.Y(n_385)
);

OAI21x1_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_292),
.B(n_256),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_251),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_333),
.B(n_260),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_R g394 ( 
.A(n_323),
.B(n_305),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_358),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_318),
.B(n_261),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_320),
.B(n_338),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_315),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_338),
.B(n_240),
.Y(n_404)
);

AND3x2_ASAP7_75t_L g405 ( 
.A(n_337),
.B(n_271),
.C(n_269),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_344),
.B(n_281),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_366),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_346),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_326),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_330),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_355),
.B(n_240),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_350),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_350),
.A2(n_290),
.B(n_286),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_361),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_336),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_375),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_388),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_403),
.B(n_418),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

OA22x2_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_311),
.B1(n_310),
.B2(n_291),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_380),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_229),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_296),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_426),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_422),
.B(n_300),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_403),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_395),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_392),
.B(n_408),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_415),
.B(n_392),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_378),
.B(n_224),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_385),
.B(n_235),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_370),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_385),
.B(n_236),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_401),
.Y(n_463)
);

AND3x2_ASAP7_75t_L g464 ( 
.A(n_379),
.B(n_241),
.C(n_240),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_241),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_409),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_412),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_419),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_39),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_387),
.B(n_237),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_370),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_426),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_419),
.B(n_241),
.Y(n_478)
);

INVx4_ASAP7_75t_SL g479 ( 
.A(n_391),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_424),
.B(n_301),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_238),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

NOR2x1p5_ASAP7_75t_L g486 ( 
.A(n_413),
.B(n_224),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_420),
.B(n_312),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_389),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_384),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_422),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_398),
.B(n_301),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_390),
.C(n_424),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_423),
.B(n_40),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_410),
.A2(n_312),
.B1(n_239),
.B2(n_285),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_383),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_430),
.B(n_374),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_501),
.B(n_383),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_489),
.Y(n_506)
);

BUFx8_ASAP7_75t_L g507 ( 
.A(n_500),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_493),
.A2(n_301),
.B1(n_421),
.B2(n_414),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_430),
.B(n_374),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_444),
.B(n_414),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_493),
.A2(n_421),
.B1(n_297),
.B2(n_295),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_430),
.B(n_376),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_376),
.B1(n_377),
.B2(n_342),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_432),
.B(n_377),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_383),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_242),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_482),
.A2(n_396),
.B1(n_412),
.B2(n_288),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_437),
.B(n_246),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_437),
.B(n_255),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_437),
.B(n_257),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_456),
.B(n_455),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_455),
.B(n_258),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_501),
.B(n_471),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_460),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_486),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_449),
.A2(n_299),
.B1(n_262),
.B2(n_267),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

A2O1A1Ixp33_ASAP7_75t_SL g530 ( 
.A1(n_461),
.A2(n_259),
.B(n_313),
.C(n_304),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_471),
.B(n_272),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_502),
.B(n_273),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_484),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_476),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_439),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_274),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_494),
.B(n_276),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_435),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_458),
.B(n_284),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_462),
.B(n_287),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_502),
.B(n_336),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_495),
.B(n_425),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_502),
.B(n_289),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_498),
.B(n_302),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_450),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_429),
.A2(n_342),
.B1(n_352),
.B2(n_347),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_496),
.B(n_339),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_441),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_467),
.B(n_303),
.Y(n_553)
);

O2A1O1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_472),
.A2(n_352),
.B(n_347),
.C(n_343),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_429),
.A2(n_343),
.B1(n_339),
.B2(n_324),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_487),
.B(n_322),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_467),
.B(n_41),
.Y(n_558)
);

CKINVDCx8_ASAP7_75t_R g559 ( 
.A(n_470),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_478),
.A2(n_324),
.B1(n_322),
.B2(n_416),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_478),
.A2(n_416),
.B1(n_3),
.B2(n_5),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_441),
.A2(n_124),
.B1(n_214),
.B2(n_213),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_435),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_461),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_452),
.B(n_2),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_452),
.B(n_6),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_459),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_433),
.B(n_6),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_435),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_480),
.B(n_7),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_481),
.A2(n_48),
.B(n_46),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_454),
.B(n_49),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_478),
.A2(n_128),
.B1(n_212),
.B2(n_210),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_492),
.B(n_50),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_469),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_473),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_454),
.B(n_51),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_492),
.B(n_52),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_492),
.B(n_53),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_473),
.B(n_8),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_496),
.B(n_9),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_473),
.B(n_11),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_485),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_442),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_485),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_559),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_587),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_557),
.B(n_454),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_552),
.B(n_442),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_552),
.B(n_448),
.Y(n_592)
);

CKINVDCx14_ASAP7_75t_R g593 ( 
.A(n_548),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_576),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_587),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_576),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_522),
.B(n_491),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_564),
.B(n_491),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_573),
.A2(n_478),
.B1(n_488),
.B2(n_457),
.Y(n_599)
);

AOI21x1_ASAP7_75t_L g600 ( 
.A1(n_517),
.A2(n_481),
.B(n_443),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_573),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_505),
.Y(n_602)
);

BUFx4f_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_568),
.A2(n_465),
.B(n_466),
.C(n_453),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_576),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_529),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_475),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_536),
.Y(n_609)
);

OR2x2_ASAP7_75t_SL g610 ( 
.A(n_537),
.B(n_500),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_577),
.B(n_463),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_514),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_555),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_506),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_569),
.A2(n_472),
.B1(n_496),
.B2(n_478),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_524),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_525),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_543),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_578),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_578),
.B(n_483),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_550),
.Y(n_621)
);

OAI21xp33_ASAP7_75t_SL g622 ( 
.A1(n_564),
.A2(n_461),
.B(n_474),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_528),
.B(n_586),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_510),
.B(n_470),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_571),
.A2(n_542),
.B1(n_478),
.B2(n_562),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_534),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_533),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_535),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_567),
.B(n_479),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_503),
.B(n_477),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_507),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g633 ( 
.A(n_560),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_579),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_509),
.B(n_477),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_558),
.A2(n_447),
.B1(n_431),
.B2(n_443),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_518),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_551),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_513),
.B(n_472),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_570),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_507),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g642 ( 
.A(n_526),
.B(n_497),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_569),
.A2(n_474),
.B1(n_427),
.B2(n_434),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_544),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_523),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_538),
.B(n_497),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_497),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_SL g649 ( 
.A(n_563),
.B(n_499),
.C(n_464),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_553),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_SL g651 ( 
.A(n_508),
.B(n_561),
.C(n_554),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g652 ( 
.A(n_565),
.B(n_490),
.C(n_445),
.Y(n_652)
);

AND2x6_ASAP7_75t_SL g653 ( 
.A(n_549),
.B(n_12),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_600),
.A2(n_580),
.B(n_575),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_602),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_639),
.A2(n_597),
.B(n_631),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_646),
.B(n_515),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_626),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_650),
.A2(n_554),
.B(n_508),
.C(n_512),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_597),
.B(n_516),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_598),
.A2(n_581),
.B(n_572),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_598),
.A2(n_572),
.B(n_445),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_589),
.A2(n_447),
.B(n_431),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_595),
.A2(n_520),
.B(n_519),
.Y(n_664)
);

AOI21x1_ASAP7_75t_SL g665 ( 
.A1(n_631),
.A2(n_541),
.B(n_540),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_592),
.B(n_591),
.Y(n_666)
);

OA22x2_ASAP7_75t_L g667 ( 
.A1(n_612),
.A2(n_566),
.B1(n_583),
.B2(n_549),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_590),
.B(n_504),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_615),
.A2(n_512),
.B1(n_539),
.B2(n_561),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_614),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_635),
.B(n_591),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_639),
.A2(n_521),
.B(n_532),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_622),
.A2(n_539),
.B(n_582),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_635),
.A2(n_546),
.B(n_545),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_601),
.A2(n_438),
.B(n_530),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_648),
.B(n_544),
.Y(n_676)
);

AO21x1_ASAP7_75t_L g677 ( 
.A1(n_636),
.A2(n_563),
.B(n_584),
.Y(n_677)
);

AO31x2_ASAP7_75t_L g678 ( 
.A1(n_605),
.A2(n_468),
.A3(n_440),
.B(n_427),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_623),
.B(n_527),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_607),
.A2(n_574),
.B(n_468),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_608),
.B(n_633),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_601),
.A2(n_438),
.B(n_583),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_607),
.A2(n_609),
.B(n_604),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_623),
.B(n_527),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_617),
.Y(n_685)
);

AOI21x1_ASAP7_75t_SL g686 ( 
.A1(n_620),
.A2(n_583),
.B(n_479),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_615),
.A2(n_531),
.B(n_434),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_626),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_609),
.A2(n_440),
.B(n_436),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_588),
.Y(n_690)
);

NAND2x1p5_ASAP7_75t_L g691 ( 
.A(n_601),
.B(n_490),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_651),
.A2(n_490),
.B(n_436),
.C(n_428),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_651),
.A2(n_428),
.B(n_438),
.C(n_451),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_647),
.A2(n_479),
.B1(n_438),
.B2(n_428),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_625),
.A2(n_438),
.B(n_451),
.C(n_479),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_618),
.A2(n_134),
.B(n_215),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_628),
.B(n_451),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_594),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_594),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_594),
.Y(n_700)
);

BUFx12f_ASAP7_75t_L g701 ( 
.A(n_653),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_629),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_590),
.B(n_54),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_644),
.A2(n_451),
.B(n_133),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_621),
.A2(n_136),
.B(n_209),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_596),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_640),
.A2(n_130),
.B(n_208),
.Y(n_708)
);

OAI21x1_ASAP7_75t_SL g709 ( 
.A1(n_704),
.A2(n_599),
.B(n_644),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_690),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_680),
.A2(n_634),
.B(n_627),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_669),
.A2(n_645),
.B1(n_637),
.B2(n_613),
.Y(n_712)
);

CKINVDCx11_ASAP7_75t_R g713 ( 
.A(n_701),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_703),
.B(n_601),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_662),
.A2(n_619),
.B(n_638),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_707),
.Y(n_716)
);

AOI221xp5_ASAP7_75t_L g717 ( 
.A1(n_669),
.A2(n_593),
.B1(n_649),
.B2(n_624),
.C(n_616),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_670),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_702),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_664),
.A2(n_619),
.B(n_638),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_663),
.A2(n_619),
.B(n_643),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_679),
.A2(n_616),
.B(n_649),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_683),
.A2(n_619),
.B(n_643),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_679),
.A2(n_652),
.B(n_620),
.Y(n_724)
);

OAI21x1_ASAP7_75t_SL g725 ( 
.A1(n_704),
.A2(n_603),
.B(n_610),
.Y(n_725)
);

AO21x2_ASAP7_75t_L g726 ( 
.A1(n_693),
.A2(n_652),
.B(n_611),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_658),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_656),
.A2(n_603),
.B(n_611),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_666),
.B(n_596),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_655),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_685),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_678),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_707),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_688),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_678),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_660),
.B(n_596),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_671),
.B(n_606),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_665),
.A2(n_689),
.B(n_654),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_667),
.A2(n_681),
.B1(n_657),
.B2(n_684),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_706),
.Y(n_740)
);

OA21x2_ASAP7_75t_L g741 ( 
.A1(n_661),
.A2(n_630),
.B(n_451),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_696),
.A2(n_606),
.B(n_642),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_656),
.A2(n_12),
.B(n_13),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_698),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_660),
.B(n_606),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_706),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_705),
.A2(n_642),
.B(n_138),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_699),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_684),
.A2(n_671),
.B1(n_659),
.B2(n_657),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_668),
.Y(n_750)
);

AOI211x1_ASAP7_75t_L g751 ( 
.A1(n_677),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_708),
.A2(n_137),
.B(n_186),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_674),
.A2(n_624),
.B(n_641),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_707),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

AOI21x1_ASAP7_75t_L g756 ( 
.A1(n_672),
.A2(n_127),
.B(n_206),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_SL g757 ( 
.A1(n_695),
.A2(n_125),
.B(n_205),
.C(n_204),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_697),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_675),
.A2(n_122),
.B(n_203),
.Y(n_759)
);

AOI22x1_ASAP7_75t_L g760 ( 
.A1(n_725),
.A2(n_674),
.B1(n_673),
.B2(n_682),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_717),
.A2(n_667),
.B1(n_676),
.B2(n_673),
.Y(n_761)
);

CKINVDCx14_ASAP7_75t_R g762 ( 
.A(n_713),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_712),
.B(n_668),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_722),
.A2(n_694),
.B1(n_687),
.B2(n_697),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_739),
.A2(n_703),
.B1(n_700),
.B2(n_687),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_714),
.B(n_692),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_718),
.Y(n_767)
);

AOI221xp5_ASAP7_75t_L g768 ( 
.A1(n_749),
.A2(n_632),
.B1(n_691),
.B2(n_16),
.C(n_17),
.Y(n_768)
);

BUFx4_ASAP7_75t_SL g769 ( 
.A(n_733),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_725),
.A2(n_691),
.B1(n_686),
.B2(n_17),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_734),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_709),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_709),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_753),
.A2(n_743),
.B1(n_724),
.B2(n_745),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_728),
.A2(n_20),
.B(n_21),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_716),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_736),
.B(n_22),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_718),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_736),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_745),
.B(n_23),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_727),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_714),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_729),
.B(n_24),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_719),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_729),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_710),
.B(n_55),
.Y(n_786)
);

INVx6_ASAP7_75t_L g787 ( 
.A(n_710),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_SL g788 ( 
.A(n_737),
.B(n_28),
.C(n_30),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_730),
.B(n_31),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_755),
.A2(n_31),
.A3(n_32),
.B(n_33),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_710),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_730),
.B(n_32),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_751),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_731),
.B(n_34),
.Y(n_794)
);

AO21x2_ASAP7_75t_L g795 ( 
.A1(n_738),
.A2(n_755),
.B(n_715),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_757),
.A2(n_758),
.B(n_719),
.C(n_731),
.Y(n_796)
);

CKINVDCx6p67_ASAP7_75t_R g797 ( 
.A(n_710),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_714),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_714),
.B(n_57),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_758),
.A2(n_35),
.B1(n_59),
.B2(n_61),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_750),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_711),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_744),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_716),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_750),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_744),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_743),
.A2(n_201),
.B1(n_86),
.B2(n_87),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_711),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_740),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_726),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_748),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_732),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_726),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_716),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_750),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_SL g816 ( 
.A1(n_751),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_812),
.Y(n_817)
);

AOI222xp33_ASAP7_75t_L g818 ( 
.A1(n_793),
.A2(n_748),
.B1(n_750),
.B2(n_740),
.C1(n_746),
.C2(n_732),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_784),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_768),
.A2(n_726),
.B1(n_740),
.B2(n_746),
.Y(n_820)
);

OAI221xp5_ASAP7_75t_L g821 ( 
.A1(n_775),
.A2(n_740),
.B1(n_746),
.B2(n_743),
.C(n_756),
.Y(n_821)
);

NAND2x1_ASAP7_75t_L g822 ( 
.A(n_787),
.B(n_735),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_761),
.A2(n_746),
.B1(n_754),
.B2(n_733),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_787),
.B(n_735),
.Y(n_824)
);

INVx11_ASAP7_75t_L g825 ( 
.A(n_769),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_771),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_763),
.A2(n_733),
.B1(n_716),
.B2(n_743),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_741),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_781),
.B(n_779),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_760),
.A2(n_738),
.B(n_715),
.Y(n_830)
);

CKINVDCx11_ASAP7_75t_R g831 ( 
.A(n_797),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_811),
.A2(n_716),
.B1(n_756),
.B2(n_741),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_816),
.A2(n_759),
.B1(n_741),
.B2(n_752),
.Y(n_833)
);

OAI221xp5_ASAP7_75t_L g834 ( 
.A1(n_772),
.A2(n_773),
.B1(n_785),
.B2(n_788),
.C(n_770),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_782),
.A2(n_741),
.B1(n_759),
.B2(n_742),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_764),
.B(n_720),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_766),
.A2(n_752),
.B1(n_742),
.B2(n_747),
.Y(n_837)
);

OAI211xp5_ASAP7_75t_L g838 ( 
.A1(n_788),
.A2(n_807),
.B(n_777),
.C(n_780),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_767),
.B(n_720),
.Y(n_839)
);

OAI22xp33_ASAP7_75t_L g840 ( 
.A1(n_783),
.A2(n_765),
.B1(n_791),
.B2(n_800),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_778),
.B(n_747),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_790),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_766),
.A2(n_723),
.B1(n_721),
.B2(n_102),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_798),
.A2(n_723),
.B1(n_721),
.B2(n_107),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_803),
.A2(n_96),
.B1(n_101),
.B2(n_109),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_802),
.A2(n_114),
.B(n_115),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_798),
.A2(n_118),
.B1(n_129),
.B2(n_139),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_774),
.B(n_140),
.Y(n_848)
);

OA21x2_ASAP7_75t_L g849 ( 
.A1(n_808),
.A2(n_142),
.B(n_143),
.Y(n_849)
);

OA21x2_ASAP7_75t_L g850 ( 
.A1(n_807),
.A2(n_144),
.B(n_147),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_810),
.A2(n_148),
.B(n_150),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_799),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_796),
.A2(n_158),
.B(n_160),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_790),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_809),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_787),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_774),
.B(n_161),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_799),
.A2(n_786),
.B1(n_805),
.B2(n_815),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_790),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_776),
.Y(n_860)
);

OAI221xp5_ASAP7_75t_SL g861 ( 
.A1(n_801),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.C(n_165),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_SL g862 ( 
.A1(n_762),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.C(n_169),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_824),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_828),
.B(n_813),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_828),
.B(n_813),
.Y(n_866)
);

AOI211xp5_ASAP7_75t_L g867 ( 
.A1(n_834),
.A2(n_862),
.B(n_838),
.C(n_861),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_842),
.B(n_810),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_854),
.B(n_795),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_839),
.B(n_795),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_818),
.A2(n_764),
.B1(n_794),
.B2(n_792),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_840),
.B(n_789),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_824),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_817),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_859),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_856),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_817),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_836),
.A2(n_830),
.B(n_835),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_836),
.B(n_790),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_829),
.B(n_814),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_819),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_841),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_841),
.B(n_848),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_819),
.B(n_796),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_830),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_824),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_848),
.B(n_814),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_857),
.B(n_804),
.Y(n_888)
);

NOR2x1_ASAP7_75t_SL g889 ( 
.A(n_824),
.B(n_804),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_855),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_855),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_827),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_855),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_849),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_856),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_857),
.A2(n_850),
.B1(n_858),
.B2(n_820),
.Y(n_896)
);

OAI211xp5_ASAP7_75t_SL g897 ( 
.A1(n_867),
.A2(n_826),
.B(n_831),
.C(n_837),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_883),
.B(n_856),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_872),
.A2(n_850),
.B1(n_821),
.B2(n_823),
.Y(n_899)
);

INVx5_ASAP7_75t_L g900 ( 
.A(n_894),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_SL g901 ( 
.A1(n_872),
.A2(n_850),
.B1(n_856),
.B2(n_831),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_874),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_876),
.Y(n_903)
);

AO21x1_ASAP7_75t_SL g904 ( 
.A1(n_879),
.A2(n_833),
.B(n_843),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_874),
.Y(n_905)
);

NAND2xp33_ASAP7_75t_R g906 ( 
.A(n_880),
.B(n_849),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_863),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_R g908 ( 
.A(n_880),
.B(n_849),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_895),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_880),
.B(n_883),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_883),
.B(n_856),
.Y(n_911)
);

AOI21xp33_ASAP7_75t_L g912 ( 
.A1(n_867),
.A2(n_846),
.B(n_853),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_SL g913 ( 
.A1(n_889),
.A2(n_846),
.B1(n_853),
.B2(n_845),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_874),
.Y(n_914)
);

AOI221xp5_ASAP7_75t_L g915 ( 
.A1(n_892),
.A2(n_806),
.B1(n_832),
.B2(n_852),
.C(n_847),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_910),
.B(n_863),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_907),
.B(n_882),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_898),
.B(n_892),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_901),
.B(n_896),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_897),
.A2(n_896),
.B1(n_871),
.B2(n_888),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_902),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_906),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_911),
.B(n_866),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_905),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_914),
.B(n_882),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_899),
.B(n_866),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_909),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_908),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_900),
.B(n_863),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_900),
.B(n_882),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_900),
.B(n_863),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_924),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_922),
.B(n_882),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_921),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_928),
.B(n_870),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_924),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_931),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_925),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_925),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_935),
.B(n_917),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_938),
.B(n_926),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_934),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_933),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_934),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_933),
.B(n_918),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_935),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_936),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_932),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_SL g949 ( 
.A1(n_946),
.A2(n_919),
.B1(n_889),
.B2(n_937),
.Y(n_949)
);

OAI221xp5_ASAP7_75t_SL g950 ( 
.A1(n_943),
.A2(n_920),
.B1(n_871),
.B2(n_915),
.C(n_919),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_944),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_942),
.Y(n_952)
);

AOI221xp5_ASAP7_75t_L g953 ( 
.A1(n_950),
.A2(n_951),
.B1(n_949),
.B2(n_952),
.C(n_942),
.Y(n_953)
);

OAI32xp33_ASAP7_75t_L g954 ( 
.A1(n_951),
.A2(n_941),
.A3(n_937),
.B1(n_945),
.B2(n_879),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_952),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_949),
.B(n_940),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_955),
.Y(n_957)
);

INVxp33_ASAP7_75t_L g958 ( 
.A(n_956),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_953),
.A2(n_941),
.B(n_947),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_954),
.Y(n_960)
);

OAI211xp5_ASAP7_75t_L g961 ( 
.A1(n_953),
.A2(n_912),
.B(n_913),
.C(n_948),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_957),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_958),
.B(n_940),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_959),
.B(n_937),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_961),
.B(n_912),
.C(n_927),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_958),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_961),
.A2(n_903),
.B1(n_878),
.B2(n_939),
.Y(n_968)
);

OAI221xp5_ASAP7_75t_L g969 ( 
.A1(n_961),
.A2(n_879),
.B1(n_932),
.B2(n_929),
.C(n_931),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_967),
.Y(n_970)
);

AOI211xp5_ASAP7_75t_L g971 ( 
.A1(n_965),
.A2(n_825),
.B(n_930),
.C(n_888),
.Y(n_971)
);

AOI211xp5_ASAP7_75t_L g972 ( 
.A1(n_966),
.A2(n_825),
.B(n_930),
.C(n_888),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_SL g973 ( 
.A1(n_968),
.A2(n_887),
.B(n_895),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_963),
.B(n_964),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_962),
.B(n_917),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_969),
.A2(n_846),
.B(n_878),
.C(n_894),
.Y(n_976)
);

AOI222xp33_ASAP7_75t_L g977 ( 
.A1(n_967),
.A2(n_900),
.B1(n_894),
.B2(n_887),
.C1(n_884),
.C2(n_876),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_970),
.A2(n_878),
.B1(n_895),
.B2(n_876),
.C(n_887),
.Y(n_978)
);

OAI211xp5_ASAP7_75t_L g979 ( 
.A1(n_972),
.A2(n_851),
.B(n_769),
.C(n_844),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_SL g980 ( 
.A1(n_974),
.A2(n_884),
.B(n_864),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_977),
.B(n_909),
.Y(n_981)
);

NAND4xp75_ASAP7_75t_SL g982 ( 
.A(n_973),
.B(n_904),
.C(n_869),
.D(n_865),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_975),
.Y(n_983)
);

OAI221xp5_ASAP7_75t_L g984 ( 
.A1(n_971),
.A2(n_916),
.B1(n_923),
.B2(n_822),
.C(n_864),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_976),
.B(n_916),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_970),
.Y(n_986)
);

AND4x2_ASAP7_75t_L g987 ( 
.A(n_978),
.B(n_860),
.C(n_776),
.D(n_175),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_986),
.B(n_885),
.C(n_875),
.Y(n_988)
);

NAND5xp2_ASAP7_75t_L g989 ( 
.A(n_980),
.B(n_873),
.C(n_866),
.D(n_865),
.E(n_893),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_885),
.C(n_875),
.Y(n_990)
);

OAI22x1_ASAP7_75t_L g991 ( 
.A1(n_981),
.A2(n_873),
.B1(n_886),
.B2(n_870),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_985),
.B(n_170),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_979),
.B(n_870),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_982),
.Y(n_994)
);

OAI221xp5_ASAP7_75t_SL g995 ( 
.A1(n_984),
.A2(n_886),
.B1(n_868),
.B2(n_885),
.C(n_893),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_L g996 ( 
.A(n_994),
.B(n_995),
.C(n_993),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_990),
.A2(n_868),
.B1(n_870),
.B2(n_860),
.Y(n_997)
);

AOI221x1_ASAP7_75t_L g998 ( 
.A1(n_991),
.A2(n_860),
.B1(n_869),
.B2(n_881),
.C(n_870),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_SL g999 ( 
.A1(n_992),
.A2(n_860),
.B1(n_869),
.B2(n_890),
.Y(n_999)
);

NAND4xp25_ASAP7_75t_L g1000 ( 
.A(n_989),
.B(n_865),
.C(n_868),
.D(n_881),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_988),
.B(n_881),
.C(n_877),
.Y(n_1001)
);

OR3x1_ASAP7_75t_L g1002 ( 
.A(n_987),
.B(n_860),
.C(n_178),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_1002),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_999),
.Y(n_1005)
);

NAND4xp25_ASAP7_75t_L g1006 ( 
.A(n_1000),
.B(n_877),
.C(n_891),
.D(n_890),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_997),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1004),
.A2(n_1001),
.B1(n_998),
.B2(n_878),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1003),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1005),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1007),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_SL g1012 ( 
.A1(n_1011),
.A2(n_1006),
.B1(n_891),
.B2(n_890),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1013),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1012),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_1014),
.A2(n_1009),
.B1(n_1008),
.B2(n_891),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1015),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_1017),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_1016),
.A2(n_877),
.B1(n_179),
.B2(n_180),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1018),
.A2(n_172),
.B1(n_184),
.B2(n_185),
.Y(n_1020)
);

AOI221xp5_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_1019),
.B1(n_188),
.B2(n_189),
.C(n_190),
.Y(n_1021)
);

AOI211xp5_ASAP7_75t_L g1022 ( 
.A1(n_1021),
.A2(n_187),
.B(n_192),
.C(n_193),
.Y(n_1022)
);


endmodule