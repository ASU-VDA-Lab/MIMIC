module real_aes_6690_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g105 ( .A(n_0), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_1), .A2(n_133), .B(n_137), .C(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_2), .A2(n_167), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g509 ( .A(n_3), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_4), .B(n_234), .Y(n_253) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_5), .A2(n_167), .B(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_L g133 ( .A(n_6), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g208 ( .A(n_7), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_8), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_8), .B(n_41), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_9), .A2(n_166), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_10), .B(n_145), .Y(n_220) );
INVx1_ASAP7_75t_L g479 ( .A(n_11), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_12), .B(n_248), .Y(n_534) );
INVx1_ASAP7_75t_L g153 ( .A(n_13), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_14), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g546 ( .A(n_15), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_16), .A2(n_143), .B(n_230), .C(n_232), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_17), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_18), .B(n_497), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_19), .B(n_167), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_20), .B(n_179), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_21), .A2(n_248), .B(n_263), .C(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_22), .B(n_234), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_23), .B(n_145), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_24), .A2(n_175), .B(n_232), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_25), .B(n_145), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_26), .Y(n_184) );
INVx1_ASAP7_75t_L g141 ( .A(n_27), .Y(n_141) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_28), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_29), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_30), .B(n_145), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_31), .A2(n_78), .B1(n_458), .B2(n_740), .C1(n_743), .C2(n_744), .Y(n_457) );
INVx1_ASAP7_75t_L g743 ( .A(n_31), .Y(n_743) );
INVx1_ASAP7_75t_L g173 ( .A(n_32), .Y(n_173) );
INVx1_ASAP7_75t_L g488 ( .A(n_33), .Y(n_488) );
INVx2_ASAP7_75t_L g131 ( .A(n_34), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_35), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_36), .A2(n_248), .B(n_249), .C(n_251), .Y(n_247) );
INVxp67_ASAP7_75t_L g174 ( .A(n_37), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_38), .A2(n_137), .B(n_140), .C(n_148), .Y(n_136) );
CKINVDCx14_ASAP7_75t_R g246 ( .A(n_39), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_40), .A2(n_133), .B(n_137), .C(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g111 ( .A(n_41), .Y(n_111) );
INVx1_ASAP7_75t_L g487 ( .A(n_42), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_43), .A2(n_192), .B(n_206), .C(n_207), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_44), .B(n_145), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_45), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_46), .Y(n_169) );
INVx1_ASAP7_75t_L g261 ( .A(n_47), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_48), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_49), .B(n_167), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_50), .A2(n_137), .B1(n_265), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_51), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_52), .Y(n_506) );
CKINVDCx14_ASAP7_75t_R g204 ( .A(n_53), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_54), .A2(n_206), .B(n_251), .C(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_55), .Y(n_562) );
INVx1_ASAP7_75t_L g476 ( .A(n_56), .Y(n_476) );
INVx1_ASAP7_75t_L g134 ( .A(n_57), .Y(n_134) );
INVx1_ASAP7_75t_L g152 ( .A(n_58), .Y(n_152) );
INVx1_ASAP7_75t_SL g250 ( .A(n_59), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_60), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_61), .B(n_234), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_62), .A2(n_100), .B1(n_112), .B2(n_749), .Y(n_99) );
INVx1_ASAP7_75t_L g187 ( .A(n_63), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_SL g496 ( .A1(n_64), .A2(n_251), .B(n_497), .C(n_498), .Y(n_496) );
INVxp67_ASAP7_75t_L g499 ( .A(n_65), .Y(n_499) );
INVx1_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_67), .A2(n_167), .B(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_68), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_69), .A2(n_167), .B(n_227), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_70), .Y(n_491) );
INVx1_ASAP7_75t_L g556 ( .A(n_71), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_72), .A2(n_166), .B(n_168), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g135 ( .A(n_73), .Y(n_135) );
INVx1_ASAP7_75t_L g228 ( .A(n_74), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_75), .A2(n_133), .B(n_137), .C(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_76), .A2(n_167), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g231 ( .A(n_77), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_79), .B(n_142), .Y(n_522) );
INVx2_ASAP7_75t_L g150 ( .A(n_80), .Y(n_150) );
INVx1_ASAP7_75t_L g219 ( .A(n_81), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_82), .B(n_497), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_83), .A2(n_133), .B(n_137), .C(n_508), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_84), .B(n_105), .C(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g449 ( .A(n_84), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g461 ( .A(n_84), .B(n_451), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_84), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_85), .A2(n_137), .B(n_186), .C(n_194), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_86), .A2(n_119), .B1(n_120), .B2(n_446), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_86), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_87), .B(n_149), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_88), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_89), .A2(n_133), .B(n_137), .C(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_90), .Y(n_538) );
INVx1_ASAP7_75t_L g495 ( .A(n_91), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_92), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_93), .B(n_142), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_94), .B(n_157), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_95), .B(n_157), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g264 ( .A(n_97), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_98), .A2(n_167), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g751 ( .A(n_102), .Y(n_751) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_109), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g451 ( .A(n_105), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_456), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g748 ( .A(n_116), .Y(n_748) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_447), .B(n_453), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_121), .A2(n_459), .B1(n_462), .B2(n_466), .Y(n_458) );
INVx1_ASAP7_75t_L g741 ( .A(n_121), .Y(n_741) );
OR4x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_336), .C(n_383), .D(n_423), .Y(n_121) );
NAND3xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_282), .C(n_311), .Y(n_122) );
AOI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_197), .B(n_235), .C(n_275), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_124), .A2(n_295), .B(n_312), .C(n_316), .Y(n_311) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_159), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_126), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_SL g278 ( .A(n_126), .Y(n_278) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_126), .Y(n_290) );
AND2x4_ASAP7_75t_L g294 ( .A(n_126), .B(n_242), .Y(n_294) );
AND2x2_ASAP7_75t_L g305 ( .A(n_126), .B(n_182), .Y(n_305) );
OR2x2_ASAP7_75t_L g329 ( .A(n_126), .B(n_238), .Y(n_329) );
AND2x2_ASAP7_75t_L g342 ( .A(n_126), .B(n_243), .Y(n_342) );
AND2x2_ASAP7_75t_L g382 ( .A(n_126), .B(n_368), .Y(n_382) );
AND2x2_ASAP7_75t_L g389 ( .A(n_126), .B(n_352), .Y(n_389) );
AND2x2_ASAP7_75t_L g419 ( .A(n_126), .B(n_160), .Y(n_419) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_154), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_135), .B(n_136), .C(n_149), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_128), .A2(n_184), .B(n_185), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_128), .A2(n_216), .B(n_217), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_128), .A2(n_177), .B1(n_485), .B2(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_128), .A2(n_506), .B(n_507), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_128), .A2(n_556), .B(n_557), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
AND2x4_ASAP7_75t_L g167 ( .A(n_129), .B(n_133), .Y(n_167) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g147 ( .A(n_130), .Y(n_147) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
INVx1_ASAP7_75t_L g266 ( .A(n_131), .Y(n_266) );
INVx1_ASAP7_75t_L g139 ( .A(n_132), .Y(n_139) );
INVx3_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
INVx1_ASAP7_75t_L g497 ( .A(n_132), .Y(n_497) );
BUFx3_ASAP7_75t_L g148 ( .A(n_133), .Y(n_148) );
INVx4_ASAP7_75t_SL g177 ( .A(n_133), .Y(n_177) );
INVx5_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx3_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_138), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_144), .C(n_146), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g172 ( .A1(n_142), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_142), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_143), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_143), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_143), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
INVx4_ASAP7_75t_L g248 ( .A(n_145), .Y(n_248) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_147), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_149), .A2(n_202), .B(n_209), .Y(n_201) );
INVx1_ASAP7_75t_L g214 ( .A(n_149), .Y(n_214) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_149), .A2(n_541), .B(n_547), .Y(n_540) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_L g158 ( .A(n_150), .B(n_151), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_156), .A2(n_183), .B(n_195), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_156), .B(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g234 ( .A(n_156), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g524 ( .A(n_156), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_157), .A2(n_493), .B(n_500), .Y(n_492) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_159), .B(n_346), .Y(n_358) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_181), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_160), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g296 ( .A(n_160), .B(n_181), .Y(n_296) );
BUFx3_ASAP7_75t_L g304 ( .A(n_160), .Y(n_304) );
OR2x2_ASAP7_75t_L g325 ( .A(n_160), .B(n_200), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_160), .B(n_346), .Y(n_436) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_165), .B(n_178), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_162), .A2(n_239), .B(n_240), .Y(n_238) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_162), .A2(n_555), .B(n_561), .Y(n_554) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_SL g518 ( .A1(n_163), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_164), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_164), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_164), .A2(n_505), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
BUFx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_177), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_170), .A2(n_177), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g227 ( .A1(n_170), .A2(n_177), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_170), .A2(n_177), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_170), .A2(n_177), .B(n_261), .C(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_170), .A2(n_177), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_170), .A2(n_177), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_170), .A2(n_177), .B(n_543), .C(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_175), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_175), .B(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_175), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g189 ( .A(n_176), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_176), .A2(n_189), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g194 ( .A(n_177), .Y(n_194) );
INVx1_ASAP7_75t_L g240 ( .A(n_178), .Y(n_240) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_180), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_180), .A2(n_530), .B(n_537), .Y(n_529) );
AND2x2_ASAP7_75t_L g241 ( .A(n_181), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g289 ( .A(n_181), .Y(n_289) );
AND2x2_ASAP7_75t_L g352 ( .A(n_181), .B(n_243), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_181), .A2(n_355), .B1(n_357), .B2(n_359), .C(n_360), .Y(n_354) );
AND2x2_ASAP7_75t_L g368 ( .A(n_181), .B(n_238), .Y(n_368) );
AND2x2_ASAP7_75t_L g394 ( .A(n_181), .B(n_278), .Y(n_394) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g274 ( .A(n_182), .B(n_243), .Y(n_274) );
BUFx2_ASAP7_75t_L g408 ( .A(n_182), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_190), .C(n_191), .Y(n_186) );
O2A1O1Ixp5_ASAP7_75t_L g218 ( .A1(n_188), .A2(n_191), .B(n_219), .C(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_191), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_191), .A2(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI32xp33_ASAP7_75t_L g374 ( .A1(n_198), .A2(n_335), .A3(n_349), .B1(n_375), .B2(n_376), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
AND2x2_ASAP7_75t_L g315 ( .A(n_199), .B(n_257), .Y(n_315) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g297 ( .A(n_200), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_200), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g369 ( .A(n_200), .B(n_257), .Y(n_369) );
AND2x2_ASAP7_75t_L g380 ( .A(n_200), .B(n_272), .Y(n_380) );
BUFx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g281 ( .A(n_201), .B(n_258), .Y(n_281) );
AND2x2_ASAP7_75t_L g285 ( .A(n_201), .B(n_258), .Y(n_285) );
AND2x2_ASAP7_75t_L g320 ( .A(n_201), .B(n_271), .Y(n_320) );
AND2x2_ASAP7_75t_L g327 ( .A(n_201), .B(n_223), .Y(n_327) );
OAI211xp5_ASAP7_75t_L g332 ( .A1(n_201), .A2(n_278), .B(n_289), .C(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g386 ( .A(n_201), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_201), .B(n_212), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_210), .B(n_269), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_210), .B(n_285), .Y(n_375) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g280 ( .A(n_211), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
AND2x2_ASAP7_75t_L g272 ( .A(n_212), .B(n_224), .Y(n_272) );
OR2x2_ASAP7_75t_L g287 ( .A(n_212), .B(n_224), .Y(n_287) );
AND2x2_ASAP7_75t_L g310 ( .A(n_212), .B(n_271), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_212), .Y(n_314) );
AND2x2_ASAP7_75t_L g333 ( .A(n_212), .B(n_270), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_212), .A2(n_298), .B1(n_344), .B2(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_212), .B(n_386), .Y(n_410) );
AND2x2_ASAP7_75t_L g425 ( .A(n_212), .B(n_285), .Y(n_425) );
INVx4_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx3_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
AND2x2_ASAP7_75t_L g299 ( .A(n_213), .B(n_224), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_213), .B(n_257), .Y(n_301) );
AND3x2_ASAP7_75t_L g363 ( .A(n_213), .B(n_327), .C(n_364), .Y(n_363) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_214), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_214), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_214), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g398 ( .A(n_223), .B(n_270), .Y(n_398) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g257 ( .A(n_224), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_224), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_224), .B(n_269), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_224), .B(n_310), .C(n_386), .Y(n_438) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_233), .Y(n_224) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_225), .A2(n_244), .B(n_253), .Y(n_243) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_225), .A2(n_259), .B(n_267), .Y(n_258) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_234), .A2(n_474), .B(n_480), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_254), .B1(n_268), .B2(n_273), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_241), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_238), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g350 ( .A(n_238), .Y(n_350) );
OAI31xp33_ASAP7_75t_L g366 ( .A1(n_241), .A2(n_367), .A3(n_368), .B(n_369), .Y(n_366) );
AND2x2_ASAP7_75t_L g391 ( .A(n_241), .B(n_278), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_241), .B(n_304), .Y(n_437) );
AND2x2_ASAP7_75t_L g346 ( .A(n_242), .B(n_278), .Y(n_346) );
AND2x2_ASAP7_75t_L g407 ( .A(n_242), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g277 ( .A(n_243), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g335 ( .A(n_243), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_248), .B(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_252), .Y(n_535) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_255), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_256), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AOI221x1_ASAP7_75t_SL g323 ( .A1(n_257), .A2(n_324), .B1(n_326), .B2(n_328), .C(n_330), .Y(n_323) );
INVx2_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
INVx2_ASAP7_75t_L g511 ( .A(n_265), .Y(n_511) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g353 ( .A(n_268), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_269), .B(n_286), .Y(n_378) );
INVx1_ASAP7_75t_SL g441 ( .A(n_269), .Y(n_441) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g359 ( .A(n_272), .B(n_285), .Y(n_359) );
INVx1_ASAP7_75t_L g427 ( .A(n_273), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_273), .B(n_356), .Y(n_440) );
INVx2_ASAP7_75t_SL g279 ( .A(n_274), .Y(n_279) );
AND2x2_ASAP7_75t_L g322 ( .A(n_274), .B(n_278), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_274), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_274), .B(n_349), .Y(n_376) );
AOI21xp33_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_279), .B(n_280), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_277), .B(n_349), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_277), .B(n_304), .Y(n_445) );
OR2x2_ASAP7_75t_L g317 ( .A(n_278), .B(n_296), .Y(n_317) );
AND2x2_ASAP7_75t_L g416 ( .A(n_278), .B(n_407), .Y(n_416) );
OAI22xp5_ASAP7_75t_SL g291 ( .A1(n_279), .A2(n_292), .B1(n_297), .B2(n_300), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_279), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g339 ( .A(n_281), .B(n_287), .Y(n_339) );
INVx1_ASAP7_75t_L g403 ( .A(n_281), .Y(n_403) );
AOI311xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_288), .A3(n_290), .B(n_291), .C(n_302), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_286), .A2(n_418), .B1(n_430), .B2(n_433), .C(n_435), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_286), .B(n_441), .Y(n_443) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g340 ( .A(n_288), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g330 ( .A1(n_289), .A2(n_331), .B(n_332), .C(n_334), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_SL g399 ( .A1(n_293), .A2(n_295), .B(n_400), .C(n_401), .Y(n_399) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_294), .B(n_368), .Y(n_434) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_297), .A2(n_317), .B1(n_318), .B2(n_321), .C(n_323), .Y(n_316) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g319 ( .A(n_299), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g402 ( .A(n_299), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g360 ( .A1(n_303), .A2(n_361), .B(n_362), .C(n_366), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_304), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_304), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g326 ( .A(n_310), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_314), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g428 ( .A(n_317), .Y(n_428) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_320), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g355 ( .A(n_320), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g432 ( .A(n_320), .Y(n_432) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g373 ( .A(n_322), .B(n_349), .Y(n_373) );
INVx1_ASAP7_75t_SL g367 ( .A(n_329), .Y(n_367) );
INVx1_ASAP7_75t_L g344 ( .A(n_335), .Y(n_344) );
NAND3xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_354), .C(n_370), .Y(n_336) );
AOI322xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .A3(n_341), .B1(n_343), .B2(n_347), .C1(n_351), .C2(n_353), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g390 ( .A1(n_338), .A2(n_391), .B(n_392), .C(n_399), .Y(n_390) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_341), .A2(n_362), .B1(n_393), .B2(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g351 ( .A(n_349), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g388 ( .A(n_349), .B(n_389), .Y(n_388) );
AOI32xp33_ASAP7_75t_L g439 ( .A1(n_349), .A2(n_440), .A3(n_441), .B1(n_442), .B2(n_444), .Y(n_439) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g361 ( .A(n_352), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_352), .A2(n_405), .B1(n_409), .B2(n_411), .C(n_414), .Y(n_404) );
AND2x2_ASAP7_75t_L g418 ( .A(n_352), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g421 ( .A(n_356), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g431 ( .A(n_356), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g422 ( .A(n_365), .B(n_386), .Y(n_422) );
AOI211xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B(n_374), .C(n_377), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_387), .B(n_390), .C(n_404), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_398), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g413 ( .A(n_410), .Y(n_413) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B(n_420), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI211xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_426), .B(n_429), .C(n_439), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g455 ( .A(n_449), .Y(n_455) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_450), .B(n_465), .Y(n_746) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g464 ( .A(n_451), .B(n_465), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_453), .A2(n_457), .B(n_747), .Y(n_456) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22x1_ASAP7_75t_L g740 ( .A1(n_459), .A2(n_462), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g742 ( .A(n_467), .Y(n_742) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND3x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_662), .C(n_707), .Y(n_468) );
NOR4xp25_ASAP7_75t_L g469 ( .A(n_470), .B(n_585), .C(n_626), .D(n_643), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_501), .B(n_515), .C(n_548), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_472), .B(n_502), .Y(n_501) );
NOR4xp25_ASAP7_75t_L g609 ( .A(n_472), .B(n_603), .C(n_610), .D(n_616), .Y(n_609) );
AND2x2_ASAP7_75t_L g682 ( .A(n_472), .B(n_571), .Y(n_682) );
AND2x2_ASAP7_75t_L g701 ( .A(n_472), .B(n_647), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_472), .B(n_696), .Y(n_710) );
AND2x2_ASAP7_75t_L g723 ( .A(n_472), .B(n_514), .Y(n_723) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_SL g568 ( .A(n_473), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_473), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g625 ( .A(n_473), .B(n_482), .Y(n_625) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_473), .B(n_571), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_473), .B(n_482), .Y(n_640) );
AND2x2_ASAP7_75t_L g649 ( .A(n_473), .B(n_574), .Y(n_649) );
BUFx2_ASAP7_75t_L g672 ( .A(n_473), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_473), .B(n_492), .Y(n_676) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
AND2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_492), .Y(n_514) );
BUFx2_ASAP7_75t_L g578 ( .A(n_482), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_482), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_610) );
OR2x2_ASAP7_75t_L g632 ( .A(n_482), .B(n_504), .Y(n_632) );
AND2x2_ASAP7_75t_L g696 ( .A(n_482), .B(n_574), .Y(n_696) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g564 ( .A(n_483), .B(n_504), .Y(n_564) );
AND2x2_ASAP7_75t_L g571 ( .A(n_483), .B(n_492), .Y(n_571) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_483), .Y(n_613) );
OR2x2_ASAP7_75t_L g648 ( .A(n_483), .B(n_503), .Y(n_648) );
INVx1_ASAP7_75t_L g567 ( .A(n_492), .Y(n_567) );
INVx3_ASAP7_75t_L g576 ( .A(n_492), .Y(n_576) );
BUFx2_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
AND2x2_ASAP7_75t_L g633 ( .A(n_492), .B(n_568), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_501), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_503), .B(n_576), .Y(n_580) );
INVx1_ASAP7_75t_L g608 ( .A(n_503), .Y(n_608) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
INVx1_ASAP7_75t_L g586 ( .A(n_514), .Y(n_586) );
NAND2x1_ASAP7_75t_SL g515 ( .A(n_516), .B(n_526), .Y(n_515) );
AND2x2_ASAP7_75t_L g584 ( .A(n_516), .B(n_539), .Y(n_584) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_516), .Y(n_658) );
AND2x2_ASAP7_75t_L g685 ( .A(n_516), .B(n_605), .Y(n_685) );
AND2x2_ASAP7_75t_L g693 ( .A(n_516), .B(n_655), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_516), .B(n_551), .Y(n_720) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g552 ( .A(n_517), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g569 ( .A(n_517), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g590 ( .A(n_517), .Y(n_590) );
INVx1_ASAP7_75t_L g596 ( .A(n_517), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_517), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g629 ( .A(n_517), .B(n_554), .Y(n_629) );
OR2x2_ASAP7_75t_L g667 ( .A(n_517), .B(n_622), .Y(n_667) );
AOI32xp33_ASAP7_75t_L g679 ( .A1(n_517), .A2(n_680), .A3(n_683), .B1(n_684), .B2(n_685), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_517), .B(n_655), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_517), .B(n_615), .Y(n_730) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g641 ( .A(n_527), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
INVx1_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
AND2x2_ASAP7_75t_L g605 ( .A(n_528), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_528), .B(n_553), .Y(n_622) );
AND2x2_ASAP7_75t_L g655 ( .A(n_528), .B(n_631), .Y(n_655) );
AND2x2_ASAP7_75t_L g692 ( .A(n_528), .B(n_554), .Y(n_692) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g551 ( .A(n_529), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_529), .B(n_553), .Y(n_582) );
AND2x2_ASAP7_75t_L g589 ( .A(n_529), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g630 ( .A(n_529), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_539), .B(n_553), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_539), .B(n_597), .Y(n_678) );
INVx1_ASAP7_75t_L g700 ( .A(n_539), .Y(n_700) );
INVx1_ASAP7_75t_L g717 ( .A(n_539), .Y(n_717) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g570 ( .A(n_540), .B(n_553), .Y(n_570) );
AND2x2_ASAP7_75t_L g592 ( .A(n_540), .B(n_554), .Y(n_592) );
INVx1_ASAP7_75t_L g631 ( .A(n_540), .Y(n_631) );
AOI221x1_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_563), .B1(n_569), .B2(n_571), .C(n_572), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_549), .A2(n_636), .B1(n_703), .B2(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g594 ( .A(n_550), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g689 ( .A(n_550), .B(n_569), .Y(n_689) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g645 ( .A(n_551), .B(n_570), .Y(n_645) );
INVx1_ASAP7_75t_L g657 ( .A(n_552), .Y(n_657) );
AND2x2_ASAP7_75t_L g668 ( .A(n_552), .B(n_655), .Y(n_668) );
AND2x2_ASAP7_75t_L g735 ( .A(n_552), .B(n_630), .Y(n_735) );
INVx2_ASAP7_75t_L g597 ( .A(n_553), .Y(n_597) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_564), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g687 ( .A(n_564), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_565), .B(n_648), .Y(n_651) );
INVx3_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_566), .A2(n_687), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_SL g709 ( .A(n_569), .B(n_595), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_570), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g661 ( .A(n_570), .B(n_589), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_570), .B(n_596), .Y(n_738) );
AND2x2_ASAP7_75t_L g607 ( .A(n_571), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g674 ( .A(n_571), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B(n_581), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_574), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g623 ( .A(n_574), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g635 ( .A(n_574), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_574), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g659 ( .A(n_575), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_575), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_575), .B(n_578), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_578), .A2(n_617), .B(n_647), .C(n_649), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_578), .A2(n_665), .B1(n_668), .B2(n_669), .C(n_673), .Y(n_664) );
AND2x2_ASAP7_75t_L g660 ( .A(n_579), .B(n_613), .Y(n_660) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g620 ( .A(n_584), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g691 ( .A(n_584), .B(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_593), .C(n_618), .Y(n_585) );
NAND3xp33_ASAP7_75t_SL g704 ( .A(n_586), .B(n_705), .C(n_706), .Y(n_704) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
OR2x2_ASAP7_75t_L g677 ( .A(n_588), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_601), .B2(n_607), .C(n_609), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_595), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_595), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g617 ( .A(n_600), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_600), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
OR2x2_ASAP7_75t_L g737 ( .A(n_600), .B(n_648), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVxp67_ASAP7_75t_L g711 ( .A(n_603), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_605), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g612 ( .A(n_606), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_608), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_608), .B(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_608), .B(n_675), .Y(n_714) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_612), .Y(n_638) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g728 ( .A(n_617), .B(n_648), .Y(n_728) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g706 ( .A(n_623), .Y(n_706) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI322xp33_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_632), .A3(n_633), .B1(n_634), .B2(n_637), .C1(n_639), .C2(n_641), .Y(n_626) );
OAI322xp33_ASAP7_75t_L g708 ( .A1(n_627), .A2(n_709), .A3(n_710), .B1(n_711), .B2(n_712), .C1(n_713), .C2(n_715), .Y(n_708) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx4_ASAP7_75t_L g642 ( .A(n_629), .Y(n_642) );
AND2x2_ASAP7_75t_L g703 ( .A(n_629), .B(n_655), .Y(n_703) );
AND2x2_ASAP7_75t_L g716 ( .A(n_629), .B(n_717), .Y(n_716) );
CKINVDCx16_ASAP7_75t_R g727 ( .A(n_632), .Y(n_727) );
INVx1_ASAP7_75t_L g705 ( .A(n_633), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_635), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g722 ( .A(n_635), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_635), .B(n_676), .Y(n_733) );
OR2x2_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
INVxp33_ASAP7_75t_L g683 ( .A(n_638), .Y(n_683) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_642), .A2(n_644), .B1(n_646), .B2(n_650), .C(n_652), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g699 ( .A(n_642), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g726 ( .A(n_642), .Y(n_726) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_649), .A2(n_674), .A3(n_691), .B1(n_693), .B2(n_694), .C1(n_697), .C2(n_701), .Y(n_690) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_660), .B2(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_686), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_679), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_667), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NAND2xp33_ASAP7_75t_SL g684 ( .A(n_670), .B(n_681), .Y(n_684) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g724 ( .A1(n_672), .A2(n_725), .A3(n_727), .B1(n_728), .B2(n_729), .C1(n_731), .C2(n_734), .Y(n_724) );
AOI21xp33_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_682), .B(n_730), .Y(n_739) );
OAI211xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_688), .B(n_690), .C(n_702), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_718), .C(n_724), .D(n_736), .Y(n_707) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx14_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
OAI21xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_738), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
endmodule