module real_jpeg_14064_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_33),
.B1(n_52),
.B2(n_56),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_68),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_5),
.A2(n_52),
.B1(n_56),
.B2(n_68),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_5),
.A2(n_25),
.B1(n_31),
.B2(n_68),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_52),
.B1(n_56),
.B2(n_70),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_25),
.B1(n_31),
.B2(n_70),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_36),
.B(n_37),
.C(n_43),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_8),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_8),
.B(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_40),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_40),
.B(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_8),
.B(n_25),
.C(n_86),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_39),
.B1(n_52),
.B2(n_56),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_8),
.A2(n_24),
.B1(n_27),
.B2(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_8),
.B(n_62),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_49),
.B1(n_52),
.B2(n_56),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_9),
.A2(n_25),
.B1(n_31),
.B2(n_49),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_30),
.B1(n_52),
.B2(n_56),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_13),
.A2(n_25),
.B1(n_31),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_13),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_52),
.B1(n_56),
.B2(n_80),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_14),
.A2(n_25),
.B1(n_31),
.B2(n_61),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_14),
.A2(n_52),
.B1(n_56),
.B2(n_61),
.Y(n_118)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_110),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_47),
.C(n_63),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_21),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_34),
.B1(n_35),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_22),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_23),
.A2(n_77),
.B(n_98),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_23),
.A2(n_28),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_24),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_24),
.A2(n_27),
.B1(n_191),
.B2(n_199),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_24),
.A2(n_76),
.B(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_25),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_25),
.A2(n_31),
.B1(n_86),
.B2(n_87),
.Y(n_89)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_27),
.B(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_27),
.B(n_39),
.Y(n_197)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_28),
.B(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_28),
.A2(n_29),
.B(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_31),
.B(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B(n_40),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_39),
.B(n_89),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_57)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_SL g163 ( 
.A(n_41),
.B(n_54),
.C(n_56),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_63),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_50),
.A2(n_60),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_50),
.A2(n_51),
.B1(n_122),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_50),
.A2(n_51),
.B1(n_146),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_56),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_52),
.A2(n_55),
.B(n_161),
.C(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_52),
.B(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_62),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_65),
.B1(n_69),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_67),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_93),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_81),
.B2(n_92),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_89),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_84),
.A2(n_90),
.B1(n_156),
.B2(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_84),
.A2(n_90),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_84),
.A2(n_90),
.B1(n_178),
.B2(n_188),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_118),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_99),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.C(n_128),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_111),
.B(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_113),
.B(n_128),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.C(n_123),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_119),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_155),
.B(n_157),
.Y(n_154)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_227),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_222),
.B(n_223),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_166),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_151),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_136),
.B(n_151),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_149),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_140),
.B1(n_147),
.B2(n_148),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_140),
.B(n_147),
.C(n_149),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_158),
.B1(n_159),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_164),
.B1(n_165),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_179),
.B(n_221),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_177),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_215),
.B(n_220),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_205),
.B(n_214),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_194),
.B(n_204),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_189),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B(n_203),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_210),
.C(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_226),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);


endmodule