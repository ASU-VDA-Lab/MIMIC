module fake_jpeg_31212_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_52),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_26),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_60),
.Y(n_109)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_63),
.Y(n_160)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_67),
.B(n_72),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_30),
.B(n_6),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_79),
.B(n_83),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_10),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_10),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_88),
.B(n_41),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_100),
.Y(n_139)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_103),
.Y(n_151)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_105),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_27),
.B1(n_63),
.B2(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_106),
.A2(n_122),
.B1(n_152),
.B2(n_47),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_41),
.B(n_24),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_107),
.A2(n_47),
.B(n_48),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_108),
.B(n_115),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_51),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_21),
.B1(n_42),
.B2(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_118),
.A2(n_136),
.B1(n_147),
.B2(n_122),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_53),
.A2(n_94),
.B1(n_70),
.B2(n_68),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_120),
.A2(n_153),
.B1(n_166),
.B2(n_33),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_27),
.B1(n_23),
.B2(n_32),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_52),
.A2(n_51),
.B1(n_49),
.B2(n_36),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_37),
.B(n_39),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_78),
.A2(n_21),
.B1(n_42),
.B2(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_80),
.B(n_49),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_159),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_62),
.A2(n_21),
.B1(n_42),
.B2(n_23),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_23),
.B1(n_21),
.B2(n_42),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_65),
.A2(n_38),
.B1(n_36),
.B2(n_45),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_86),
.A2(n_38),
.B1(n_37),
.B2(n_45),
.Y(n_166)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_169),
.A2(n_170),
.B(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_176),
.Y(n_243)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_87),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_183),
.Y(n_244)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

AO22x2_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_102),
.B1(n_99),
.B2(n_82),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_112),
.Y(n_183)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_188),
.Y(n_251)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_109),
.B(n_40),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_191),
.B(n_192),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_40),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_211),
.B1(n_182),
.B2(n_177),
.Y(n_220)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_208),
.Y(n_218)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_204),
.B1(n_209),
.B2(n_210),
.Y(n_221)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_201),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_39),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_202),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_91),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_203),
.B(n_215),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_154),
.A2(n_75),
.B1(n_110),
.B2(n_140),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_121),
.A2(n_91),
.B(n_89),
.C(n_17),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_207),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_124),
.B1(n_165),
.B2(n_163),
.Y(n_229)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_125),
.A2(n_96),
.B1(n_95),
.B2(n_92),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_136),
.B1(n_116),
.B2(n_118),
.Y(n_224)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_17),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_217),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_150),
.A2(n_106),
.B(n_89),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_149),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_28),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_224),
.A2(n_144),
.B1(n_167),
.B2(n_163),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_229),
.A2(n_179),
.B1(n_167),
.B2(n_165),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_182),
.A2(n_147),
.B(n_157),
.C(n_161),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_232),
.A2(n_236),
.B(n_206),
.C(n_201),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_177),
.A2(n_149),
.B1(n_157),
.B2(n_131),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_177),
.B(n_112),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_170),
.B(n_113),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_246),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_217),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_200),
.B1(n_185),
.B2(n_182),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_256),
.B1(n_279),
.B2(n_221),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_210),
.B1(n_117),
.B2(n_189),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_242),
.C(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_276),
.C(n_284),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_218),
.B(n_199),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_262),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_228),
.A2(n_205),
.B(n_213),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_238),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_184),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_178),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_282),
.B1(n_232),
.B2(n_229),
.Y(n_297)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_171),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_281),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_251),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_275),
.A2(n_234),
.B1(n_144),
.B2(n_253),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_207),
.C(n_208),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_234),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_225),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_244),
.A2(n_183),
.B1(n_181),
.B2(n_168),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_242),
.B(n_227),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_280),
.B(n_223),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_251),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_237),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_180),
.C(n_175),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_187),
.C(n_190),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_228),
.C(n_220),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_174),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_290),
.A2(n_295),
.B1(n_301),
.B2(n_304),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_257),
.B(n_244),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_293),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_224),
.B1(n_232),
.B2(n_219),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_308),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_219),
.B1(n_246),
.B2(n_237),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_219),
.B1(n_231),
.B2(n_243),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_243),
.B1(n_254),
.B2(n_253),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_281),
.A2(n_132),
.B1(n_131),
.B2(n_146),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_231),
.B1(n_132),
.B2(n_146),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_156),
.B1(n_223),
.B2(n_238),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_310),
.A2(n_275),
.B1(n_285),
.B2(n_265),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_253),
.B1(n_156),
.B2(n_250),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_279),
.B1(n_283),
.B2(n_284),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_314),
.B(n_317),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_226),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_283),
.Y(n_321)
);

OR2x6_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_280),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_247),
.C(n_226),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_319),
.B(n_334),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_296),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_328),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_268),
.C(n_262),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_335),
.Y(n_372)
);

BUFx12f_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_325),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_326),
.A2(n_345),
.B1(n_349),
.B2(n_305),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_296),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_283),
.Y(n_330)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_276),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g356 ( 
.A(n_333),
.B(n_316),
.C(n_306),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_267),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_287),
.B(n_263),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_339),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_297),
.A2(n_300),
.B1(n_298),
.B2(n_286),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_344),
.B1(n_252),
.B2(n_235),
.Y(n_376)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_342),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_271),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_343),
.B(n_347),
.Y(n_359)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_270),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_346),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_312),
.B(n_308),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_295),
.A2(n_272),
.B1(n_258),
.B2(n_261),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_351),
.A2(n_367),
.B(n_331),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_314),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_361),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_327),
.A2(n_293),
.B1(n_317),
.B2(n_292),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_375),
.B1(n_376),
.B2(n_345),
.Y(n_384)
);

BUFx12f_ASAP7_75t_SL g400 ( 
.A(n_356),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_292),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_357),
.B(n_333),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_291),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_313),
.C(n_309),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_363),
.B(n_364),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_320),
.B(n_313),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_325),
.A2(n_306),
.B(n_309),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_303),
.C(n_306),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_368),
.B(n_378),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_278),
.B(n_277),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_373),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_374),
.A2(n_381),
.B1(n_362),
.B2(n_354),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_327),
.A2(n_301),
.B1(n_274),
.B2(n_266),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_333),
.B(n_264),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_378),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_247),
.C(n_264),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_348),
.B1(n_339),
.B2(n_318),
.Y(n_380)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_380),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_324),
.A2(n_241),
.B1(n_264),
.B2(n_250),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_384),
.A2(n_388),
.B1(n_374),
.B2(n_385),
.Y(n_412)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_387),
.B(n_403),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_324),
.B1(n_322),
.B2(n_333),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_371),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_399),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_330),
.B(n_325),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_390),
.A2(n_410),
.B(n_245),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_359),
.B(n_346),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_394),
.Y(n_426)
);

XNOR2x1_ASAP7_75t_SL g393 ( 
.A(n_356),
.B(n_333),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_377),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_365),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_235),
.Y(n_396)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_396),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_318),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_329),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_405),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_363),
.B(n_344),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_402),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_338),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_407),
.B1(n_351),
.B2(n_350),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_325),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_337),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_362),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_342),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_409),
.B(n_245),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_412),
.A2(n_415),
.B1(n_421),
.B2(n_394),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_428),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_357),
.C(n_355),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_420),
.C(n_423),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_385),
.A2(n_381),
.B1(n_350),
.B2(n_360),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_432),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_361),
.C(n_353),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_379),
.B1(n_370),
.B2(n_358),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_358),
.C(n_379),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_424),
.Y(n_444)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_427),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_384),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_410),
.A2(n_214),
.B(n_173),
.Y(n_430)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_430),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_233),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_417),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_426),
.B(n_389),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_442),
.Y(n_456)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_445),
.Y(n_468)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_433),
.A2(n_406),
.B1(n_405),
.B2(n_382),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_397),
.B1(n_431),
.B2(n_407),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_387),
.C(n_400),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_448),
.C(n_449),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_428),
.C(n_420),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_388),
.C(n_390),
.Y(n_449)
);

BUFx24_ASAP7_75t_SL g450 ( 
.A(n_434),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_450),
.B(n_451),
.Y(n_460)
);

AOI21xp33_ASAP7_75t_L g451 ( 
.A1(n_422),
.A2(n_391),
.B(n_395),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_452),
.B(n_455),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_401),
.C(n_408),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_454),
.C(n_418),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_391),
.C(n_399),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_462),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_412),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_465),
.Y(n_478)
);

OAI321xp33_ASAP7_75t_L g461 ( 
.A1(n_444),
.A2(n_429),
.A3(n_397),
.B1(n_418),
.B2(n_424),
.C(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_416),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_463),
.B(n_12),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_415),
.C(n_413),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_436),
.C(n_447),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_407),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_467),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_393),
.B(n_217),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_439),
.A2(n_217),
.B(n_241),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_471),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_241),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_435),
.A2(n_250),
.B1(n_233),
.B2(n_212),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_473),
.B1(n_198),
.B2(n_194),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_441),
.A2(n_449),
.B1(n_453),
.B2(n_454),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_475),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_456),
.B(n_193),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_233),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_481),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_482),
.B(n_483),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_463),
.B(n_12),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_134),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_486),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_196),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_470),
.A2(n_28),
.B1(n_12),
.B2(n_4),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_487),
.A2(n_13),
.B(n_15),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_28),
.C(n_196),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_28),
.C(n_19),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_468),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_496),
.Y(n_503)
);

OAI221xp5_ASAP7_75t_L g491 ( 
.A1(n_476),
.A2(n_469),
.B1(n_467),
.B2(n_464),
.C(n_465),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_491),
.A2(n_478),
.B(n_485),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_4),
.Y(n_508)
);

NOR3xp33_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_458),
.C(n_462),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_489),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_499),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_19),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_5),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_19),
.C(n_28),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_488),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_504),
.A2(n_506),
.B(n_510),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_507),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_493),
.A2(n_480),
.B(n_487),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_497),
.A2(n_5),
.B1(n_13),
.B2(n_11),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_509),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_5),
.Y(n_510)
);

NAND4xp25_ASAP7_75t_SL g513 ( 
.A(n_511),
.B(n_496),
.C(n_492),
.D(n_495),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_513),
.B(n_510),
.C(n_498),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_503),
.A2(n_501),
.B(n_500),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_15),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_517),
.A2(n_518),
.B(n_519),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_5),
.C(n_13),
.Y(n_518)
);

OAI311xp33_ASAP7_75t_L g521 ( 
.A1(n_517),
.A2(n_516),
.A3(n_514),
.B1(n_3),
.C1(n_1),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_521),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_520),
.C(n_1),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_3),
.B(n_0),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_0),
.B(n_1),
.Y(n_526)
);


endmodule