module fake_aes_1329_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
NAND3xp33_ASAP7_75t_L g3 ( .A(n_1), .B(n_0), .C(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_0), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_7) );
OR2x6_ASAP7_75t_SL g8 ( .A(n_5), .B(n_0), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_8), .B(n_1), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_1), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_7), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_9), .B(n_3), .Y(n_12) );
OAI322xp33_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_2), .A3(n_3), .B1(n_6), .B2(n_7), .C1(n_10), .C2(n_11), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
A2O1A1Ixp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_2), .B(n_6), .C(n_13), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_2), .B1(n_6), .B2(n_12), .Y(n_16) );
OA21x2_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_2), .B(n_16), .Y(n_17) );
INVxp67_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
endmodule