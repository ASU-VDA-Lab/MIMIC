module fake_jpeg_29880_n_202 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_20),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_28),
.B1(n_11),
.B2(n_9),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_26),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_50),
.Y(n_66)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_64),
.B(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_16),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_30),
.B(n_29),
.C(n_16),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_61),
.B(n_83),
.C(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_30),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_20),
.B1(n_29),
.B2(n_33),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_90),
.B1(n_86),
.B2(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_39),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_28),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_92),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_3),
.C(n_4),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_66),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_117),
.C(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_98),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_91),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_107),
.Y(n_125)
);

NAND2x1p5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_68),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_82),
.B1(n_66),
.B2(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_106),
.B1(n_112),
.B2(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_63),
.B1(n_70),
.B2(n_68),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_118),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_71),
.C(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_71),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_102),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_138),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_95),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_93),
.B1(n_112),
.B2(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_154),
.B1(n_123),
.B2(n_134),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_158),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_116),
.B1(n_104),
.B2(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_152),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_142),
.A2(n_100),
.B1(n_111),
.B2(n_120),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_130),
.B(n_132),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_94),
.B1(n_107),
.B2(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_132),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_146),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_126),
.B1(n_127),
.B2(n_136),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_141),
.B1(n_122),
.B2(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_125),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_147),
.C(n_157),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_149),
.B1(n_145),
.B2(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_178),
.B1(n_179),
.B2(n_167),
.Y(n_183)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_153),
.B1(n_135),
.B2(n_128),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_177),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_163),
.C(n_170),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_182),
.C(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_163),
.C(n_166),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_172),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_171),
.B(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_186),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_173),
.C(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_179),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_175),
.B1(n_176),
.B2(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_139),
.A3(n_174),
.B1(n_176),
.B2(n_177),
.C1(n_182),
.C2(n_195),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_194),
.C(n_174),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_196),
.B(n_139),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule