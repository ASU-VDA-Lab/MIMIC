module real_jpeg_11433_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_63),
.B1(n_65),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_3),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_3),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_71),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_5),
.A2(n_36),
.B1(n_68),
.B2(n_69),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_5),
.A2(n_36),
.B1(n_63),
.B2(n_65),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_6),
.A2(n_63),
.B1(n_65),
.B2(n_82),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_82),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_129),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_7),
.B(n_30),
.C(n_46),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_104),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_27),
.B1(n_33),
.B2(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_7),
.B(n_110),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_11),
.A2(n_63),
.B1(n_65),
.B2(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_73),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_12),
.A2(n_63),
.B1(n_65),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_12),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_12),
.A2(n_68),
.B1(n_69),
.B2(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_114),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_51),
.B1(n_68),
.B2(n_69),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_13),
.A2(n_51),
.B1(n_63),
.B2(n_65),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_14),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_14),
.A2(n_40),
.B1(n_68),
.B2(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_14),
.A2(n_40),
.B1(n_63),
.B2(n_65),
.Y(n_271)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_333),
.C(n_339),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_331),
.B(n_336),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_319),
.B(n_330),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_281),
.B(n_316),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_258),
.B(n_280),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_140),
.B(n_257),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_115),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_23),
.B(n_115),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_85),
.C(n_95),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_24),
.B(n_85),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_57),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_25),
.B(n_58),
.C(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_26),
.B(n_41),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_34),
.B(n_37),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_27),
.A2(n_33),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_27),
.A2(n_33),
.B1(n_215),
.B2(n_223),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_27),
.A2(n_90),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_28),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_28),
.A2(n_32),
.B1(n_35),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_28),
.A2(n_38),
.B(n_91),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_28),
.A2(n_32),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_30),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_29),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_32),
.B(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_33),
.A2(n_88),
.B(n_101),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_33),
.B(n_104),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_52),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_42),
.A2(n_47),
.B1(n_55),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_42),
.A2(n_55),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_42),
.B(n_104),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_42),
.A2(n_55),
.B1(n_187),
.B2(n_212),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_42),
.A2(n_55),
.B(n_151),
.Y(n_294)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_43),
.B(n_53),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_43),
.A2(n_54),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_43),
.B(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_56)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OA22x2_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_49),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_48),
.B(n_69),
.C(n_79),
.Y(n_183)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_49),
.A2(n_78),
.B(n_182),
.C(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_49),
.B(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_52),
.B(n_197),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_55),
.A2(n_94),
.B(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_55),
.A2(n_137),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_55),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_74),
.B2(n_75),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_67),
.B1(n_70),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_60),
.A2(n_72),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_60),
.B(n_271),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_69),
.B(n_103),
.C(n_105),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_104),
.CON(n_103),
.SN(n_103)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_66),
.C(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_67),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_69),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g182 ( 
.A(n_69),
.B(n_104),
.CON(n_182),
.SN(n_182)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_81),
.B(n_83),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_76),
.A2(n_110),
.B1(n_159),
.B2(n_182),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_76),
.A2(n_110),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_76),
.A2(n_81),
.B(n_110),
.Y(n_326)
);

AND2x4_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_80),
.A2(n_107),
.B1(n_108),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_80),
.A2(n_108),
.B1(n_149),
.B2(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_83),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_93),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_95),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_106),
.C(n_111),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_97),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_113),
.B1(n_129),
.B2(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_111),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_108),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_109),
.B(n_125),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_139),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_131),
.B2(n_132),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_117),
.B(n_132),
.C(n_139),
.Y(n_279)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_119),
.B(n_123),
.C(n_127),
.Y(n_261)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_124),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_128),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_129),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_129),
.A2(n_145),
.B1(n_287),
.B2(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_129),
.A2(n_130),
.B(n_145),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_130),
.A2(n_145),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_133),
.A2(n_134),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_134),
.B(n_136),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_134),
.A2(n_266),
.B(n_269),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_136),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_170),
.B(n_252),
.C(n_256),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_163),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_163),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.C(n_156),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_143),
.B(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.C(n_152),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_145),
.A2(n_270),
.B(n_305),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_157),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_164),
.B(n_168),
.C(n_169),
.Y(n_253)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_246),
.B(n_251),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_201),
.B(n_245),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_189),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_175),
.B(n_189),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.C(n_185),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_176),
.A2(n_177),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_185),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_190),
.B(n_195),
.C(n_199),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_200),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_239),
.B(n_244),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_229),
.B(n_238),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_218),
.B(n_228),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_213),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_213),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_227),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_243),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_279),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_279),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_264),
.C(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_273),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B(n_278),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_284),
.C(n_298),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_278),
.A2(n_284),
.B1(n_285),
.B2(n_315),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_311),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_282),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_299),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_289),
.B1(n_296),
.B2(n_297),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_291),
.C(n_294),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_296),
.B1(n_303),
.B2(n_309),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_295),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_304),
.C(n_308),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_300),
.C(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_310),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_321),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_325),
.C(n_327),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule