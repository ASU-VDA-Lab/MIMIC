module fake_jpeg_32065_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_50),
.Y(n_52)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_27),
.B(n_0),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_37),
.B1(n_28),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_57),
.B1(n_28),
.B2(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_37),
.B1(n_28),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_30),
.B1(n_23),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_98)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_28),
.B1(n_23),
.B2(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_30),
.B1(n_23),
.B2(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_26),
.Y(n_79)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_23),
.B1(n_35),
.B2(n_32),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_20),
.B(n_24),
.C(n_29),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_27),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_50),
.B(n_42),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_97),
.C(n_104),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_39),
.B1(n_42),
.B2(n_46),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_78),
.B1(n_92),
.B2(n_73),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_43),
.B(n_44),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_48),
.C(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_82),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_40),
.B1(n_46),
.B2(n_45),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_31),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_87),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_88),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_89),
.B(n_68),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_103),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_39),
.B1(n_24),
.B2(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_102),
.Y(n_119)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_31),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_29),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_20),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_27),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_73),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_71),
.C(n_44),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_110),
.C(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_43),
.C(n_36),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_104),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_127),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_97),
.Y(n_142)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_69),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_79),
.B(n_77),
.C(n_95),
.D(n_96),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_83),
.C(n_91),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_60),
.B1(n_61),
.B2(n_20),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_43),
.C(n_47),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_97),
.B1(n_101),
.B2(n_68),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_61),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_89),
.B1(n_81),
.B2(n_98),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_121),
.B1(n_135),
.B2(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_131),
.B(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_103),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_102),
.B(n_104),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_106),
.B(n_124),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_99),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_159),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_158),
.B1(n_127),
.B2(n_113),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_24),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_67),
.B1(n_66),
.B2(n_101),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_94),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_33),
.B1(n_21),
.B2(n_25),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_25),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_109),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_129),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_134),
.C(n_108),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_194),
.C(n_196),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_173),
.B1(n_182),
.B2(n_147),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_118),
.B1(n_116),
.B2(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_192),
.B1(n_198),
.B2(n_166),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_178),
.B(n_181),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_152),
.B1(n_157),
.B2(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_106),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_191),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_117),
.B(n_33),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_189),
.B(n_144),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_126),
.B(n_21),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_133),
.B(n_60),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_133),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_136),
.A2(n_101),
.B1(n_67),
.B2(n_90),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_67),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_165),
.C(n_148),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_129),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_23),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_160),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_141),
.A2(n_90),
.B1(n_100),
.B2(n_53),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_158),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_205),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_164),
.B1(n_151),
.B2(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_143),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_215),
.C(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_228),
.B1(n_202),
.B2(n_200),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_139),
.C(n_140),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_139),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_167),
.C(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_160),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_192),
.B1(n_174),
.B2(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_179),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

OAI22x1_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_126),
.B1(n_138),
.B2(n_129),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_138),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_163),
.C(n_156),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_168),
.C(n_175),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_173),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_12),
.Y(n_229)
);

OAI322xp33_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_174),
.A3(n_171),
.B1(n_183),
.B2(n_178),
.C1(n_15),
.C2(n_9),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_247),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_180),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_239),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_200),
.B(n_225),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_172),
.B1(n_182),
.B2(n_194),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_245),
.B1(n_48),
.B2(n_53),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_171),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_188),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_253),
.C(n_255),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_175),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_198),
.B1(n_169),
.B2(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_169),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_251),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_195),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_187),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_206),
.A2(n_187),
.B1(n_90),
.B2(n_100),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_216),
.B1(n_214),
.B2(n_212),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_126),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_48),
.A3(n_53),
.B1(n_9),
.B2(n_16),
.C1(n_14),
.C2(n_13),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_205),
.A3(n_222),
.B1(n_220),
.B2(n_208),
.C1(n_209),
.C2(n_48),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_260),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_223),
.B(n_226),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_273),
.B(n_245),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_262),
.A2(n_255),
.B1(n_244),
.B2(n_241),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_234),
.B1(n_249),
.B2(n_231),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_212),
.C(n_228),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_269),
.C(n_270),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_224),
.C(n_84),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_243),
.C(n_251),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_16),
.B(n_14),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_48),
.B1(n_18),
.B2(n_2),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_287),
.C(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_232),
.C(n_248),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_257),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_84),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_84),
.C(n_48),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_295),
.C(n_272),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_259),
.B1(n_1),
.B2(n_2),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_18),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_18),
.C(n_16),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_258),
.B1(n_274),
.B2(n_261),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_299),
.B(n_306),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_258),
.B1(n_278),
.B2(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_0),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_257),
.C(n_264),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_286),
.C(n_290),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_276),
.B1(n_262),
.B2(n_266),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_291),
.B(n_285),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_284),
.A2(n_275),
.B(n_10),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_295),
.B(n_1),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_0),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_281),
.B1(n_292),
.B2(n_279),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_312),
.A2(n_308),
.B(n_301),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_310),
.B(n_280),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_324),
.B(n_293),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_318),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_323),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_307),
.B(n_297),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_311),
.C(n_306),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_325),
.A2(n_328),
.B(n_333),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_320),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_319),
.C(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_331),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_18),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_312),
.A2(n_1),
.B(n_3),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_332),
.B(n_334),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_3),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_341),
.B(n_8),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_325),
.A2(n_330),
.B(n_329),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g345 ( 
.A1(n_336),
.A2(n_339),
.B(n_4),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_325),
.A2(n_320),
.B1(n_5),
.B2(n_6),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_18),
.B(n_5),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_344),
.B(n_340),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_337),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_346),
.A2(n_342),
.B1(n_347),
.B2(n_7),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_5),
.Y(n_349)
);


endmodule