module fake_aes_2547_n_495 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_495);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_495;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_479;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_70), .B(n_101), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_82), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_49), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_94), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_56), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_105), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_66), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_63), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_9), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_2), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_60), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_55), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_18), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_40), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_89), .Y(n_131) );
INVxp67_ASAP7_75t_SL g132 ( .A(n_97), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_43), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_95), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_109), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_39), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_108), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_69), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_103), .Y(n_140) );
BUFx5_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
INVxp33_ASAP7_75t_L g142 ( .A(n_44), .Y(n_142) );
INVxp33_ASAP7_75t_SL g143 ( .A(n_67), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_62), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_39), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_53), .B(n_28), .Y(n_146) );
INVxp67_ASAP7_75t_SL g147 ( .A(n_17), .Y(n_147) );
INVx2_ASAP7_75t_SL g148 ( .A(n_76), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_30), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_16), .Y(n_151) );
INVxp33_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_41), .Y(n_153) );
INVxp33_ASAP7_75t_SL g154 ( .A(n_23), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_19), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_48), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_79), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_13), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_75), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_61), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_92), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_77), .B(n_45), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_32), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_4), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_64), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_90), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_24), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_31), .Y(n_168) );
INVxp33_ASAP7_75t_L g169 ( .A(n_107), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_71), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_52), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_41), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_68), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_2), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_104), .Y(n_175) );
INVxp33_ASAP7_75t_SL g176 ( .A(n_84), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_42), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_57), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_96), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_78), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_54), .Y(n_181) );
NOR2xp67_ASAP7_75t_L g182 ( .A(n_106), .B(n_100), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_81), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_14), .Y(n_184) );
INVxp33_ASAP7_75t_L g185 ( .A(n_102), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_181), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_116), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_116), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_116), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_116), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_128), .B(n_0), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_116), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_124), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_124), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_142), .B(n_1), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
INVx5_ASAP7_75t_L g204 ( .A(n_140), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_115), .A2(n_1), .B(n_3), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_141), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_141), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_117), .B(n_3), .Y(n_217) );
BUFx8_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_177), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_184), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_209), .B(n_170), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_204), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_212), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_216), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_194), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_212), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_212), .B(n_148), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_194), .B(n_119), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_207), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_212), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_189), .B(n_148), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_209), .A2(n_134), .B1(n_113), .B2(n_120), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_204), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_217), .B(n_152), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_207), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_189), .B(n_145), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_211), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
NOR2x1p5_ASAP7_75t_L g246 ( .A(n_186), .B(n_130), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_217), .B(n_152), .Y(n_248) );
BUFx6f_ASAP7_75t_SL g249 ( .A(n_197), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_189), .B(n_170), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_195), .B(n_169), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
NAND3x1_ASAP7_75t_L g253 ( .A(n_195), .B(n_170), .C(n_134), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_214), .Y(n_254) );
INVx8_ASAP7_75t_L g255 ( .A(n_192), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_255), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_255), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_255), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_242), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_227), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_253), .B(n_202), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_255), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_238), .B(n_118), .Y(n_263) );
INVx4_ASAP7_75t_SL g264 ( .A(n_249), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_238), .A2(n_218), .B1(n_209), .B2(n_192), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_228), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_248), .B(n_218), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_223), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_255), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_253), .B(n_145), .Y(n_272) );
NAND2xp33_ASAP7_75t_L g273 ( .A(n_223), .B(n_141), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_240), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_251), .B(n_192), .Y(n_275) );
INVx5_ASAP7_75t_L g276 ( .A(n_224), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_240), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_231), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_231), .B(n_218), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_240), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_250), .B(n_206), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_246), .A2(n_154), .B1(n_112), .B2(n_123), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_234), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_236), .B(n_206), .Y(n_284) );
AND2x6_ASAP7_75t_SL g285 ( .A(n_230), .B(n_110), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_236), .A2(n_209), .B1(n_210), .B2(n_206), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_225), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_249), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_229), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_229), .B(n_206), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_233), .B(n_210), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_224), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_232), .Y(n_293) );
BUFx12f_ASAP7_75t_L g294 ( .A(n_226), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_232), .Y(n_295) );
INVx3_ASAP7_75t_SL g296 ( .A(n_232), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_235), .A2(n_157), .B1(n_183), .B2(n_122), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_235), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_235), .B(n_210), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_296), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_288), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_267), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_260), .B(n_137), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_283), .B(n_151), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_278), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_284), .A2(n_197), .B(n_198), .C(n_214), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_288), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_296), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_256), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_263), .A2(n_198), .B(n_219), .C(n_215), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_257), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_275), .B(n_143), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_266), .A2(n_215), .B(n_219), .C(n_190), .Y(n_315) );
AOI21xp33_ASAP7_75t_L g316 ( .A1(n_279), .A2(n_185), .B(n_176), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_264), .B(n_147), .Y(n_317) );
CKINVDCx11_ASAP7_75t_R g318 ( .A(n_285), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_257), .Y(n_320) );
OAI22x1_ASAP7_75t_L g321 ( .A1(n_298), .A2(n_209), .B1(n_150), .B2(n_164), .Y(n_321) );
BUFx4f_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_273), .A2(n_243), .B(n_239), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_258), .Y(n_324) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_277), .A2(n_219), .B(n_215), .C(n_201), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_261), .A2(n_176), .B1(n_243), .B2(n_239), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_272), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_281), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
NOR2xp67_ASAP7_75t_R g331 ( .A(n_262), .B(n_125), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_268), .B(n_245), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_258), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_272), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_282), .B(n_208), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_300), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_270), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_289), .B(n_252), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_289), .B(n_252), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_264), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_259), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_297), .B(n_213), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_291), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_291), .B(n_172), .Y(n_348) );
INVx6_ASAP7_75t_L g349 ( .A(n_294), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_287), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_328), .A2(n_286), .B1(n_269), .B2(n_271), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_330), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_323), .A2(n_269), .B(n_265), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_322), .A2(n_174), .B1(n_153), .B2(n_156), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_301), .B(n_265), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_301), .B1(n_326), .B2(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_348), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_303), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_346), .Y(n_359) );
AO31x2_ASAP7_75t_L g360 ( .A1(n_315), .A2(n_188), .A3(n_193), .B(n_187), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_316), .B(n_201), .C(n_200), .Y(n_361) );
NOR2x1_ASAP7_75t_R g362 ( .A(n_318), .B(n_166), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_304), .B(n_200), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_350), .B(n_292), .Y(n_364) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_182), .B(n_187), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_310), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_350), .B(n_292), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_163), .B1(n_168), .B2(n_167), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g369 ( .A1(n_314), .A2(n_222), .B1(n_221), .B2(n_220), .C(n_132), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_305), .B(n_306), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g371 ( .A1(n_311), .A2(n_115), .B(n_139), .C(n_127), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_321), .A2(n_126), .B1(n_129), .B2(n_121), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_349), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_339), .B(n_276), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_327), .A2(n_114), .B1(n_162), .B2(n_146), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_335), .A2(n_133), .B1(n_135), .B2(n_131), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_317), .A2(n_138), .B1(n_144), .B2(n_136), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_341), .A2(n_160), .B1(n_161), .B2(n_159), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_307), .A2(n_188), .A3(n_193), .B(n_187), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_312), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_342), .A2(n_173), .B1(n_175), .B2(n_171), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_332), .A2(n_179), .B1(n_180), .B2(n_178), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_319), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_331), .B(n_237), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_325), .A2(n_244), .B(n_241), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_320), .B1(n_324), .B2(n_313), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_359), .A2(n_344), .B1(n_302), .B2(n_308), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_361), .A2(n_345), .B1(n_338), .B2(n_337), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_361), .A2(n_337), .B1(n_340), .B2(n_334), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_372), .B(n_111), .C(n_196), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_358), .B(n_5), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_363), .A2(n_308), .B1(n_333), .B2(n_329), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_354), .A2(n_196), .B1(n_199), .B2(n_247), .Y(n_396) );
OAI21x1_ASAP7_75t_SL g397 ( .A1(n_356), .A2(n_199), .B(n_6), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_377), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_379), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_373), .B(n_7), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_357), .Y(n_402) );
AO31x2_ASAP7_75t_L g403 ( .A1(n_351), .A2(n_205), .A3(n_203), .B(n_8), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_369), .A2(n_205), .B1(n_226), .B2(n_10), .Y(n_404) );
AO31x2_ASAP7_75t_L g405 ( .A1(n_353), .A2(n_13), .A3(n_11), .B(n_12), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_382), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_353), .A2(n_51), .B(n_50), .Y(n_407) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_362), .A2(n_368), .B1(n_378), .B2(n_380), .C1(n_383), .C2(n_376), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_20), .B(n_21), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_375), .B(n_22), .C(n_23), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_384), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_367), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_374), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_364), .Y(n_415) );
AO31x2_ASAP7_75t_L g416 ( .A1(n_387), .A2(n_33), .A3(n_34), .B(n_35), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_367), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_408), .A2(n_365), .B(n_386), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_389), .B(n_381), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_410), .A2(n_360), .B1(n_46), .B2(n_47), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_394), .B(n_65), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_401), .B(n_74), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_402), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_412), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_409), .A2(n_98), .B(n_99), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_407), .A2(n_397), .B(n_392), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_405), .Y(n_434) );
AOI33xp33_ASAP7_75t_L g435 ( .A1(n_413), .A2(n_417), .A3(n_396), .B1(n_415), .B2(n_404), .B3(n_388), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_398), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_393), .A2(n_391), .B(n_414), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_416), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_434), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_437), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_420), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_419), .A2(n_395), .B(n_390), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_439), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_422), .B(n_403), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_423), .B(n_403), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_427), .B(n_418), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_428), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_436), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_438), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_438), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_426), .B(n_421), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_435), .B(n_425), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_433), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_433), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_433), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_431), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_429), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_430), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_446), .B(n_447), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_443), .B(n_440), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_451), .B(n_450), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_441), .B(n_442), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_448), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_445), .B(n_461), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_449), .B(n_455), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_452), .B(n_453), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_458), .B(n_457), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_454), .B(n_460), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_458), .B(n_456), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_466), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_468), .B(n_444), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_462), .B(n_459), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_471), .B(n_459), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_472), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_464), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_467), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_473), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_475), .B(n_469), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_479), .B(n_463), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_478), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_474), .B(n_465), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_476), .B(n_470), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_477), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_483), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_487), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_488), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_489), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_490), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_491), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_492), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_493), .A2(n_480), .B(n_484), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_494), .A2(n_486), .B1(n_482), .B2(n_485), .C(n_481), .Y(n_495) );
endmodule