module real_jpeg_29262_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI221xp5_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_8),
.B1(n_13),
.B2(n_20),
.C(n_22),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g9 ( 
.A(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_4),
.B(n_17),
.Y(n_33)
);

OR2x2_ASAP7_75t_SL g11 ( 
.A(n_5),
.B(n_12),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_28),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

OR2x2_ASAP7_75t_SL g42 ( 
.A(n_12),
.B(n_37),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_23),
.B(n_25),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_16),
.B(n_17),
.Y(n_13)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_35),
.B1(n_38),
.B2(n_42),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);


endmodule