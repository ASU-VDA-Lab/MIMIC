module fake_netlist_6_2206_n_170 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_170);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_170;

wire n_52;
wire n_119;
wire n_91;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_85;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_66;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_22),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_1),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_2),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_7),
.B1(n_9),
.B2(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_20),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_33),
.B(n_39),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_61),
.C(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_46),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_41),
.B1(n_34),
.B2(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_40),
.A3(n_38),
.B1(n_45),
.B2(n_34),
.C(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_42),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_35),
.B(n_25),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_23),
.B(n_26),
.C(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_29),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_30),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_55),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_70),
.B(n_60),
.C(n_57),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_55),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_67),
.B(n_70),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_63),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AOI21x1_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_64),
.B(n_56),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_96),
.Y(n_106)
);

BUFx8_ASAP7_75t_SL g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_100),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_82),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_77),
.C(n_80),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_100),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_111),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_115),
.B(n_109),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_73),
.B1(n_107),
.B2(n_85),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

OR2x6_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_93),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_102),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_87),
.C(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_101),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_101),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_124),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND4xp25_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_121),
.C(n_134),
.D(n_124),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_123),
.C(n_86),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_123),
.C(n_129),
.Y(n_142)
);

NOR2x1p5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_59),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_126),
.B1(n_72),
.B2(n_59),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_57),
.C(n_72),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_147),
.B1(n_146),
.B2(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_89),
.C(n_64),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_126),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_152),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_62),
.C(n_66),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_126),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_66),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_150),
.C(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_154),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_160),
.B1(n_159),
.B2(n_157),
.Y(n_167)
);

BUFx2_ASAP7_75t_SL g168 ( 
.A(n_165),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_166),
.B(n_162),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_168),
.B1(n_162),
.B2(n_163),
.Y(n_170)
);


endmodule