module real_aes_2762_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_0), .B(n_138), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_1), .A2(n_147), .B(n_152), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_2), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_3), .B(n_154), .Y(n_192) );
INVx1_ASAP7_75t_L g145 ( .A(n_4), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_5), .B(n_154), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_6), .B(n_164), .Y(n_564) );
INVx1_ASAP7_75t_L g544 ( .A(n_7), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_8), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_9), .Y(n_510) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_10), .B(n_156), .Y(n_181) );
INVx2_ASAP7_75t_L g135 ( .A(n_11), .Y(n_135) );
AOI221x1_ASAP7_75t_L g227 ( .A1(n_12), .A2(n_24), .B1(n_138), .B2(n_147), .C(n_228), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_14), .B(n_138), .Y(n_177) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_15), .A2(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g572 ( .A(n_16), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_17), .B(n_158), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_18), .B(n_154), .Y(n_168) );
AO21x1_ASAP7_75t_L g187 ( .A1(n_19), .A2(n_138), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
INVx1_ASAP7_75t_L g570 ( .A(n_21), .Y(n_570) );
INVx1_ASAP7_75t_SL g492 ( .A(n_22), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_23), .B(n_139), .Y(n_560) );
NAND2x1_ASAP7_75t_L g200 ( .A(n_25), .B(n_154), .Y(n_200) );
AOI33xp33_ASAP7_75t_L g530 ( .A1(n_26), .A2(n_53), .A3(n_475), .B1(n_480), .B2(n_531), .B3(n_532), .Y(n_530) );
NAND2x1_ASAP7_75t_L g219 ( .A(n_27), .B(n_156), .Y(n_219) );
INVx1_ASAP7_75t_L g503 ( .A(n_28), .Y(n_503) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_29), .A2(n_88), .B(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g160 ( .A(n_29), .B(n_88), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_30), .B(n_483), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_31), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_32), .B(n_154), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_33), .B(n_156), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_34), .A2(n_147), .B(n_208), .Y(n_207) );
AOI22xp5_ASAP7_75t_SL g791 ( .A1(n_35), .A2(n_792), .B1(n_798), .B2(n_799), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_35), .Y(n_798) );
AND2x2_ASAP7_75t_L g144 ( .A(n_36), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g148 ( .A(n_36), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g474 ( .A(n_36), .Y(n_474) );
OR2x6_ASAP7_75t_L g111 ( .A(n_37), .B(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_38), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_39), .B(n_138), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_40), .B(n_483), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_41), .A2(n_133), .B1(n_164), .B2(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_42), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_43), .B(n_139), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_44), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_45), .B(n_156), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_46), .B(n_175), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_47), .B(n_139), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_48), .A2(n_147), .B(n_218), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_49), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_50), .A2(n_85), .B1(n_120), .B2(n_121), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_50), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_51), .A2(n_80), .B1(n_795), .B2(n_796), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_51), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_52), .B(n_156), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_54), .B(n_139), .Y(n_521) );
INVx1_ASAP7_75t_L g141 ( .A(n_55), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_55), .Y(n_151) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_56), .A2(n_104), .B1(n_447), .B2(n_452), .C1(n_808), .C2(n_813), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_56), .A2(n_116), .B1(n_442), .B2(n_443), .Y(n_115) );
INVxp67_ASAP7_75t_L g443 ( .A(n_56), .Y(n_443) );
AND2x2_ASAP7_75t_L g522 ( .A(n_56), .B(n_158), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_57), .A2(n_74), .B1(n_472), .B2(n_483), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_58), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_59), .B(n_154), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_60), .B(n_133), .Y(n_512) );
AOI21xp5_ASAP7_75t_SL g471 ( .A1(n_61), .A2(n_472), .B(n_477), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_62), .A2(n_147), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g567 ( .A(n_63), .Y(n_567) );
AO21x1_ASAP7_75t_L g189 ( .A1(n_64), .A2(n_147), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_65), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_66), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g520 ( .A(n_67), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_68), .B(n_138), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_69), .A2(n_472), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g212 ( .A(n_70), .B(n_159), .Y(n_212) );
INVx1_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_71), .Y(n_149) );
AND2x2_ASAP7_75t_L g223 ( .A(n_72), .B(n_132), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_73), .B(n_483), .Y(n_533) );
AND2x2_ASAP7_75t_L g494 ( .A(n_75), .B(n_132), .Y(n_494) );
INVx1_ASAP7_75t_L g568 ( .A(n_76), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_77), .A2(n_472), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_78), .A2(n_118), .B1(n_119), .B2(n_122), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_78), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_79), .A2(n_472), .B(n_525), .C(n_559), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_80), .Y(n_795) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
AND2x2_ASAP7_75t_L g131 ( .A(n_82), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_83), .B(n_138), .Y(n_170) );
AND2x2_ASAP7_75t_SL g469 ( .A(n_84), .B(n_132), .Y(n_469) );
INVx1_ASAP7_75t_L g120 ( .A(n_85), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_86), .A2(n_472), .B1(n_528), .B2(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g188 ( .A(n_87), .B(n_164), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_89), .B(n_156), .Y(n_169) );
AND2x2_ASAP7_75t_L g204 ( .A(n_90), .B(n_132), .Y(n_204) );
INVx1_ASAP7_75t_L g478 ( .A(n_91), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_92), .B(n_154), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_93), .A2(n_793), .B1(n_794), .B2(n_797), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_93), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_94), .A2(n_147), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_95), .B(n_156), .Y(n_229) );
AND2x2_ASAP7_75t_L g534 ( .A(n_96), .B(n_132), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_97), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_98), .A2(n_501), .B(n_502), .C(n_505), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_99), .Y(n_806) );
BUFx2_ASAP7_75t_L g451 ( .A(n_100), .Y(n_451) );
BUFx2_ASAP7_75t_SL g817 ( .A(n_100), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_101), .A2(n_147), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_102), .B(n_139), .Y(n_481) );
OAI21x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_115), .B(n_444), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g446 ( .A(n_108), .Y(n_446) );
BUFx2_ASAP7_75t_L g819 ( .A(n_108), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x6_ASAP7_75t_SL g456 ( .A(n_109), .B(n_111), .Y(n_456) );
OR2x6_ASAP7_75t_SL g458 ( .A(n_109), .B(n_110), .Y(n_458) );
OR2x2_ASAP7_75t_L g807 ( .A(n_109), .B(n_111), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g442 ( .A(n_116), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_123), .B1(n_440), .B2(n_441), .Y(n_116) );
INVx1_ASAP7_75t_L g440 ( .A(n_117), .Y(n_440) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g441 ( .A(n_123), .Y(n_441) );
INVx3_ASAP7_75t_L g803 ( .A(n_123), .Y(n_803) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_349), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_267), .C(n_293), .D(n_333), .Y(n_124) );
OAI211xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_182), .B(n_213), .C(n_253), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_161), .Y(n_127) );
AND2x2_ASAP7_75t_L g420 ( .A(n_128), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_129), .B(n_161), .Y(n_287) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g214 ( .A(n_130), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_130), .B(n_240), .Y(n_239) );
INVx5_ASAP7_75t_L g273 ( .A(n_130), .Y(n_273) );
NOR2x1_ASAP7_75t_SL g315 ( .A(n_130), .B(n_162), .Y(n_315) );
AND2x2_ASAP7_75t_L g371 ( .A(n_130), .B(n_174), .Y(n_371) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
INVx3_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_132), .A2(n_203), .B1(n_500), .B2(n_506), .Y(n_499) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_133), .B(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_135), .B(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g164 ( .A(n_135), .B(n_160), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_158), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g504 ( .A(n_139), .Y(n_504) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x6_ASAP7_75t_L g156 ( .A(n_140), .B(n_149), .Y(n_156) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g154 ( .A(n_142), .B(n_151), .Y(n_154) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_144), .Y(n_505) );
AND2x2_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_145), .Y(n_485) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g486 ( .A(n_148), .Y(n_486) );
INVx2_ASAP7_75t_L g476 ( .A(n_149), .Y(n_476) );
AND2x4_ASAP7_75t_L g472 ( .A(n_150), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g480 ( .A(n_151), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
INVxp67_ASAP7_75t_L g573 ( .A(n_154), .Y(n_573) );
INVxp67_ASAP7_75t_L g571 ( .A(n_156), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_157), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_157), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_157), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_157), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_157), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_157), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_157), .A2(n_229), .B(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_157), .A2(n_478), .B(n_479), .C(n_481), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_157), .A2(n_479), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_157), .A2(n_479), .B(n_520), .C(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g528 ( .A(n_157), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_157), .A2(n_479), .B(n_544), .C(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_157), .A2(n_560), .B(n_561), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_157), .B(n_164), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_158), .Y(n_222) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_158), .A2(n_227), .B(n_231), .Y(n_226) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_158), .A2(n_227), .B(n_231), .Y(n_266) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_173), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_162), .B(n_174), .Y(n_243) );
AND2x2_ASAP7_75t_L g304 ( .A(n_162), .B(n_273), .Y(n_304) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_171), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_163), .B(n_172), .Y(n_171) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_163), .A2(n_165), .B(n_171), .Y(n_257) );
INVx1_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_164), .A2(n_177), .B(n_178), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_164), .B(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_164), .A2(n_471), .B(n_482), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
AND2x2_ASAP7_75t_L g316 ( .A(n_173), .B(n_240), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_173), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g360 ( .A(n_173), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g393 ( .A(n_173), .B(n_214), .Y(n_393) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g237 ( .A(n_174), .Y(n_237) );
AND2x2_ASAP7_75t_L g270 ( .A(n_174), .B(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
OR2x2_ASAP7_75t_L g381 ( .A(n_174), .B(n_240), .Y(n_381) );
INVx2_ASAP7_75t_SL g525 ( .A(n_175), .Y(n_525) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_175), .A2(n_542), .B(n_546), .Y(n_541) );
INVx1_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_195), .Y(n_183) );
AOI211x1_ASAP7_75t_SL g310 ( .A1(n_184), .A2(n_302), .B(n_311), .C(n_313), .Y(n_310) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_184), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_184), .B(n_353), .Y(n_400) );
BUFx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g250 ( .A(n_185), .Y(n_250) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g225 ( .A(n_186), .Y(n_225) );
OAI21x1_ASAP7_75t_SL g186 ( .A1(n_187), .A2(n_189), .B(n_193), .Y(n_186) );
INVx1_ASAP7_75t_L g194 ( .A(n_188), .Y(n_194) );
AOI322xp5_ASAP7_75t_L g213 ( .A1(n_195), .A2(n_214), .A3(n_224), .B1(n_232), .B2(n_235), .C1(n_241), .C2(n_244), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_195), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
INVx2_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
INVxp67_ASAP7_75t_L g290 ( .A(n_196), .Y(n_290) );
BUFx3_ASAP7_75t_L g354 ( .A(n_196), .Y(n_354) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_203), .B(n_204), .Y(n_196) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_197), .A2(n_203), .B(n_204), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_203), .A2(n_206), .B(n_212), .Y(n_205) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_203), .A2(n_206), .B(n_212), .Y(n_252) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_203), .A2(n_516), .B(n_522), .Y(n_515) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_203), .A2(n_516), .B(n_522), .Y(n_538) );
INVx2_ASAP7_75t_L g263 ( .A(n_205), .Y(n_263) );
AND2x2_ASAP7_75t_L g312 ( .A(n_205), .B(n_226), .Y(n_312) );
AND2x2_ASAP7_75t_L g356 ( .A(n_205), .B(n_265), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_211), .Y(n_206) );
AND2x2_ASAP7_75t_L g241 ( .A(n_214), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_214), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_214), .B(n_270), .Y(n_435) );
INVx4_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
AND2x2_ASAP7_75t_L g272 ( .A(n_215), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_215), .Y(n_325) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_223), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_222), .A2(n_488), .B(n_494), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_224), .B(n_309), .Y(n_334) );
INVx1_ASAP7_75t_SL g373 ( .A(n_224), .Y(n_373) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
AND2x4_ASAP7_75t_L g264 ( .A(n_225), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_225), .B(n_263), .Y(n_332) );
AND2x2_ASAP7_75t_L g384 ( .A(n_225), .B(n_234), .Y(n_384) );
OR2x2_ASAP7_75t_L g408 ( .A(n_225), .B(n_226), .Y(n_408) );
AND2x2_ASAP7_75t_L g232 ( .A(n_226), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g282 ( .A(n_226), .B(n_263), .Y(n_282) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_226), .B(n_250), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_232), .B(n_345), .Y(n_362) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx2_ASAP7_75t_L g297 ( .A(n_234), .Y(n_297) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_234), .B(n_251), .Y(n_337) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
OR2x2_ASAP7_75t_L g285 ( .A(n_236), .B(n_239), .Y(n_285) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g254 ( .A(n_237), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g402 ( .A(n_237), .B(n_315), .Y(n_402) );
AND2x2_ASAP7_75t_L g418 ( .A(n_237), .B(n_272), .Y(n_418) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI311xp33_ASAP7_75t_L g388 ( .A1(n_239), .A2(n_327), .A3(n_389), .B(n_391), .C(n_398), .Y(n_388) );
AND2x4_ASAP7_75t_L g255 ( .A(n_240), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_240), .B(n_273), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_240), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g372 ( .A(n_240), .B(n_359), .Y(n_372) );
AND2x2_ASAP7_75t_L g258 ( .A(n_242), .B(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_243), .Y(n_276) );
OR2x2_ASAP7_75t_L g365 ( .A(n_243), .B(n_329), .Y(n_365) );
INVx1_ASAP7_75t_L g421 ( .A(n_243), .Y(n_421) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g330 ( .A(n_247), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g344 ( .A(n_247), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g419 ( .A(n_247), .B(n_292), .Y(n_419) );
BUFx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g262 ( .A(n_248), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g281 ( .A(n_248), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g343 ( .A(n_249), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_249), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_398) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g292 ( .A(n_250), .B(n_263), .Y(n_292) );
AND2x4_ASAP7_75t_L g345 ( .A(n_250), .B(n_252), .Y(n_345) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI21xp33_ASAP7_75t_SL g253 ( .A1(n_254), .A2(n_258), .B(n_260), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_254), .A2(n_340), .B1(n_344), .B2(n_346), .Y(n_339) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_255), .B(n_273), .Y(n_299) );
INVx2_ASAP7_75t_L g361 ( .A(n_255), .Y(n_361) );
AND2x2_ASAP7_75t_L g375 ( .A(n_255), .B(n_371), .Y(n_375) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g271 ( .A(n_257), .Y(n_271) );
INVx1_ASAP7_75t_L g324 ( .A(n_257), .Y(n_324) );
INVx1_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
AND3x2_ASAP7_75t_L g303 ( .A(n_259), .B(n_304), .C(n_305), .Y(n_303) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g367 ( .A(n_262), .Y(n_367) );
AND2x2_ASAP7_75t_L g295 ( .A(n_264), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g366 ( .A(n_264), .B(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_264), .A2(n_378), .B1(n_382), .B2(n_385), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_264), .B(n_412), .Y(n_416) );
BUFx2_ASAP7_75t_L g307 ( .A(n_265), .Y(n_307) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g278 ( .A(n_266), .Y(n_278) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_266), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_277), .B1(n_279), .B2(n_280), .C(n_283), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_274), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g359 ( .A(n_271), .Y(n_359) );
INVx2_ASAP7_75t_SL g348 ( .A(n_272), .Y(n_348) );
AND2x2_ASAP7_75t_L g430 ( .A(n_272), .B(n_297), .Y(n_430) );
INVx4_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
INVx1_ASAP7_75t_L g279 ( .A(n_274), .Y(n_279) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x4_ASAP7_75t_L g390 ( .A(n_278), .B(n_345), .Y(n_390) );
INVx1_ASAP7_75t_SL g429 ( .A(n_278), .Y(n_429) );
AND2x2_ASAP7_75t_L g434 ( .A(n_278), .B(n_337), .Y(n_434) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g376 ( .A(n_282), .Y(n_376) );
OAI21xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_286), .B(n_288), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g306 ( .A(n_292), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g396 ( .A(n_292), .B(n_397), .Y(n_396) );
OAI211xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_298), .B(n_300), .C(n_317), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g389 ( .A(n_296), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_297), .B(n_312), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_297), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g422 ( .A(n_297), .B(n_345), .Y(n_422) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_298), .A2(n_322), .B1(n_334), .B2(n_335), .C(n_339), .Y(n_333) );
INVx3_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g404 ( .A(n_299), .B(n_305), .Y(n_404) );
OAI32xp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_306), .A3(n_308), .B1(n_310), .B2(n_314), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_304), .Y(n_394) );
INVx2_ASAP7_75t_L g327 ( .A(n_305), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g436 ( .A1(n_305), .A2(n_357), .B(n_437), .C(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
OR2x2_ASAP7_75t_L g438 ( .A(n_307), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_311), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g399 ( .A(n_314), .Y(n_399) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
OAI21xp33_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_326), .B(n_330), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
OR2x2_ASAP7_75t_L g357 ( .A(n_320), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_321), .B(n_324), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_323), .A2(n_355), .B1(n_424), .B2(n_427), .C(n_431), .Y(n_423) );
INVx2_ASAP7_75t_L g426 ( .A(n_323), .Y(n_426) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
OR2x2_ASAP7_75t_L g347 ( .A(n_327), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g414 ( .A(n_327), .B(n_372), .Y(n_414) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g412 ( .A(n_337), .Y(n_412) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_345), .B(n_375), .Y(n_432) );
INVx2_ASAP7_75t_L g439 ( .A(n_345), .Y(n_439) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_347), .A2(n_410), .B1(n_413), .B2(n_415), .C(n_417), .Y(n_409) );
AND5x1_ASAP7_75t_L g349 ( .A(n_350), .B(n_388), .C(n_403), .D(n_423), .E(n_433), .Y(n_349) );
NOR2xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_368), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_357), .B1(n_360), .B2(n_362), .C(n_363), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI221xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_373), .B1(n_374), .B2(n_376), .C(n_377), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_373), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
OR2x2_ASAP7_75t_L g386 ( .A(n_381), .B(n_387), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_395), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_422), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_419), .A2(n_434), .B(n_435), .C(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22x1_ASAP7_75t_L g453 ( .A1(n_441), .A2(n_454), .B1(n_457), .B2(n_459), .Y(n_453) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g809 ( .A(n_446), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_SL g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx2_ASAP7_75t_L g812 ( .A(n_449), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_449), .A2(n_815), .B(n_818), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_451), .B(n_812), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_791), .B(n_800), .Y(n_452) );
INVx3_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_456), .Y(n_455) );
CKINVDCx11_ASAP7_75t_R g804 ( .A(n_456), .Y(n_804) );
INVx1_ASAP7_75t_SL g802 ( .A(n_457), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
OAI22x1_ASAP7_75t_L g801 ( .A1(n_459), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_801) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
AND3x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_681), .C(n_744), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_645), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_586), .C(n_615), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_465), .B(n_575), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_495), .B1(n_535), .B2(n_547), .Y(n_465) );
NAND2x1_ASAP7_75t_L g730 ( .A(n_466), .B(n_576), .Y(n_730) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_487), .Y(n_467) );
INVx2_ASAP7_75t_L g549 ( .A(n_468), .Y(n_549) );
INVx4_ASAP7_75t_L g591 ( .A(n_468), .Y(n_591) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_468), .Y(n_611) );
AND2x4_ASAP7_75t_L g622 ( .A(n_468), .B(n_590), .Y(n_622) );
AND2x2_ASAP7_75t_L g628 ( .A(n_468), .B(n_552), .Y(n_628) );
NOR2x1_ASAP7_75t_SL g758 ( .A(n_468), .B(n_563), .Y(n_758) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g511 ( .A(n_472), .Y(n_511) );
NOR2x1p5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g532 ( .A(n_475), .Y(n_532) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x6_ASAP7_75t_L g479 ( .A(n_476), .B(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g501 ( .A(n_479), .Y(n_501) );
INVx2_ASAP7_75t_L g562 ( .A(n_479), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_479), .A2(n_504), .B1(n_567), .B2(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g484 ( .A(n_480), .B(n_485), .Y(n_484) );
INVxp33_ASAP7_75t_L g531 ( .A(n_480), .Y(n_531) );
INVx1_ASAP7_75t_L g513 ( .A(n_483), .Y(n_513) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g555 ( .A(n_484), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
INVx2_ASAP7_75t_L g594 ( .A(n_487), .Y(n_594) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_487), .Y(n_608) );
INVx1_ASAP7_75t_L g619 ( .A(n_487), .Y(n_619) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_487), .Y(n_631) );
AND2x2_ASAP7_75t_L g663 ( .A(n_487), .B(n_563), .Y(n_663) );
AND2x2_ASAP7_75t_L g695 ( .A(n_487), .B(n_579), .Y(n_695) );
INVx1_ASAP7_75t_L g702 ( .A(n_487), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_514), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g644 ( .A(n_497), .B(n_583), .Y(n_644) );
INVx2_ASAP7_75t_L g718 ( .A(n_497), .Y(n_718) );
AND2x2_ASAP7_75t_L g741 ( .A(n_497), .B(n_514), .Y(n_741) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_498), .B(n_538), .Y(n_582) );
INVx2_ASAP7_75t_L g603 ( .A(n_498), .Y(n_603) );
AND2x4_ASAP7_75t_L g625 ( .A(n_498), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g660 ( .A(n_498), .Y(n_660) );
AND2x2_ASAP7_75t_L g737 ( .A(n_498), .B(n_541), .Y(n_737) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_507), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g708 ( .A(n_514), .Y(n_708) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_515), .B(n_603), .Y(n_633) );
AND2x2_ASAP7_75t_L g638 ( .A(n_515), .B(n_603), .Y(n_638) );
INVx2_ASAP7_75t_L g651 ( .A(n_515), .Y(n_651) );
NOR2x1_ASAP7_75t_L g699 ( .A(n_515), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x4_ASAP7_75t_L g624 ( .A(n_523), .B(n_537), .Y(n_624) );
AND2x2_ASAP7_75t_L g639 ( .A(n_523), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g692 ( .A(n_523), .Y(n_692) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_524), .B(n_541), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_524), .B(n_538), .Y(n_696) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_534), .Y(n_524) );
AO21x2_ASAP7_75t_L g585 ( .A1(n_525), .A2(n_526), .B(n_534), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_527), .B(n_533), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVxp33_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx3_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
AND2x2_ASAP7_75t_L g767 ( .A(n_538), .B(n_768), .Y(n_767) );
INVx3_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_539), .B(n_692), .Y(n_787) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g602 ( .A(n_540), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g583 ( .A(n_541), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g626 ( .A(n_541), .Y(n_626) );
INVxp67_ASAP7_75t_L g640 ( .A(n_541), .Y(n_640) );
INVx1_ASAP7_75t_L g700 ( .A(n_541), .Y(n_700) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_541), .Y(n_768) );
INVx1_ASAP7_75t_L g752 ( .A(n_547), .Y(n_752) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_548), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g706 ( .A(n_549), .B(n_578), .Y(n_706) );
OR2x2_ASAP7_75t_L g742 ( .A(n_550), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g724 ( .A(n_551), .B(n_702), .Y(n_724) );
AND2x2_ASAP7_75t_L g776 ( .A(n_551), .B(n_611), .Y(n_776) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_563), .Y(n_551) );
AND2x4_ASAP7_75t_L g578 ( .A(n_552), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g590 ( .A(n_552), .Y(n_590) );
INVx2_ASAP7_75t_L g607 ( .A(n_552), .Y(n_607) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_552), .Y(n_785) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .Y(n_554) );
INVx3_ASAP7_75t_L g579 ( .A(n_563), .Y(n_579) );
INVx2_ASAP7_75t_L g673 ( .A(n_563), .Y(n_673) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B(n_574), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_572), .B2(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_577), .B(n_653), .Y(n_670) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_577), .B(n_591), .Y(n_712) );
INVx4_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_578), .B(n_653), .Y(n_790) );
AND2x2_ASAP7_75t_L g606 ( .A(n_579), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g620 ( .A(n_579), .Y(n_620) );
AOI22xp5_ASAP7_75t_SL g668 ( .A1(n_580), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_581), .B(n_639), .Y(n_665) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g726 ( .A(n_582), .B(n_614), .Y(n_726) );
AND2x2_ASAP7_75t_L g596 ( .A(n_583), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g632 ( .A(n_583), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g728 ( .A(n_583), .B(n_718), .Y(n_728) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g650 ( .A(n_585), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g676 ( .A(n_585), .Y(n_676) );
AND2x2_ASAP7_75t_L g766 ( .A(n_585), .B(n_603), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_595), .B1(n_599), .B2(n_604), .C(n_609), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
INVx1_ASAP7_75t_L g667 ( .A(n_589), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_589), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_589), .B(n_663), .Y(n_782) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NOR2xp67_ASAP7_75t_SL g635 ( .A(n_591), .B(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_591), .Y(n_648) );
OR2x2_ASAP7_75t_L g732 ( .A(n_591), .B(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_SL g784 ( .A(n_591), .B(n_785), .Y(n_784) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g653 ( .A(n_593), .Y(n_653) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_594), .Y(n_743) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221x1_ASAP7_75t_L g683 ( .A1(n_596), .A2(n_684), .B1(n_686), .B2(n_689), .C(n_693), .Y(n_683) );
AND2x2_ASAP7_75t_L g669 ( .A(n_597), .B(n_625), .Y(n_669) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g612 ( .A(n_600), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_600), .B(n_602), .Y(n_739) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
AND2x2_ASAP7_75t_SL g610 ( .A(n_606), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_606), .B(n_619), .Y(n_636) );
INVx2_ASAP7_75t_L g643 ( .A(n_606), .Y(n_643) );
INVx1_ASAP7_75t_L g688 ( .A(n_607), .Y(n_688) );
BUFx2_ASAP7_75t_L g777 ( .A(n_608), .Y(n_777) );
NAND2xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
OR2x6_ASAP7_75t_L g642 ( .A(n_611), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g723 ( .A(n_611), .B(n_663), .Y(n_723) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_634), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_623), .B1(n_627), .B2(n_632), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_618), .B(n_622), .Y(n_680) );
AND2x4_ASAP7_75t_L g686 ( .A(n_618), .B(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_619), .B(n_620), .Y(n_618) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_619), .Y(n_711) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_622), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_622), .B(n_653), .Y(n_685) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_622), .Y(n_769) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g716 ( .A(n_624), .B(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g677 ( .A(n_625), .Y(n_677) );
NAND2x1_ASAP7_75t_SL g721 ( .A(n_625), .B(n_676), .Y(n_721) );
AND2x2_ASAP7_75t_L g755 ( .A(n_625), .B(n_650), .Y(n_755) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_641), .B2(n_644), .Y(n_634) );
BUFx2_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_637), .A2(n_706), .B1(n_780), .B2(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_638), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g658 ( .A(n_639), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g774 ( .A(n_643), .B(n_775), .C(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g678 ( .A(n_644), .Y(n_678) );
AOI211x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_654), .B(n_656), .C(n_674), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_649), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
AND2x2_ASAP7_75t_L g736 ( .A(n_650), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_650), .B(n_717), .Y(n_748) );
AND2x2_ASAP7_75t_L g780 ( .A(n_650), .B(n_718), .Y(n_780) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g761 ( .A(n_653), .Y(n_761) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g690 ( .A(n_655), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_668), .Y(n_656) );
AOI22xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_661), .B1(n_664), .B2(n_666), .Y(n_657) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g698 ( .A(n_660), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g713 ( .A(n_660), .Y(n_713) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_SL g783 ( .A(n_663), .B(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g719 ( .A(n_672), .B(n_702), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B(n_679), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_676), .B(n_698), .Y(n_773) );
OR2x2_ASAP7_75t_L g751 ( .A(n_677), .B(n_696), .Y(n_751) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_703), .C(n_727), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_686), .A2(n_716), .B1(n_719), .B2(n_720), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_687), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g760 ( .A(n_687), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_687), .B(n_761), .Y(n_764) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI222xp33_ASAP7_75t_L g747 ( .A1(n_691), .A2(n_748), .B1(n_749), .B2(n_750), .C1(n_751), .C2(n_752), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_697), .B2(n_701), .Y(n_693) );
INVx1_ASAP7_75t_SL g733 ( .A(n_695), .Y(n_733) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g770 ( .A(n_699), .B(n_766), .Y(n_770) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_714), .Y(n_703) );
AOI21xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_713), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_722), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_721), .B(n_735), .Y(n_734) );
OAI21xp5_ASAP7_75t_SL g722 ( .A1(n_723), .A2(n_724), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g749 ( .A(n_724), .Y(n_749) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_734), .C(n_738), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B(n_742), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
NAND3x1_ASAP7_75t_L g745 ( .A(n_746), .B(n_771), .C(n_778), .Y(n_745) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_753), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_762), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_755), .B(n_756), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_757), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_765), .B1(n_769), .B2(n_770), .Y(n_762) );
AND2x4_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_772), .B(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_788), .Y(n_778) );
AOI22xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_781), .B1(n_783), .B2(n_786), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI21xp33_ASAP7_75t_L g800 ( .A1(n_791), .A2(n_801), .B(n_805), .Y(n_800) );
INVx1_ASAP7_75t_L g799 ( .A(n_792), .Y(n_799) );
INVx1_ASAP7_75t_L g797 ( .A(n_794), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
BUFx4f_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVxp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx8_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
endmodule