module real_jpeg_24155_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx6_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_19),
.B1(n_21),
.B2(n_57),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_24),
.C(n_29),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_39),
.B1(n_99),
.B2(n_104),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_19),
.B1(n_21),
.B2(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_20),
.B1(n_53),
.B2(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_19),
.B1(n_21),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_77),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_75),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_50),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_15),
.B(n_50),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.C(n_38),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_16),
.A2(n_17),
.B1(n_33),
.B2(n_34),
.Y(n_85)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_18),
.A2(n_22),
.B1(n_30),
.B2(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_19),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_21),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g52 ( 
.A1(n_19),
.A2(n_36),
.A3(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_19),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_37),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_22),
.A2(n_30),
.B1(n_31),
.B2(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_27),
.B(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_28),
.B(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_56),
.B1(n_72),
.B2(n_74),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_60),
.B(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_39),
.A2(n_90),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_40),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_68),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_57),
.CON(n_56),
.SN(n_56)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_86),
.B(n_111),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_95),
.B(n_110),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_94),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_94),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_102),
.B(n_109),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);


endmodule