module fake_netlist_6_3064_n_705 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_705);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_705;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

BUFx10_ASAP7_75t_L g130 ( 
.A(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_42),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_57),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_38),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_116),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_5),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_16),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_41),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_21),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_14),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_12),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_35),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_79),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_46),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_56),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_45),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_29),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_90),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_0),
.B(n_1),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_18),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_19),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_1),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_129),
.A2(n_2),
.B(n_3),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_3),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_20),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_4),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_22),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_137),
.B(n_24),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_138),
.B(n_6),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_141),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_159),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_155),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_143),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVxp33_ASAP7_75t_SL g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

AND3x2_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_146),
.C(n_176),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_142),
.B1(n_178),
.B2(n_156),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

NOR2x1p5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_154),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_160),
.B1(n_166),
.B2(n_146),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_200),
.B(n_171),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_179),
.B1(n_163),
.B2(n_164),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_186),
.B(n_169),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

AND3x2_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_177),
.C(n_175),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_208),
.B(n_162),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_165),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_209),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_212),
.A2(n_173),
.B1(n_172),
.B2(n_170),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_186),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_192),
.Y(n_271)
);

OAI221xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_220),
.B1(n_211),
.B2(n_197),
.C(n_194),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_227),
.Y(n_273)
);

O2A1O1Ixp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_183),
.B(n_206),
.C(n_191),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_230),
.A2(n_205),
.B1(n_212),
.B2(n_181),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

AOI221xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_211),
.B1(n_197),
.B2(n_221),
.C(n_210),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_186),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g280 ( 
.A1(n_230),
.A2(n_209),
.B1(n_189),
.B2(n_181),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_227),
.B(n_226),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_189),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_233),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_219),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_245),
.B1(n_181),
.B2(n_183),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_219),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_226),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_191),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_191),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_224),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_209),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_223),
.B(n_202),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_204),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_254),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_204),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_204),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_225),
.B(n_209),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_206),
.Y(n_302)
);

OR2x6_ASAP7_75t_L g303 ( 
.A(n_225),
.B(n_198),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_223),
.B(n_206),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_258),
.A2(n_219),
.B1(n_221),
.B2(n_217),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_222),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_219),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_248),
.B(n_199),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_229),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_250),
.B(n_199),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_232),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_235),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_250),
.B(n_213),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_213),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_274),
.A2(n_236),
.B(n_198),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_288),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_295),
.B(n_296),
.Y(n_333)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_282),
.B(n_213),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_259),
.B(n_267),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_312),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_281),
.Y(n_337)
);

OAI321xp33_ASAP7_75t_L g338 ( 
.A1(n_285),
.A2(n_213),
.A3(n_214),
.B1(n_215),
.B2(n_217),
.C(n_264),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_296),
.A2(n_302),
.B(n_298),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_298),
.A2(n_259),
.B(n_243),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_214),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_214),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_287),
.A2(n_262),
.B(n_261),
.C(n_252),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_306),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_243),
.B(n_242),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_256),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_217),
.B1(n_215),
.B2(n_214),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_256),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_215),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_280),
.A2(n_256),
.B(n_243),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_271),
.B(n_242),
.Y(n_355)
);

BUFx4f_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_291),
.A2(n_242),
.B(n_217),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_215),
.Y(n_358)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_217),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_279),
.A2(n_242),
.B(n_70),
.Y(n_360)
);

CKINVDCx10_ASAP7_75t_R g361 ( 
.A(n_303),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_272),
.B(n_313),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_277),
.B(n_7),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

AOI221xp5_ASAP7_75t_L g365 ( 
.A1(n_310),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_314),
.Y(n_366)
);

OA22x2_ASAP7_75t_L g367 ( 
.A1(n_293),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_314),
.B(n_11),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_269),
.A2(n_71),
.B(n_124),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_278),
.B(n_12),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_69),
.B(n_122),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_301),
.B(n_13),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_304),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_305),
.A2(n_73),
.B1(n_120),
.B2(n_25),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_318),
.A2(n_75),
.B(n_27),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_311),
.B(n_28),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_77),
.B(n_30),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_SL g382 ( 
.A1(n_325),
.A2(n_326),
.B(n_309),
.C(n_308),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_326),
.A2(n_81),
.B(n_31),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_286),
.A2(n_84),
.B1(n_32),
.B2(n_33),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_294),
.B(n_85),
.Y(n_385)
);

AO31x2_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_17),
.A3(n_34),
.B(n_36),
.Y(n_386)
);

AO32x2_ASAP7_75t_L g387 ( 
.A1(n_331),
.A2(n_37),
.A3(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_387)
);

AOI221x1_ASAP7_75t_L g388 ( 
.A1(n_333),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.C(n_49),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_50),
.Y(n_389)
);

AO31x2_ASAP7_75t_L g390 ( 
.A1(n_368),
.A2(n_51),
.A3(n_52),
.B(n_53),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_334),
.B(n_54),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_332),
.B(n_55),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_58),
.B(n_59),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_60),
.B(n_61),
.Y(n_395)
);

AOI21x1_ASAP7_75t_L g396 ( 
.A1(n_335),
.A2(n_62),
.B(n_63),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_L g397 ( 
.A1(n_345),
.A2(n_64),
.B(n_67),
.Y(n_397)
);

OAI21x1_ASAP7_75t_SL g398 ( 
.A1(n_371),
.A2(n_72),
.B(n_76),
.Y(n_398)
);

NAND3x1_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_86),
.C(n_88),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_366),
.A2(n_91),
.B(n_92),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_93),
.Y(n_401)
);

AOI21xp33_ASAP7_75t_L g402 ( 
.A1(n_362),
.A2(n_337),
.B(n_351),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_328),
.A2(n_340),
.B(n_346),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_342),
.B(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_99),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_103),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_367),
.Y(n_409)
);

AOI21xp33_ASAP7_75t_L g410 ( 
.A1(n_358),
.A2(n_105),
.B(n_106),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_347),
.A2(n_355),
.B(n_382),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_356),
.B(n_108),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_110),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_348),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_364),
.B(n_114),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

AO31x2_ASAP7_75t_L g420 ( 
.A1(n_377),
.A2(n_118),
.A3(n_380),
.B(n_378),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_348),
.B(n_359),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_350),
.B(n_352),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_353),
.A2(n_357),
.B(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_338),
.B(n_375),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_376),
.Y(n_425)
);

BUFx4_ASAP7_75t_SL g426 ( 
.A(n_361),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_349),
.A2(n_370),
.B(n_360),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_375),
.B(n_376),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_375),
.B(n_384),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_381),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_385),
.A2(n_295),
.B(n_333),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g434 ( 
.A1(n_403),
.A2(n_423),
.B(n_412),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

AOI21x1_ASAP7_75t_L g437 ( 
.A1(n_432),
.A2(n_401),
.B(n_424),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_413),
.A2(n_402),
.B1(n_399),
.B2(n_389),
.Y(n_438)
);

AO21x2_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_392),
.B(n_394),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_SL g440 ( 
.A(n_408),
.B(n_419),
.Y(n_440)
);

BUFx2_ASAP7_75t_R g441 ( 
.A(n_426),
.Y(n_441)
);

INVx3_ASAP7_75t_SL g442 ( 
.A(n_419),
.Y(n_442)
);

NAND2x1_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_421),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_422),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

BUFx8_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_415),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_388),
.A2(n_397),
.B(n_396),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_395),
.A2(n_400),
.B(n_428),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_406),
.B(n_414),
.Y(n_457)
);

AO31x2_ASAP7_75t_L g458 ( 
.A1(n_416),
.A2(n_386),
.A3(n_420),
.B(n_387),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_407),
.B(n_393),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_433),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_433),
.A2(n_420),
.B(n_430),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_410),
.A2(n_386),
.B(n_387),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_386),
.A2(n_387),
.B(n_390),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_390),
.A2(n_412),
.B(n_328),
.Y(n_467)
);

BUFx8_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_404),
.B(n_288),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_402),
.B(n_413),
.Y(n_470)
);

OA21x2_ASAP7_75t_L g471 ( 
.A1(n_412),
.A2(n_328),
.B(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_432),
.A2(n_295),
.B(n_333),
.Y(n_474)
);

NOR2x1_ASAP7_75t_SL g475 ( 
.A(n_408),
.B(n_359),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_421),
.B(n_419),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_435),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_454),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_457),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_454),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_472),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_470),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_461),
.A2(n_434),
.B(n_474),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_438),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_445),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_456),
.A2(n_474),
.B(n_437),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_460),
.A2(n_471),
.B(n_457),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_436),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_445),
.B(n_453),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_452),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_476),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_459),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_467),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_465),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_476),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_458),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_466),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_444),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_455),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_439),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_488),
.A2(n_439),
.B1(n_464),
.B2(n_451),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_509),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_509),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_464),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_478),
.B(n_475),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_443),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_442),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_442),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_440),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_511),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_507),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_441),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_511),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g530 ( 
.A1(n_490),
.A2(n_468),
.B(n_450),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_450),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_468),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_508),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_441),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_481),
.A2(n_500),
.B1(n_499),
.B2(n_507),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_489),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_487),
.B(n_506),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_504),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_484),
.B(n_479),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_477),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_483),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_494),
.B(n_493),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_494),
.B(n_493),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_497),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_497),
.B(n_483),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_495),
.B(n_491),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_502),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_504),
.B(n_505),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_481),
.B(n_505),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_501),
.B(n_514),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_500),
.B(n_512),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_518),
.B(n_513),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_547),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_550),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_526),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_513),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_529),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_552),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_514),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_531),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_527),
.A2(n_500),
.B1(n_512),
.B2(n_489),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_552),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_556),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_531),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_557),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_557),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_538),
.B(n_486),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_526),
.B(n_489),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_550),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_534),
.B(n_486),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_548),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_537),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_548),
.B(n_551),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_523),
.B(n_498),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_486),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_542),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_515),
.B(n_530),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_534),
.Y(n_587)
);

AOI221xp5_ASAP7_75t_L g588 ( 
.A1(n_540),
.A2(n_498),
.B1(n_492),
.B2(n_490),
.C(n_486),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_553),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_542),
.B(n_492),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_524),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_519),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_580),
.B(n_519),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_571),
.B(n_539),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_539),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_563),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_525),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_590),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_573),
.B(n_516),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_560),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_589),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_565),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_559),
.B(n_528),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_559),
.B(n_528),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_589),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_582),
.B(n_549),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_582),
.B(n_523),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_564),
.B(n_525),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_564),
.B(n_517),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_585),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_522),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_573),
.B(n_522),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_568),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_576),
.B(n_530),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_575),
.B(n_517),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_584),
.B(n_554),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_572),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_587),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_574),
.B(n_521),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_584),
.B(n_554),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_613),
.A2(n_569),
.B(n_586),
.C(n_527),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_599),
.B(n_574),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_562),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_602),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_620),
.B(n_579),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_595),
.B(n_530),
.Y(n_631)
);

XOR2x2_ASAP7_75t_L g632 ( 
.A(n_609),
.B(n_535),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_595),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_597),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_579),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_621),
.B(n_567),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_593),
.B(n_562),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_621),
.B(n_567),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_594),
.B(n_587),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_600),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_591),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_605),
.B(n_562),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_603),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_634),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_641),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_626),
.A2(n_533),
.B(n_532),
.C(n_535),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_628),
.B(n_598),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_626),
.A2(n_614),
.B(n_624),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_632),
.A2(n_536),
.B1(n_586),
.B2(n_558),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_630),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_629),
.B(n_615),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_631),
.A2(n_618),
.B(n_608),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_627),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_629),
.B(n_598),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_647),
.B(n_619),
.C(n_623),
.Y(n_656)
);

AOI21xp33_ASAP7_75t_L g657 ( 
.A1(n_653),
.A2(n_631),
.B(n_640),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_654),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_645),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_652),
.B(n_638),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_646),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_651),
.B(n_637),
.Y(n_662)
);

NAND2x1_ASAP7_75t_L g663 ( 
.A(n_658),
.B(n_655),
.Y(n_663)
);

OAI21xp33_ASAP7_75t_L g664 ( 
.A1(n_656),
.A2(n_650),
.B(n_649),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_657),
.A2(n_651),
.B(n_633),
.C(n_642),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_659),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_660),
.B(n_661),
.Y(n_667)
);

NOR2xp67_ASAP7_75t_L g668 ( 
.A(n_666),
.B(n_662),
.Y(n_668)
);

AOI211xp5_ASAP7_75t_L g669 ( 
.A1(n_664),
.A2(n_521),
.B(n_558),
.C(n_577),
.Y(n_669)
);

NAND3x1_ASAP7_75t_L g670 ( 
.A(n_667),
.B(n_648),
.C(n_642),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_665),
.B(n_577),
.C(n_541),
.Y(n_671)
);

AOI211xp5_ASAP7_75t_L g672 ( 
.A1(n_663),
.A2(n_558),
.B(n_592),
.C(n_520),
.Y(n_672)
);

AOI211x1_ASAP7_75t_L g673 ( 
.A1(n_671),
.A2(n_639),
.B(n_637),
.C(n_596),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_672),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_669),
.B(n_643),
.Y(n_675)
);

NAND3x1_ASAP7_75t_L g676 ( 
.A(n_675),
.B(n_670),
.C(n_639),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_674),
.A2(n_618),
.B1(n_636),
.B2(n_644),
.C(n_520),
.Y(n_677)
);

AOI221xp5_ASAP7_75t_L g678 ( 
.A1(n_673),
.A2(n_644),
.B1(n_611),
.B2(n_604),
.C(n_622),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_675),
.Y(n_679)
);

XOR2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_555),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_676),
.B(n_596),
.Y(n_681)
);

NAND4xp25_ASAP7_75t_L g682 ( 
.A(n_677),
.B(n_555),
.C(n_588),
.D(n_543),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_678),
.Y(n_683)
);

NOR2x1p5_ASAP7_75t_L g684 ( 
.A(n_679),
.B(n_635),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_679),
.Y(n_685)
);

AO22x2_ASAP7_75t_L g686 ( 
.A1(n_683),
.A2(n_546),
.B1(n_616),
.B2(n_617),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_685),
.A2(n_561),
.B1(n_578),
.B2(n_601),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_685),
.Y(n_688)
);

XNOR2xp5_ASAP7_75t_L g689 ( 
.A(n_684),
.B(n_576),
.Y(n_689)
);

XNOR2x1_ASAP7_75t_L g690 ( 
.A(n_680),
.B(n_541),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_681),
.A2(n_625),
.B1(n_612),
.B2(n_610),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_688),
.B(n_682),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_686),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_687),
.A2(n_541),
.B1(n_610),
.B2(n_606),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_691),
.A2(n_607),
.B1(n_541),
.B2(n_606),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_693),
.B(n_689),
.Y(n_696)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_695),
.A2(n_690),
.B(n_607),
.Y(n_697)
);

XNOR2xp5_ASAP7_75t_L g698 ( 
.A(n_694),
.B(n_576),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_692),
.A2(n_541),
.B1(n_570),
.B2(n_566),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_612),
.B(n_605),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_698),
.A2(n_581),
.B1(n_570),
.B2(n_566),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_700),
.A2(n_697),
.B(n_699),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_591),
.C(n_545),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_702),
.A2(n_545),
.B(n_544),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_704),
.A2(n_703),
.B1(n_581),
.B2(n_544),
.Y(n_705)
);


endmodule