module fake_jpeg_22881_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.C(n_1),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_14),
.B(n_15),
.Y(n_20)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

AOI21xp33_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_18),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_11),
.B1(n_8),
.B2(n_2),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_8),
.B(n_12),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_27),
.B(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_15),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_30),
.B1(n_19),
.B2(n_5),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_19),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_26),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_34),
.C(n_33),
.Y(n_36)
);


endmodule