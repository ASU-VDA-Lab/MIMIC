module fake_ibex_1374_n_1930 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_1930);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_1930;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_504;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_1036;
wire n_974;
wire n_1831;
wire n_608;
wire n_864;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_878;
wire n_474;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1894;
wire n_961;
wire n_634;
wire n_1331;
wire n_1349;
wire n_991;
wire n_1223;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_423;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_1928;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1900;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_9),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_306),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_138),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_293),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_236),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_105),
.Y(n_418)
);

BUFx2_ASAP7_75t_SL g419 ( 
.A(n_394),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_23),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_323),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_96),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_314),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_4),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_343),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_346),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_352),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_23),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_120),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_241),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_225),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_324),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_327),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_18),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_295),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_255),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_8),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_407),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_402),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_300),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_251),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_288),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_28),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_332),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_90),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_30),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_175),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_357),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_379),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_205),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_294),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_315),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_319),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_309),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_32),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_256),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_356),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_335),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_214),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_162),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_17),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_122),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_90),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_85),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_54),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_354),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_57),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_208),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_70),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_230),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_393),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_15),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_382),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_270),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_49),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_32),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_301),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_186),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_21),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_53),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_68),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_291),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_72),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_68),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_333),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_19),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_97),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_163),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_289),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_365),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_52),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_311),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_296),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_74),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_184),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_336),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_137),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_259),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_131),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_199),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_140),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_108),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_351),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_18),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_409),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_286),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_238),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_227),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_272),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_396),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_223),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_363),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_292),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_312),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_104),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_339),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_371),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_235),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_250),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_326),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_318),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_387),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_349),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_395),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_317),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_374),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_231),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_252),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_405),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_207),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_340),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_61),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_329),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_384),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_211),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_342),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_216),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_322),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_98),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_105),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_167),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_248),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_358),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_362),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_258),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_96),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_174),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_16),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_341),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_313),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_298),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_284),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_117),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_165),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_287),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_350),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_260),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_147),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_360),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_280),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_321),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_228),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_53),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_242),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_74),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_316),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_247),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_117),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_120),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_367),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_347),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_397),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_93),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_299),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_121),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_244),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_388),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_310),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_253),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_157),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_361),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_337),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_106),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_274),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_403),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_85),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_121),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_148),
.Y(n_593)
);

BUFx5_ASAP7_75t_L g594 ( 
.A(n_386),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_348),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_2),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_159),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_304),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_297),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_385),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_40),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_239),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_49),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_217),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_201),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_12),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_375),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_123),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_62),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_113),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_122),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_331),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_139),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_380),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_369),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_33),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_328),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_263),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_0),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_104),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_188),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_80),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_7),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_408),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_404),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_206),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_392),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_142),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_376),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_41),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_302),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_25),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_308),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_218),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_364),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_372),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_325),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_209),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_285),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_282),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_29),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_200),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_278),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_52),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_307),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_13),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_70),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_132),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_330),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_73),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_283),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_158),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_203),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_305),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_273),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_257),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_249),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_193),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_377),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_212),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_320),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_366),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_98),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_368),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_303),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_54),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_79),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_411),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_389),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_400),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_391),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_370),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_399),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_179),
.Y(n_674)
);

BUFx5_ASAP7_75t_L g675 ( 
.A(n_338),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_43),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_47),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_91),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_189),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_213),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_373),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_78),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_197),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_398),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_118),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_355),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_48),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_204),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_103),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_38),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_160),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_46),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_345),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_390),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_378),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_65),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_344),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_47),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_28),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_196),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_84),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_134),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_383),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_125),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_22),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_359),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_59),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_30),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_495),
.B(n_0),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_555),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_499),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_530),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_494),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_490),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_681),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_424),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_473),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_481),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_702),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_591),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_591),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_490),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_650),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_650),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_689),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_689),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_528),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_467),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_472),
.B(n_1),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_565),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_708),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_497),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_426),
.B(n_1),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_708),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_597),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_430),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_698),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_698),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_701),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_701),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_578),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_655),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_497),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_632),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_429),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_447),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_465),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_466),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_475),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_487),
.Y(n_751)
);

BUFx2_ASAP7_75t_SL g752 ( 
.A(n_459),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_489),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_519),
.B(n_2),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_573),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_570),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_459),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_588),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_574),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_574),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_427),
.B(n_3),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_592),
.Y(n_762)
);

CKINVDCx14_ASAP7_75t_R g763 ( 
.A(n_434),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_601),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_540),
.B(n_3),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_608),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_L g767 ( 
.A(n_609),
.B(n_4),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_610),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_R g769 ( 
.A(n_414),
.B(n_126),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_620),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_630),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_641),
.Y(n_772)
);

INVxp33_ASAP7_75t_SL g773 ( 
.A(n_430),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_666),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_667),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_480),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_676),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_574),
.Y(n_778)
);

INVxp33_ASAP7_75t_SL g779 ( 
.A(n_413),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_677),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_480),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_418),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_690),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_570),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_692),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_547),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_434),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_682),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_594),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_434),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_584),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_584),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_547),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_590),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_590),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_631),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_584),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_631),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_688),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_640),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_594),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_420),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_688),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_688),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_421),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_454),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_440),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_454),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_714),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_789),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_742),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_806),
.B(n_579),
.Y(n_812)
);

AND2x6_ASAP7_75t_L g813 ( 
.A(n_787),
.B(n_455),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_745),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_752),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_789),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_801),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_720),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_714),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_757),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_776),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_721),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_723),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_724),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_725),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_726),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_735),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_808),
.B(n_561),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_801),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_790),
.B(n_705),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_738),
.Y(n_831)
);

INVx6_ASAP7_75t_L g832 ( 
.A(n_759),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_737),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_805),
.B(n_585),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_763),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_739),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_740),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_763),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_781),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_732),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_730),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_807),
.B(n_683),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_795),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_729),
.B(n_682),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_796),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_798),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_800),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_R g848 ( 
.A(n_716),
.B(n_640),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_741),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_746),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_791),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_782),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_794),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_747),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_748),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_749),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_751),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_773),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_786),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_753),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_755),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_758),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_792),
.B(n_561),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_722),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_762),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_764),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_797),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_766),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_768),
.B(n_441),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_770),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_771),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_774),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_780),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_783),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_802),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_785),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_786),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_765),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_793),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_734),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_722),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_793),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_744),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_744),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_713),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_750),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_734),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_799),
.B(n_522),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_713),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_803),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_772),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_804),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_717),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_775),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_777),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_756),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_718),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_728),
.B(n_682),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_778),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_761),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_727),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_761),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_709),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_754),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_731),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_767),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_736),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_709),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_760),
.B(n_707),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_710),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_711),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_743),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_756),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_712),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_784),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_715),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_719),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_788),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_769),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_779),
.B(n_455),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_769),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_784),
.B(n_453),
.C(n_442),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_733),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_789),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_714),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_806),
.B(n_423),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_752),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_742),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_752),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_752),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_720),
.B(n_533),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_789),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_742),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_789),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_789),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_789),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_714),
.Y(n_937)
);

INVx6_ASAP7_75t_L g938 ( 
.A(n_759),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_742),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_742),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_742),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_752),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_789),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_742),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_789),
.A2(n_477),
.B(n_441),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_737),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_789),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_752),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_752),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_789),
.A2(n_520),
.B(n_477),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_742),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_806),
.B(n_520),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_789),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_806),
.B(n_527),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_742),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_789),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_714),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_720),
.B(n_669),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_742),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_806),
.B(n_527),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_742),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_789),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_752),
.Y(n_963)
);

OA21x2_ASAP7_75t_L g964 ( 
.A1(n_789),
.A2(n_598),
.B(n_562),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_878),
.B(n_417),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_875),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_959),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_959),
.Y(n_968)
);

AO22x2_ASAP7_75t_L g969 ( 
.A1(n_922),
.A2(n_568),
.B1(n_703),
.B2(n_674),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_836),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_893),
.B(n_674),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_961),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_L g973 ( 
.A(n_813),
.B(n_594),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_961),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_841),
.B(n_436),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_811),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_836),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_814),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_836),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_848),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_830),
.B(n_703),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_830),
.B(n_425),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_828),
.B(n_900),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_835),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_837),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_916),
.A2(n_438),
.B1(n_445),
.B2(n_435),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_885),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_899),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_837),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_910),
.B(n_448),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_837),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_832),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_832),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_894),
.B(n_415),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_838),
.B(n_458),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_852),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_895),
.B(n_416),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_920),
.B(n_464),
.Y(n_998)
);

OAI22x1_ASAP7_75t_L g999 ( 
.A1(n_859),
.A2(n_468),
.B1(n_478),
.B2(n_470),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_928),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_920),
.B(n_479),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_933),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_938),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_889),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_918),
.B(n_474),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_831),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_849),
.Y(n_1007)
);

AND2x6_ASAP7_75t_L g1008 ( 
.A(n_902),
.B(n_485),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_851),
.B(n_476),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_867),
.B(n_482),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_880),
.B(n_422),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_858),
.B(n_483),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_945),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_922),
.B(n_486),
.C(n_484),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_851),
.B(n_496),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_833),
.B(n_506),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_886),
.B(n_525),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_939),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_940),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_880),
.B(n_428),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_941),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_944),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_950),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_844),
.B(n_485),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_853),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_816),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_938),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_926),
.B(n_431),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_890),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_892),
.B(n_432),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_815),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_951),
.Y(n_1032)
);

NAND3xp33_ASAP7_75t_L g1033 ( 
.A(n_946),
.B(n_537),
.C(n_508),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_955),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_816),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_898),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_818),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_891),
.A2(n_419),
.B1(n_469),
.B2(n_457),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_822),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_816),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_909),
.B(n_503),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_911),
.B(n_914),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_823),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_850),
.B(n_433),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_840),
.B(n_544),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_964),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_824),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_825),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_880),
.B(n_437),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_826),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_855),
.B(n_439),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_856),
.B(n_443),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_817),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_827),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_854),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_927),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_862),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_865),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_964),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_872),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_887),
.B(n_444),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_857),
.B(n_860),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_817),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_817),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_929),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_930),
.Y(n_1066)
);

BUFx4_ASAP7_75t_L g1067 ( 
.A(n_917),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_876),
.B(n_545),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_861),
.B(n_446),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_863),
.B(n_552),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_866),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_868),
.B(n_551),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_935),
.Y(n_1073)
);

AND2x6_ASAP7_75t_L g1074 ( 
.A(n_887),
.B(n_503),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_931),
.B(n_553),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_870),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_871),
.Y(n_1077)
);

BUFx10_ASAP7_75t_L g1078 ( 
.A(n_942),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_923),
.Y(n_1079)
);

AND2x6_ASAP7_75t_L g1080 ( 
.A(n_887),
.B(n_514),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_935),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_903),
.B(n_908),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_948),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_873),
.B(n_558),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_874),
.B(n_580),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_869),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_903),
.A2(n_492),
.B1(n_498),
.B2(n_491),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_935),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_812),
.B(n_449),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_963),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_869),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_952),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_820),
.B(n_596),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_897),
.B(n_603),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_956),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_888),
.B(n_635),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_952),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_956),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_954),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_903),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_954),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_901),
.B(n_606),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_809),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_960),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_821),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_956),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_812),
.B(n_450),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_960),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_904),
.Y(n_1110)
);

AO22x2_ASAP7_75t_L g1111 ( 
.A1(n_906),
.A2(n_505),
.B1(n_507),
.B2(n_501),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_834),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_834),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_931),
.B(n_958),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_810),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_842),
.Y(n_1116)
);

INVxp33_ASAP7_75t_L g1117 ( 
.A(n_908),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_908),
.A2(n_616),
.B1(n_619),
.B2(n_611),
.Y(n_1118)
);

BUFx10_ASAP7_75t_L g1119 ( 
.A(n_905),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_842),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_819),
.Y(n_1121)
);

AO22x2_ASAP7_75t_L g1122 ( 
.A1(n_877),
.A2(n_521),
.B1(n_524),
.B2(n_511),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_839),
.B(n_622),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_907),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_912),
.B(n_623),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_958),
.B(n_451),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_843),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_919),
.B(n_452),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_813),
.A2(n_535),
.B1(n_539),
.B2(n_538),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_921),
.B(n_456),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_829),
.B(n_460),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_813),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_924),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_932),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_845),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_813),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_846),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_934),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_847),
.B(n_644),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_936),
.B(n_514),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_943),
.B(n_461),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_864),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_947),
.B(n_462),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_879),
.B(n_646),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_953),
.B(n_463),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_962),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_962),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_962),
.B(n_471),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_882),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_881),
.B(n_647),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_883),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_957),
.B(n_488),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_884),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_896),
.B(n_493),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_913),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_915),
.B(n_500),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_925),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_937),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_836),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_959),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_959),
.Y(n_1161)
);

NAND3x1_ASAP7_75t_L g1162 ( 
.A(n_809),
.B(n_554),
.C(n_549),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_832),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_832),
.B(n_567),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_836),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_916),
.A2(n_685),
.B1(n_687),
.B2(n_678),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_875),
.B(n_696),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_899),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_832),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_959),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_841),
.B(n_502),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_878),
.B(n_504),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_959),
.Y(n_1173)
);

AND2x6_ASAP7_75t_L g1174 ( 
.A(n_841),
.B(n_571),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_959),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_878),
.B(n_509),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_841),
.B(n_699),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_832),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_878),
.B(n_510),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_836),
.Y(n_1180)
);

INVx8_ASAP7_75t_L g1181 ( 
.A(n_815),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_841),
.B(n_512),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_836),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_841),
.B(n_513),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_878),
.B(n_515),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_875),
.B(n_571),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_878),
.B(n_516),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_959),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_979),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1112),
.A2(n_1116),
.B1(n_1120),
.B2(n_1113),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1086),
.B(n_517),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_SL g1192 ( 
.A(n_1025),
.B(n_523),
.C(n_518),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_966),
.B(n_529),
.C(n_526),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_996),
.B(n_531),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1092),
.B(n_532),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1093),
.A2(n_586),
.B1(n_599),
.B2(n_593),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_996),
.B(n_5),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1167),
.B(n_5),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1098),
.B(n_534),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_988),
.B(n_1168),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1100),
.B(n_536),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1013),
.A2(n_983),
.B(n_1062),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_984),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1177),
.B(n_6),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1163),
.B(n_605),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1102),
.Y(n_1206)
);

AO22x1_ASAP7_75t_L g1207 ( 
.A1(n_1127),
.A2(n_542),
.B1(n_543),
.B2(n_541),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1105),
.B(n_546),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1109),
.A2(n_602),
.B1(n_604),
.B2(n_600),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_SL g1210 ( 
.A(n_971),
.B(n_548),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1034),
.B(n_1042),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1067),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_976),
.A2(n_613),
.B1(n_615),
.B2(n_607),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_965),
.B(n_550),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_975),
.B(n_556),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1068),
.B(n_557),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_L g1217 ( 
.A(n_1174),
.B(n_594),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_979),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1177),
.A2(n_617),
.B1(n_627),
.B2(n_624),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1071),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_978),
.B(n_559),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_979),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1000),
.A2(n_648),
.B1(n_657),
.B2(n_633),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1010),
.B(n_560),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1124),
.B(n_563),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1036),
.B(n_564),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1010),
.B(n_706),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1076),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1077),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1002),
.B(n_566),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1180),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1018),
.A2(n_661),
.B(n_664),
.C(n_660),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1014),
.A2(n_679),
.B1(n_691),
.B2(n_673),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1019),
.A2(n_697),
.B(n_695),
.C(n_598),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1136),
.B(n_1176),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1185),
.B(n_569),
.Y(n_1236)
);

AND2x6_ASAP7_75t_SL g1237 ( 
.A(n_1151),
.B(n_6),
.Y(n_1237)
);

NOR3xp33_ASAP7_75t_L g1238 ( 
.A(n_1142),
.B(n_575),
.C(n_572),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1021),
.A2(n_652),
.B1(n_562),
.B2(n_594),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_981),
.B(n_1127),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_993),
.Y(n_1241)
);

O2A1O1Ixp5_ASAP7_75t_L g1242 ( 
.A1(n_1011),
.A2(n_652),
.B(n_605),
.C(n_634),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_998),
.B(n_576),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1180),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_992),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_981),
.Y(n_1246)
);

BUFx4f_ASAP7_75t_L g1247 ( 
.A(n_1181),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1187),
.B(n_577),
.Y(n_1248)
);

NOR3xp33_ASAP7_75t_L g1249 ( 
.A(n_1152),
.B(n_582),
.C(n_581),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1111),
.A2(n_634),
.B1(n_675),
.B2(n_594),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1022),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1032),
.B(n_583),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_998),
.B(n_587),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1111),
.A2(n_594),
.B1(n_675),
.B2(n_595),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1037),
.Y(n_1255)
);

AND2x2_ASAP7_75t_SL g1256 ( 
.A(n_1106),
.B(n_7),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_990),
.A2(n_675),
.B1(n_612),
.B2(n_614),
.Y(n_1257)
);

NOR2x2_ASAP7_75t_L g1258 ( 
.A(n_1164),
.B(n_1104),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1180),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1072),
.B(n_589),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_990),
.B(n_8),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1066),
.B(n_704),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1084),
.B(n_618),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1119),
.B(n_621),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1101),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1001),
.B(n_625),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1039),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1001),
.B(n_626),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1043),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1119),
.B(n_628),
.Y(n_1270)
);

INVx4_ASAP7_75t_L g1271 ( 
.A(n_984),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1090),
.B(n_700),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_982),
.A2(n_675),
.B1(n_636),
.B2(n_637),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1085),
.B(n_629),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1164),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1172),
.B(n_1179),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1089),
.B(n_638),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_SL g1278 ( 
.A1(n_1070),
.A2(n_642),
.B(n_643),
.C(n_639),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1121),
.A2(n_649),
.B1(n_651),
.B2(n_645),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1056),
.B(n_1065),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_982),
.A2(n_675),
.B1(n_654),
.B2(n_656),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1031),
.B(n_1091),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1101),
.A2(n_675),
.B1(n_658),
.B2(n_659),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1108),
.B(n_653),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1047),
.B(n_662),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1056),
.B(n_9),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1065),
.B(n_694),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1083),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1082),
.A2(n_675),
.B1(n_668),
.B2(n_670),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1023),
.A2(n_671),
.B(n_665),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1082),
.A2(n_680),
.B1(n_684),
.B2(n_672),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1048),
.B(n_686),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1012),
.B(n_693),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1050),
.B(n_10),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1017),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1016),
.B(n_11),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1054),
.B(n_13),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1055),
.B(n_14),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1156),
.B(n_14),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1181),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_993),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1058),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1060),
.B(n_15),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1174),
.B(n_16),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1079),
.B(n_1024),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1083),
.B(n_17),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_967),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1174),
.B(n_19),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1169),
.Y(n_1309)
);

INVx8_ASAP7_75t_L g1310 ( 
.A(n_1074),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1178),
.Y(n_1311)
);

AND2x6_ASAP7_75t_L g1312 ( 
.A(n_1132),
.B(n_127),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1006),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_968),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1135),
.B(n_20),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_969),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1045),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1057),
.B(n_24),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1129),
.B(n_26),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1157),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1007),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_972),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_995),
.B(n_27),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1117),
.B(n_27),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1186),
.B(n_29),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_974),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1160),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1094),
.B(n_31),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_SL g1329 ( 
.A(n_1137),
.B(n_31),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1161),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1170),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_969),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_SL g1333 ( 
.A(n_1178),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1173),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1147),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1175),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1123),
.B(n_34),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_980),
.B(n_35),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1029),
.B(n_36),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1023),
.A2(n_129),
.B(n_128),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1122),
.A2(n_1188),
.B1(n_1133),
.B2(n_1138),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1027),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1009),
.B(n_36),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1114),
.B(n_37),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1110),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1078),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1149),
.B(n_37),
.Y(n_1347)
);

INVx8_ASAP7_75t_L g1348 ( 
.A(n_1074),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1115),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1153),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1015),
.B(n_39),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1095),
.B(n_41),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1041),
.B(n_42),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1075),
.B(n_42),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1075),
.B(n_43),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1103),
.B(n_44),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1040),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1008),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1038),
.B(n_1114),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1005),
.A2(n_1134),
.B(n_1097),
.C(n_973),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_994),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1008),
.B(n_45),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1008),
.B(n_48),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1078),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1155),
.Y(n_1365)
);

NOR3xp33_ASAP7_75t_L g1366 ( 
.A(n_1157),
.B(n_50),
.C(n_51),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_997),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1044),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1028),
.B(n_1118),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_986),
.B(n_50),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1166),
.B(n_51),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1146),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1046),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1051),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1052),
.B(n_55),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1003),
.B(n_55),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1069),
.B(n_56),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1040),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1125),
.B(n_56),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1171),
.B(n_1182),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1206),
.Y(n_1381)
);

AOI211xp5_ASAP7_75t_L g1382 ( 
.A1(n_1356),
.A2(n_1379),
.B(n_1366),
.C(n_1296),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1247),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1220),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1247),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1240),
.A2(n_1122),
.B1(n_1139),
.B2(n_1144),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1245),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1228),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1229),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1251),
.Y(n_1390)
);

AO22x1_ASAP7_75t_L g1391 ( 
.A1(n_1212),
.A2(n_1004),
.B1(n_987),
.B2(n_1074),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1346),
.B(n_1184),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1310),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1200),
.B(n_1150),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1300),
.B(n_1346),
.Y(n_1395)
);

BUFx2_ASAP7_75t_SL g1396 ( 
.A(n_1300),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1246),
.A2(n_999),
.B1(n_1033),
.B2(n_1154),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1357),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1255),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1320),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1225),
.B(n_1030),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1276),
.A2(n_1087),
.B(n_1126),
.C(n_1130),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1267),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1275),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1190),
.A2(n_1059),
.B1(n_1046),
.B2(n_1162),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1333),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1264),
.B(n_1270),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1269),
.B(n_1080),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1307),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1314),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1309),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1368),
.B(n_1080),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1342),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1288),
.B(n_1143),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1322),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1329),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1256),
.B(n_1158),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1331),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1374),
.B(n_1080),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1336),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1361),
.B(n_1128),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1367),
.B(n_1020),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1211),
.B(n_1049),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1302),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1326),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1357),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1378),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_SL g1428 ( 
.A(n_1193),
.B(n_1061),
.C(n_1131),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1376),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1327),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1320),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1310),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1341),
.B(n_1145),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1330),
.Y(n_1434)
);

OR2x2_ASAP7_75t_SL g1435 ( 
.A(n_1258),
.B(n_1059),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1345),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1334),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1310),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1341),
.B(n_1140),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1365),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1348),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1313),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1294),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1197),
.B(n_1141),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1297),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1194),
.B(n_1040),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1348),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1241),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1364),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1376),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1378),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1305),
.A2(n_1140),
.B1(n_1148),
.B2(n_977),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1321),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1280),
.B(n_970),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1298),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1348),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1198),
.B(n_1140),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1335),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1202),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1373),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1303),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1350),
.B(n_985),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1189),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1359),
.A2(n_1023),
.B1(n_1096),
.B2(n_1081),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1318),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1282),
.B(n_1096),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1203),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1344),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1301),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1344),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1218),
.Y(n_1471)
);

NOR3xp33_ASAP7_75t_SL g1472 ( 
.A(n_1210),
.B(n_57),
.C(n_58),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1339),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1204),
.B(n_1096),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1261),
.B(n_989),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_R g1476 ( 
.A(n_1333),
.B(n_58),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1315),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1203),
.B(n_1081),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1271),
.Y(n_1479)
);

BUFx8_ASAP7_75t_L g1480 ( 
.A(n_1311),
.Y(n_1480)
);

CKINVDCx16_ASAP7_75t_R g1481 ( 
.A(n_1376),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1325),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1271),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1237),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1349),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1355),
.Y(n_1486)
);

NOR3xp33_ASAP7_75t_SL g1487 ( 
.A(n_1224),
.B(n_59),
.C(n_60),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1323),
.A2(n_1293),
.B1(n_1337),
.B2(n_1328),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1282),
.B(n_1081),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1222),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1231),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1316),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1316),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1352),
.B(n_991),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1335),
.Y(n_1495)
);

AND3x1_ASAP7_75t_L g1496 ( 
.A(n_1192),
.B(n_1165),
.C(n_1159),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1219),
.B(n_1183),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1244),
.Y(n_1498)
);

NOR3xp33_ASAP7_75t_SL g1499 ( 
.A(n_1227),
.B(n_1253),
.C(n_1243),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1370),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1196),
.B(n_1099),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1279),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_L g1503 ( 
.A(n_1354),
.B(n_60),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1266),
.B(n_1026),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1205),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1209),
.B(n_1099),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1380),
.B(n_1035),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1286),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_R g1509 ( 
.A(n_1217),
.B(n_1312),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1213),
.B(n_1099),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1259),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1265),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1312),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1213),
.B(n_1053),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_R g1515 ( 
.A(n_1312),
.B(n_61),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1223),
.B(n_1063),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1223),
.B(n_1107),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1369),
.A2(n_1073),
.B(n_1064),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1312),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_L g1520 ( 
.A(n_1265),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1372),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1371),
.Y(n_1522)
);

NOR2xp67_ASAP7_75t_L g1523 ( 
.A(n_1268),
.B(n_62),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1272),
.B(n_1088),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1207),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1353),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1287),
.B(n_63),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1332),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1242),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1402),
.A2(n_1360),
.B(n_1232),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1459),
.A2(n_1377),
.B(n_1375),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1393),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1400),
.Y(n_1533)
);

INVx3_ASAP7_75t_SL g1534 ( 
.A(n_1383),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1500),
.A2(n_1208),
.B(n_1199),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1459),
.A2(n_1235),
.B(n_1343),
.Y(n_1536)
);

NOR2x1_ASAP7_75t_L g1537 ( 
.A(n_1396),
.B(n_1306),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1518),
.A2(n_1351),
.B(n_1340),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1387),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1513),
.A2(n_1239),
.B(n_1304),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1492),
.B(n_1299),
.Y(n_1541)
);

AO21x1_ASAP7_75t_L g1542 ( 
.A1(n_1405),
.A2(n_1362),
.B(n_1363),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1493),
.A2(n_1234),
.A3(n_1347),
.B(n_1308),
.Y(n_1543)
);

OA22x2_ASAP7_75t_L g1544 ( 
.A1(n_1528),
.A2(n_1324),
.B1(n_1239),
.B2(n_1262),
.Y(n_1544)
);

AO31x2_ASAP7_75t_L g1545 ( 
.A1(n_1464),
.A2(n_1290),
.A3(n_1195),
.B(n_1191),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1529),
.A2(n_1250),
.B(n_1254),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1381),
.B(n_1260),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1478),
.A2(n_1319),
.B(n_1358),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1384),
.Y(n_1549)
);

AO31x2_ASAP7_75t_L g1550 ( 
.A1(n_1461),
.A2(n_1230),
.A3(n_1252),
.B(n_1221),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1386),
.B(n_1226),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1381),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1422),
.B(n_1249),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1439),
.A2(n_1317),
.B(n_1295),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1470),
.A2(n_1257),
.B1(n_1281),
.B2(n_1273),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1384),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1403),
.Y(n_1557)
);

AOI211x1_ASAP7_75t_L g1558 ( 
.A1(n_1485),
.A2(n_1201),
.B(n_1248),
.C(n_1236),
.Y(n_1558)
);

NOR2x1_ASAP7_75t_L g1559 ( 
.A(n_1406),
.B(n_1338),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1394),
.B(n_1263),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1481),
.B(n_1413),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1388),
.B(n_1274),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1461),
.A2(n_1233),
.B(n_1285),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1389),
.B(n_1216),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1465),
.A2(n_1292),
.B(n_1284),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1488),
.A2(n_1508),
.B1(n_1450),
.B2(n_1429),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1463),
.A2(n_1289),
.B(n_1283),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1471),
.A2(n_1491),
.B(n_1490),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1509),
.A2(n_1278),
.B(n_1277),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1465),
.A2(n_1215),
.B(n_1214),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1435),
.A2(n_1291),
.B1(n_1238),
.B2(n_65),
.Y(n_1571)
);

O2A1O1Ixp5_ASAP7_75t_L g1572 ( 
.A1(n_1446),
.A2(n_133),
.B(n_135),
.C(n_130),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1406),
.B(n_63),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1498),
.A2(n_1511),
.B(n_1408),
.Y(n_1574)
);

AOI21xp33_ASAP7_75t_L g1575 ( 
.A1(n_1382),
.A2(n_64),
.B(n_66),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1417),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1522),
.A2(n_67),
.B(n_69),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1510),
.A2(n_141),
.B(n_136),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1501),
.A2(n_144),
.B(n_143),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1390),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1443),
.A2(n_72),
.B(n_69),
.C(n_71),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1482),
.A2(n_71),
.B(n_73),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1480),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1445),
.A2(n_75),
.B(n_76),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1506),
.A2(n_146),
.B(n_145),
.Y(n_1585)
);

AOI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1433),
.A2(n_150),
.B(n_149),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1455),
.A2(n_152),
.B(n_151),
.Y(n_1587)
);

CKINVDCx6p67_ASAP7_75t_R g1588 ( 
.A(n_1505),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1473),
.A2(n_154),
.B(n_153),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1399),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1480),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1473),
.A2(n_156),
.B(n_155),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1401),
.A2(n_1419),
.B(n_1412),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1514),
.A2(n_75),
.B(n_76),
.Y(n_1594)
);

BUFx12f_ASAP7_75t_L g1595 ( 
.A(n_1431),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1436),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1489),
.A2(n_164),
.B(n_161),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1486),
.A2(n_168),
.B(n_166),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1424),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1502),
.B(n_77),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1422),
.B(n_77),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1398),
.A2(n_170),
.B(n_169),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1453),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1398),
.A2(n_172),
.B(n_171),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1391),
.B(n_78),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1393),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1426),
.A2(n_176),
.B(n_173),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1515),
.B(n_79),
.Y(n_1608)
);

O2A1O1Ixp5_ASAP7_75t_SL g1609 ( 
.A1(n_1407),
.A2(n_290),
.B(n_410),
.C(n_406),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1444),
.B(n_80),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1426),
.A2(n_178),
.B(n_177),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1425),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1427),
.A2(n_181),
.B(n_180),
.Y(n_1613)
);

OAI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1472),
.A2(n_81),
.B(n_82),
.Y(n_1614)
);

BUFx4f_ASAP7_75t_SL g1615 ( 
.A(n_1449),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1468),
.B(n_1430),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1494),
.A2(n_183),
.B(n_182),
.Y(n_1617)
);

AO31x2_ASAP7_75t_L g1618 ( 
.A1(n_1516),
.A2(n_81),
.A3(n_82),
.B(n_83),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1517),
.A2(n_83),
.B(n_84),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1560),
.B(n_1612),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1549),
.B(n_1434),
.Y(n_1621)
);

AO21x1_ASAP7_75t_L g1622 ( 
.A1(n_1619),
.A2(n_1594),
.B(n_1584),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1539),
.B(n_1404),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1614),
.A2(n_1487),
.B(n_1416),
.C(n_1523),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1542),
.A2(n_1457),
.B(n_1503),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1532),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1603),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1541),
.A2(n_1484),
.B1(n_1476),
.B2(n_1397),
.C(n_1499),
.Y(n_1629)
);

OR2x6_ASAP7_75t_L g1630 ( 
.A(n_1605),
.B(n_1513),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1535),
.A2(n_1423),
.B1(n_1525),
.B2(n_1477),
.C(n_1421),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1601),
.A2(n_1513),
.B1(n_1519),
.B2(n_1527),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1574),
.A2(n_1451),
.B(n_1427),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1588),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1519),
.B1(n_1527),
.B2(n_1440),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1538),
.A2(n_1451),
.B(n_1456),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1531),
.A2(n_1519),
.B(n_1497),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1579),
.A2(n_1585),
.B(n_1578),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1586),
.A2(n_1456),
.B(n_1410),
.Y(n_1639)
);

AO31x2_ASAP7_75t_L g1640 ( 
.A1(n_1536),
.A2(n_1437),
.A3(n_1415),
.B(n_1418),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1558),
.B(n_1428),
.C(n_1526),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1532),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1603),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1601),
.A2(n_1442),
.B1(n_1420),
.B2(n_1409),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1549),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1576),
.A2(n_1467),
.B1(n_1469),
.B2(n_1448),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1551),
.A2(n_1504),
.B1(n_1414),
.B2(n_1392),
.Y(n_1647)
);

NOR2x1_ASAP7_75t_SL g1648 ( 
.A(n_1532),
.B(n_1393),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1552),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1557),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1580),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1573),
.A2(n_1467),
.B1(n_1474),
.B2(n_1479),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1587),
.A2(n_1496),
.B(n_1495),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1615),
.A2(n_1467),
.B1(n_1483),
.B2(n_1452),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1593),
.A2(n_1495),
.B(n_1458),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1544),
.A2(n_1392),
.B1(n_1462),
.B2(n_1454),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1530),
.A2(n_1460),
.B(n_1475),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1599),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1556),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1553),
.B(n_1385),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1590),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1561),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1596),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1582),
.A2(n_1577),
.B1(n_1566),
.B2(n_1608),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1665)
);

INVx11_ASAP7_75t_L g1666 ( 
.A(n_1595),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1630),
.B(n_1606),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1644),
.A2(n_1571),
.B1(n_1575),
.B2(n_1583),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1651),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_1634),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1666),
.Y(n_1672)
);

INVx6_ASAP7_75t_L g1673 ( 
.A(n_1630),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1649),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1644),
.A2(n_1610),
.B1(n_1547),
.B2(n_1563),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1632),
.A2(n_1540),
.B(n_1598),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1620),
.B(n_1600),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1664),
.A2(n_1563),
.B1(n_1553),
.B2(n_1565),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1664),
.A2(n_1570),
.B1(n_1537),
.B2(n_1555),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1661),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1632),
.A2(n_1581),
.B1(n_1559),
.B2(n_1564),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1630),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1639),
.A2(n_1609),
.B(n_1592),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1662),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1622),
.A2(n_1631),
.B1(n_1656),
.B2(n_1647),
.Y(n_1685)
);

NAND3x1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.B(n_1533),
.C(n_1616),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1638),
.A2(n_1604),
.B(n_1602),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_R g1688 ( 
.A(n_1626),
.B(n_1598),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1645),
.B(n_1606),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1663),
.B(n_1562),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1628),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1631),
.A2(n_1629),
.B1(n_1641),
.B2(n_1635),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1624),
.B(n_1534),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1623),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1660),
.A2(n_1395),
.B1(n_1466),
.B2(n_1554),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1659),
.B(n_1550),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1645),
.A2(n_1607),
.B1(n_1613),
.B2(n_1611),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1650),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1673),
.A2(n_1621),
.B1(n_1626),
.B2(n_1648),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1669),
.A2(n_1646),
.B1(n_1667),
.B2(n_1665),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1691),
.B(n_1695),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1670),
.B(n_1665),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1698),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1669),
.A2(n_1667),
.B1(n_1654),
.B2(n_1652),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1700),
.B(n_1658),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1680),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1674),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1685),
.A2(n_1625),
.B1(n_1621),
.B2(n_1657),
.C(n_1466),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1692),
.A2(n_1642),
.B1(n_1627),
.B2(n_1606),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1675),
.A2(n_1637),
.B(n_1657),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1694),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1692),
.A2(n_1686),
.B1(n_1684),
.B2(n_1685),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1677),
.B(n_1618),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1690),
.B(n_1618),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1633),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1679),
.A2(n_1627),
.B1(n_1642),
.B2(n_1458),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1679),
.A2(n_1589),
.B1(n_1637),
.B2(n_1617),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1696),
.B(n_1618),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1678),
.A2(n_1512),
.B(n_1411),
.C(n_1521),
.Y(n_1723)
);

OAI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1693),
.A2(n_1432),
.B1(n_1438),
.B2(n_1441),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1681),
.A2(n_1546),
.B1(n_1569),
.B2(n_1548),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1673),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1668),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1675),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1703),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1678),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1705),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1713),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1704),
.B(n_1676),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1701),
.B(n_1682),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1697),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1716),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1715),
.B(n_1707),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1703),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1709),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1708),
.B(n_1543),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1708),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1709),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1717),
.B(n_1673),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1716),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1714),
.A2(n_1668),
.B1(n_1699),
.B2(n_1636),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1722),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1722),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1718),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1727),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1718),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1718),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1728),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1732),
.Y(n_1753)
);

CKINVDCx12_ASAP7_75t_R g1754 ( 
.A(n_1737),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1741),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1732),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1730),
.A2(n_1745),
.B1(n_1734),
.B2(n_1735),
.Y(n_1757)
);

AND2x6_ASAP7_75t_SL g1758 ( 
.A(n_1730),
.B(n_1671),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1731),
.Y(n_1759)
);

AO22x1_ASAP7_75t_L g1760 ( 
.A1(n_1736),
.A2(n_1672),
.B1(n_1726),
.B2(n_1719),
.Y(n_1760)
);

AOI222xp33_ASAP7_75t_L g1761 ( 
.A1(n_1733),
.A2(n_1728),
.B1(n_1710),
.B2(n_1702),
.C1(n_1706),
.C2(n_1719),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1736),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1734),
.A2(n_1723),
.B(n_1724),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1752),
.B(n_1729),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1744),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1741),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1738),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_SL g1768 ( 
.A(n_1744),
.B(n_1672),
.Y(n_1768)
);

OAI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1743),
.A2(n_1711),
.B1(n_1725),
.B2(n_1726),
.C(n_1721),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1749),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1764),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1753),
.B(n_1748),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1757),
.B(n_1752),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1764),
.B(n_1737),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1756),
.B(n_1748),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1762),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1759),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1762),
.B(n_1750),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1756),
.B(n_1750),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1755),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1770),
.B(n_1751),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1765),
.Y(n_1782)
);

INVx5_ASAP7_75t_L g1783 ( 
.A(n_1758),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1766),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1761),
.B(n_1733),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1765),
.B(n_1735),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1760),
.B(n_1746),
.Y(n_1788)
);

OAI322xp33_ASAP7_75t_L g1789 ( 
.A1(n_1769),
.A2(n_1751),
.A3(n_1747),
.B1(n_1746),
.B2(n_1740),
.C1(n_1731),
.C2(n_1739),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1754),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1783),
.B(n_1768),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1786),
.B(n_1747),
.Y(n_1792)
);

NAND4xp25_ASAP7_75t_L g1793 ( 
.A(n_1790),
.B(n_1763),
.C(n_1769),
.D(n_1726),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1790),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1782),
.B(n_1720),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1774),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1774),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1771),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1791),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1796),
.Y(n_1800)
);

INVx5_ASAP7_75t_L g1801 ( 
.A(n_1793),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1797),
.B(n_1773),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1792),
.B(n_1783),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1802),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1800),
.Y(n_1805)
);

OAI32xp33_ASAP7_75t_L g1806 ( 
.A1(n_1803),
.A2(n_1794),
.A3(n_1782),
.B1(n_1776),
.B2(n_1788),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1799),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1805),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1806),
.B(n_1801),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1804),
.B(n_1801),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1810),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1809),
.B(n_1795),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1807),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1808),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1807),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1810),
.Y(n_1816)
);

AOI211x1_ASAP7_75t_L g1817 ( 
.A1(n_1810),
.A2(n_1798),
.B(n_1787),
.C(n_1783),
.Y(n_1817)
);

INVx8_ASAP7_75t_L g1818 ( 
.A(n_1816),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1813),
.B(n_1783),
.Y(n_1819)
);

OR3x1_ASAP7_75t_L g1820 ( 
.A(n_1815),
.B(n_1783),
.C(n_1785),
.Y(n_1820)
);

AOI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1811),
.A2(n_1789),
.B(n_1778),
.C(n_1779),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1814),
.B(n_1784),
.C(n_1438),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1812),
.B(n_1775),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1817),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1813),
.B(n_1775),
.Y(n_1825)
);

NAND2x1_ASAP7_75t_L g1826 ( 
.A(n_1812),
.B(n_1778),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1814),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1811),
.Y(n_1828)
);

A2O1A1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1824),
.A2(n_1779),
.B(n_1778),
.C(n_1520),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1828),
.A2(n_1520),
.B(n_1772),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1819),
.A2(n_1725),
.B1(n_1699),
.B2(n_1777),
.C(n_1780),
.Y(n_1831)
);

OAI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1818),
.A2(n_1438),
.B(n_1441),
.C(n_1432),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1818),
.B(n_1780),
.Y(n_1833)
);

A2O1A1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1827),
.A2(n_1822),
.B(n_1826),
.C(n_1825),
.Y(n_1834)
);

AOI321xp33_ASAP7_75t_L g1835 ( 
.A1(n_1823),
.A2(n_1772),
.A3(n_1781),
.B1(n_1777),
.B2(n_1524),
.C(n_1739),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1820),
.A2(n_1781),
.B1(n_1688),
.B2(n_1712),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1821),
.B(n_86),
.Y(n_1837)
);

OAI21xp33_ASAP7_75t_L g1838 ( 
.A1(n_1819),
.A2(n_1742),
.B(n_1441),
.Y(n_1838)
);

AOI221xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1828),
.A2(n_1447),
.B1(n_1432),
.B2(n_1742),
.C(n_89),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1818),
.A2(n_1712),
.B1(n_1524),
.B2(n_1447),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1828),
.A2(n_1572),
.B(n_1447),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1827),
.B(n_86),
.C(n_87),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1828),
.A2(n_1653),
.B(n_1597),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1818),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1824),
.A2(n_1687),
.B(n_1655),
.C(n_1683),
.Y(n_1845)
);

OAI221xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1828),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_91),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1844),
.B(n_88),
.Y(n_1847)
);

A2O1A1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1834),
.A2(n_1567),
.B(n_93),
.C(n_94),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1839),
.A2(n_1833),
.B1(n_1837),
.B2(n_1842),
.C(n_1838),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1832),
.A2(n_1688),
.B1(n_1712),
.B2(n_1546),
.Y(n_1850)
);

OAI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1846),
.A2(n_92),
.B(n_94),
.C(n_95),
.Y(n_1851)
);

XNOR2x1_ASAP7_75t_L g1852 ( 
.A(n_1830),
.B(n_92),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1841),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1831),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1829),
.B(n_1840),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_R g1856 ( 
.A(n_1835),
.B(n_95),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1845),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1836),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1843),
.A2(n_1568),
.B1(n_1460),
.B2(n_100),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1844),
.B(n_97),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1844),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1844),
.B(n_99),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_R g1863 ( 
.A(n_1844),
.B(n_99),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1847),
.B(n_100),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1861),
.B(n_1853),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1861),
.B(n_101),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1860),
.B(n_101),
.C(n_102),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_R g1868 ( 
.A(n_1862),
.B(n_102),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1858),
.B(n_103),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1863),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1851),
.A2(n_1460),
.B1(n_107),
.B2(n_108),
.Y(n_1871)
);

NOR2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1854),
.B(n_106),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1852),
.Y(n_1873)
);

NOR3xp33_ASAP7_75t_L g1874 ( 
.A(n_1848),
.B(n_107),
.C(n_109),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1857),
.B(n_109),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1859),
.B(n_110),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1855),
.B(n_110),
.Y(n_1877)
);

AND2x2_ASAP7_75t_SL g1878 ( 
.A(n_1849),
.B(n_111),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1856),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_1879)
);

OAI21xp33_ASAP7_75t_SL g1880 ( 
.A1(n_1850),
.A2(n_112),
.B(n_114),
.Y(n_1880)
);

INVxp33_ASAP7_75t_L g1881 ( 
.A(n_1861),
.Y(n_1881)
);

AND3x4_ASAP7_75t_L g1882 ( 
.A(n_1874),
.B(n_114),
.C(n_115),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1865),
.B(n_115),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1877),
.B(n_116),
.Y(n_1884)
);

NOR4xp25_ASAP7_75t_L g1885 ( 
.A(n_1870),
.B(n_116),
.C(n_118),
.D(n_119),
.Y(n_1885)
);

AOI211x1_ASAP7_75t_L g1886 ( 
.A1(n_1867),
.A2(n_119),
.B(n_123),
.C(n_124),
.Y(n_1886)
);

AOI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1881),
.A2(n_124),
.B1(n_1550),
.B2(n_1545),
.C(n_190),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1879),
.A2(n_1550),
.B1(n_1545),
.B2(n_1640),
.Y(n_1888)
);

NAND3xp33_ASAP7_75t_SL g1889 ( 
.A(n_1868),
.B(n_185),
.C(n_187),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1869),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1875),
.B(n_1545),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1866),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1872),
.B(n_1640),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1878),
.A2(n_1640),
.B1(n_192),
.B2(n_194),
.Y(n_1894)
);

CKINVDCx16_ASAP7_75t_R g1895 ( 
.A(n_1889),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1890),
.B(n_1873),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1885),
.B(n_1871),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1884),
.Y(n_1898)
);

INVx5_ASAP7_75t_L g1899 ( 
.A(n_1883),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1892),
.B(n_1864),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1886),
.Y(n_1901)
);

CKINVDCx20_ASAP7_75t_R g1902 ( 
.A(n_1891),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1893),
.B(n_1876),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1894),
.B(n_1880),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1882),
.A2(n_191),
.B1(n_195),
.B2(n_198),
.Y(n_1905)
);

NOR3xp33_ASAP7_75t_L g1906 ( 
.A(n_1887),
.B(n_202),
.C(n_210),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1901),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1896),
.Y(n_1908)
);

OAI22x1_ASAP7_75t_L g1909 ( 
.A1(n_1905),
.A2(n_1888),
.B1(n_219),
.B2(n_220),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1897),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1900),
.Y(n_1911)
);

OAI221xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1906),
.A2(n_215),
.B1(n_221),
.B2(n_222),
.C(n_224),
.Y(n_1912)
);

OAI22x1_ASAP7_75t_L g1913 ( 
.A1(n_1904),
.A2(n_226),
.B1(n_229),
.B2(n_232),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1898),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1908),
.B(n_1895),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1910),
.A2(n_1899),
.B(n_1903),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1911),
.Y(n_1917)
);

OAI22x1_ASAP7_75t_L g1918 ( 
.A1(n_1907),
.A2(n_1914),
.B1(n_1899),
.B2(n_1909),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1917),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1915),
.Y(n_1920)
);

OAI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1916),
.A2(n_1912),
.B1(n_1913),
.B2(n_1902),
.C(n_240),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1919),
.A2(n_1918),
.B(n_1920),
.Y(n_1922)
);

AOI21xp33_ASAP7_75t_L g1923 ( 
.A1(n_1921),
.A2(n_233),
.B(n_234),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1922),
.A2(n_237),
.B1(n_243),
.B2(n_245),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1923),
.A2(n_246),
.B(n_254),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1922),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1925),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1924),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_R g1929 ( 
.A1(n_1927),
.A2(n_1926),
.B1(n_275),
.B2(n_276),
.C(n_277),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1928),
.B1(n_279),
.B2(n_281),
.Y(n_1930)
);


endmodule