module real_jpeg_10863_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_3),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g32 ( 
.A(n_1),
.B(n_33),
.CON(n_32),
.SN(n_32)
);

HAxp5_ASAP7_75t_SL g35 ( 
.A(n_1),
.B(n_11),
.CON(n_35),
.SN(n_35)
);

AOI22xp5_ASAP7_75t_SL g9 ( 
.A1(n_2),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_9)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_13),
.Y(n_24)
);

OA21x2_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_16),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_4),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_11)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_18),
.B(n_28),
.C(n_36),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_15),
.B(n_17),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B(n_24),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_22),
.B(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_26),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_29),
.B(n_30),
.Y(n_28)
);

BUFx24_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);


endmodule