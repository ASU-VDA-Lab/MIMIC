module fake_jpeg_10883_n_536 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_536);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_1),
.B(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_66),
.Y(n_135)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_67),
.Y(n_156)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_103),
.Y(n_105)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_34),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_82),
.B(n_97),
.Y(n_139)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_38),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_87),
.B(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g164 ( 
.A(n_91),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_2),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_3),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_3),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_43),
.B(n_30),
.C(n_49),
.Y(n_127)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_22),
.B(n_3),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_50),
.B1(n_23),
.B2(n_52),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_147),
.B1(n_150),
.B2(n_25),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_66),
.A2(n_52),
.B1(n_37),
.B2(n_50),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_140),
.B1(n_151),
.B2(n_84),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_159),
.Y(n_185)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_132),
.Y(n_220)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_70),
.A2(n_50),
.B1(n_30),
.B2(n_20),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_36),
.B1(n_26),
.B2(n_29),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_74),
.A2(n_52),
.B1(n_37),
.B2(n_47),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_51),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_26),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_32),
.C(n_49),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_40),
.C(n_95),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_51),
.B1(n_25),
.B2(n_46),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_85),
.A2(n_36),
.B1(n_46),
.B2(n_45),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_57),
.A2(n_47),
.B1(n_32),
.B2(n_42),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_42),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_168),
.A2(n_176),
.B1(n_191),
.B2(n_122),
.Y(n_242)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

BUFx2_ASAP7_75t_SL g261 ( 
.A(n_169),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_94),
.B1(n_92),
.B2(n_89),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_164),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_179),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_181),
.Y(n_276)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_183),
.A2(n_188),
.B1(n_198),
.B2(n_118),
.Y(n_258)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_187),
.B(n_204),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_29),
.B1(n_40),
.B2(n_45),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_190),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_101),
.B1(n_77),
.B2(n_81),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_107),
.A2(n_58),
.B1(n_69),
.B2(n_59),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_226),
.B1(n_106),
.B2(n_114),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_140),
.A2(n_64),
.B1(n_91),
.B2(n_59),
.Y(n_196)
);

AO22x1_ASAP7_75t_SL g253 ( 
.A1(n_196),
.A2(n_214),
.B1(n_14),
.B2(n_15),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_135),
.A2(n_129),
.B(n_105),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_197),
.A2(n_11),
.B(n_13),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_130),
.A2(n_86),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_111),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_199),
.B(n_205),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_137),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_203),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_116),
.A2(n_86),
.B1(n_5),
.B2(n_7),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_201),
.A2(n_108),
.B1(n_136),
.B2(n_132),
.Y(n_244)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_125),
.A2(n_4),
.B(n_5),
.C(n_8),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_4),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_115),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_206),
.Y(n_280)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_218),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_126),
.B(n_8),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_213),
.B(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_9),
.Y(n_213)
);

AO22x2_ASAP7_75t_L g214 ( 
.A1(n_130),
.A2(n_18),
.B1(n_10),
.B2(n_11),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_18),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_9),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_219),
.Y(n_270)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_131),
.Y(n_221)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_9),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_227),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_110),
.Y(n_223)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_225),
.Y(n_273)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_120),
.B(n_10),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_133),
.B(n_11),
.C(n_13),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_228),
.B(n_217),
.CI(n_203),
.CON(n_272),
.SN(n_272)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_231),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_245),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_242),
.B1(n_276),
.B2(n_198),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_114),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_131),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_248),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_148),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_249),
.B(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_185),
.B(n_117),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_266),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_214),
.B1(n_196),
.B2(n_176),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_117),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_179),
.B(n_171),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_257),
.B(n_278),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_262),
.B1(n_220),
.B2(n_223),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_14),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_214),
.B(n_228),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_183),
.A2(n_118),
.B1(n_141),
.B2(n_128),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_128),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_196),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_141),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_214),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_168),
.A2(n_148),
.B1(n_15),
.B2(n_16),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_179),
.B(n_14),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_282),
.B(n_324),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_283),
.A2(n_235),
.B1(n_247),
.B2(n_234),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_284),
.A2(n_303),
.B(n_316),
.Y(n_355)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_232),
.A2(n_190),
.B(n_191),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_299),
.B(n_235),
.Y(n_343)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_298),
.B1(n_304),
.B2(n_318),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

BUFx24_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_294),
.Y(n_342)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_177),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_297),
.B(n_319),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_246),
.A2(n_173),
.B(n_216),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_310),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_305),
.Y(n_331)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

AOI32xp33_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_193),
.A3(n_226),
.B1(n_195),
.B2(n_175),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_276),
.B1(n_263),
.B2(n_253),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_209),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_309),
.B(n_312),
.Y(n_350)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_229),
.Y(n_310)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_315),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_236),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_317),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_243),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_266),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_248),
.B(n_221),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_259),
.A2(n_219),
.B1(n_215),
.B2(n_220),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_243),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_230),
.B(n_180),
.C(n_172),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_328),
.C(n_271),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_260),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_322),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_240),
.B(n_215),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_323),
.B(n_325),
.Y(n_335)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_245),
.B(n_169),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_329),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_253),
.A2(n_178),
.B1(n_170),
.B2(n_174),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_327),
.A2(n_261),
.B1(n_234),
.B2(n_233),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_245),
.B(n_193),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_250),
.B(n_17),
.Y(n_329)
);

XNOR2x2_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_259),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_330),
.A2(n_338),
.B(n_346),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_311),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_334),
.A2(n_344),
.B1(n_354),
.B2(n_318),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_301),
.A2(n_241),
.B1(n_237),
.B2(n_250),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_359),
.B1(n_363),
.B2(n_327),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_288),
.A2(n_247),
.B(n_260),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_343),
.A2(n_361),
.B(n_362),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_241),
.C(n_237),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_352),
.C(n_357),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_267),
.B(n_254),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_294),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_356),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_254),
.C(n_252),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_283),
.A2(n_279),
.B1(n_238),
.B2(n_252),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_294),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_238),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_298),
.A2(n_279),
.B1(n_269),
.B2(n_274),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_304),
.A2(n_280),
.B(n_274),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_316),
.A2(n_265),
.B(n_269),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_292),
.A2(n_265),
.B1(n_267),
.B2(n_17),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_15),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_368),
.A2(n_320),
.B(n_282),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_329),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_307),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_371),
.A2(n_404),
.B1(n_369),
.B2(n_337),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_328),
.C(n_286),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_380),
.C(n_383),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_366),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_353),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_377),
.Y(n_406)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_365),
.Y(n_376)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_370),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_378),
.Y(n_421)
);

XOR2x2_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_295),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_330),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_295),
.C(n_299),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_392),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_285),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_382),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_285),
.C(n_325),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_323),
.C(n_317),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_398),
.C(n_400),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_386),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_332),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_393),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_359),
.B1(n_361),
.B2(n_364),
.Y(n_426)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_391),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g392 ( 
.A1(n_331),
.A2(n_309),
.B(n_314),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_335),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_331),
.A2(n_306),
.B1(n_320),
.B2(n_287),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_395),
.A2(n_340),
.B1(n_363),
.B2(n_355),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_335),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_396),
.Y(n_411)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_356),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_289),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_399),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_324),
.C(n_313),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_350),
.A2(n_296),
.B(n_302),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_394),
.B(n_385),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_336),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_403),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_348),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_362),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_373),
.C(n_380),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_371),
.A2(n_334),
.B1(n_337),
.B2(n_354),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_410),
.A2(n_416),
.B1(n_419),
.B2(n_391),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_413),
.B(n_372),
.Y(n_436)
);

OAI22x1_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_344),
.B1(n_340),
.B2(n_355),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_414),
.Y(n_445)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_399),
.A2(n_350),
.B1(n_370),
.B2(n_348),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_395),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_426),
.A2(n_428),
.B(n_432),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_372),
.B(n_405),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_382),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_392),
.A2(n_330),
.B1(n_364),
.B2(n_347),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_430),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_381),
.A2(n_368),
.B(n_342),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_388),
.A2(n_358),
.B1(n_367),
.B2(n_360),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_436),
.B(n_444),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_456),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_398),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_440),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_384),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_415),
.Y(n_442)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_443),
.A2(n_460),
.B1(n_426),
.B2(n_433),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_383),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_452),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_400),
.C(n_379),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_455),
.C(n_459),
.Y(n_464)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_385),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_448),
.B(n_461),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_451),
.Y(n_467)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_413),
.Y(n_452)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_411),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_458),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_382),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_425),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_389),
.C(n_376),
.Y(n_459)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_408),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_440),
.B(n_446),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_465),
.B(n_470),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_410),
.B1(n_431),
.B2(n_423),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_472),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_459),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_439),
.B(n_414),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_441),
.A2(n_428),
.B(n_412),
.Y(n_474)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_R g475 ( 
.A(n_457),
.B(n_424),
.C(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_475),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_478),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_479),
.A2(n_453),
.B1(n_438),
.B2(n_386),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_437),
.B(n_425),
.C(n_424),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_482),
.C(n_455),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_449),
.A2(n_431),
.B1(n_423),
.B2(n_389),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_401),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_401),
.C(n_435),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_456),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_487),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_485),
.A2(n_339),
.B1(n_478),
.B2(n_471),
.Y(n_511)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

OAI221xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_452),
.B1(n_409),
.B2(n_397),
.C(n_402),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_489),
.A2(n_493),
.B1(n_496),
.B2(n_351),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_360),
.Y(n_490)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_490),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_409),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_495),
.C(n_498),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_421),
.B1(n_417),
.B2(n_358),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_462),
.B(n_421),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_469),
.A2(n_417),
.B1(n_367),
.B2(n_378),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_473),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_497),
.A2(n_342),
.B1(n_390),
.B2(n_366),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_368),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_488),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_501),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_476),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_502),
.Y(n_519)
);

OAI321xp33_ASAP7_75t_L g505 ( 
.A1(n_492),
.A2(n_481),
.A3(n_468),
.B1(n_475),
.B2(n_472),
.C(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_505),
.B(n_510),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_483),
.A2(n_494),
.B1(n_486),
.B2(n_491),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_508),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_466),
.B1(n_464),
.B2(n_477),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_498),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_484),
.B(n_464),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_511),
.A2(n_339),
.B1(n_291),
.B2(n_308),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_512),
.B(n_487),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_504),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_471),
.C(n_499),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_SL g522 ( 
.A(n_514),
.B(n_516),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_518),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_503),
.Y(n_525)
);

OAI21x1_ASAP7_75t_SL g527 ( 
.A1(n_522),
.A2(n_523),
.B(n_525),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_501),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_526),
.A2(n_521),
.B(n_514),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_524),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_529),
.B(n_516),
.Y(n_530)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_530),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_519),
.C(n_503),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_531),
.B(n_519),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_507),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_507),
.C(n_506),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_511),
.B1(n_16),
.B2(n_17),
.Y(n_536)
);


endmodule