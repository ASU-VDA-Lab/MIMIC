module fake_jpeg_12639_n_519 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_55),
.Y(n_111)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_65),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_0),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_78),
.Y(n_135)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_0),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_85),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_100),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_102),
.B(n_126),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_65),
.A2(n_18),
.B1(n_30),
.B2(n_42),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_108),
.A2(n_31),
.B1(n_84),
.B2(n_75),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_52),
.A2(n_18),
.B1(n_42),
.B2(n_23),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_119),
.A2(n_140),
.B1(n_157),
.B2(n_31),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_29),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_49),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_139),
.B(n_158),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_53),
.A2(n_23),
.B1(n_18),
.B2(n_46),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_62),
.B(n_50),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_141),
.B(n_154),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_98),
.B(n_27),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_62),
.B(n_25),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_164),
.Y(n_231)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_193),
.Y(n_225)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_169),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_192),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_177),
.B(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_49),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_121),
.B(n_111),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_205),
.C(n_183),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_114),
.B(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_183),
.B(n_196),
.Y(n_253)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_186),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_48),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_187),
.B(n_190),
.Y(n_259)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_48),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_122),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_45),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_45),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_127),
.A2(n_77),
.B1(n_97),
.B2(n_101),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g245 ( 
.A1(n_198),
.A2(n_143),
.B1(n_137),
.B2(n_155),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_117),
.B1(n_148),
.B2(n_128),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_40),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_215),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_140),
.A2(n_92),
.B1(n_94),
.B2(n_72),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_202),
.A2(n_203),
.B1(n_213),
.B2(n_51),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_105),
.B(n_88),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_212),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_33),
.C(n_40),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_130),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_123),
.B(n_33),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_145),
.A2(n_39),
.B1(n_85),
.B2(n_88),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_117),
.B1(n_128),
.B2(n_143),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_214),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_124),
.A2(n_64),
.B1(n_74),
.B2(n_73),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_134),
.B(n_39),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_124),
.B(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_3),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_248),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_219),
.A2(n_193),
.B1(n_179),
.B2(n_188),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_236),
.Y(n_277)
);

XNOR2x2_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_196),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_238),
.A2(n_193),
.B1(n_194),
.B2(n_192),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_191),
.A2(n_100),
.B(n_57),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_242),
.A2(n_11),
.B(n_12),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_68),
.B1(n_58),
.B2(n_66),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_202),
.B1(n_180),
.B2(n_169),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_54),
.C(n_150),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_244),
.B(n_10),
.Y(n_298)
);

AO21x2_ASAP7_75t_L g290 ( 
.A1(n_245),
.A2(n_252),
.B(n_5),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_204),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_198),
.A2(n_137),
.B1(n_155),
.B2(n_150),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_204),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_255),
.A2(n_12),
.B(n_14),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_268),
.A2(n_273),
.B1(n_222),
.B2(n_251),
.Y(n_337)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_176),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_270),
.B(n_271),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_200),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_215),
.B1(n_198),
.B2(n_205),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_272),
.B(n_278),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_168),
.B1(n_167),
.B2(n_163),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_290),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_229),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_162),
.B1(n_164),
.B2(n_186),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_160),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_282),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_242),
.A2(n_170),
.B1(n_181),
.B2(n_161),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_286),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_195),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_165),
.B(n_195),
.C(n_212),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_294),
.B(n_267),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_16),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_250),
.Y(n_287)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_296),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_227),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_228),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_234),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_297),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_258),
.B(n_230),
.C(n_236),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_7),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_295),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_225),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_258),
.Y(n_311)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_254),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_306),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_301),
.A2(n_260),
.B(n_263),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_225),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_264),
.B1(n_231),
.B2(n_232),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_224),
.B(n_11),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_293),
.C(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_15),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_311),
.B(n_321),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_316),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_313),
.A2(n_302),
.B(n_305),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_275),
.A2(n_264),
.B1(n_232),
.B2(n_261),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_290),
.A2(n_261),
.B1(n_256),
.B2(n_231),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_324),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_256),
.B1(n_220),
.B2(n_222),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_241),
.C(n_262),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_334),
.C(n_340),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_260),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_283),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_282),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_338),
.B(n_339),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_307),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_278),
.B(n_262),
.C(n_235),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_285),
.A2(n_239),
.B(n_218),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_344),
.A2(n_299),
.B(n_280),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_268),
.A2(n_218),
.B1(n_239),
.B2(n_235),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_276),
.B1(n_290),
.B2(n_308),
.Y(n_371)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

AO22x1_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_290),
.B1(n_288),
.B2(n_272),
.Y(n_354)
);

OAI31xp33_ASAP7_75t_SL g389 ( 
.A1(n_354),
.A2(n_309),
.A3(n_317),
.B(n_329),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_341),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_367),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_357),
.A2(n_378),
.B1(n_324),
.B2(n_315),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_286),
.Y(n_358)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_323),
.Y(n_361)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_301),
.B(n_285),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_362),
.A2(n_376),
.B(n_380),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_291),
.Y(n_363)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_298),
.C(n_294),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_327),
.C(n_318),
.Y(n_400)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_320),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_369),
.Y(n_387)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_265),
.A3(n_271),
.B1(n_279),
.B2(n_274),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_326),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_317),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_382),
.Y(n_411)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_287),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_312),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_328),
.A2(n_290),
.B1(n_300),
.B2(n_287),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_303),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_379),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_318),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_381),
.Y(n_398)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_331),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_384),
.C(n_396),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_311),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_368),
.A2(n_328),
.B1(n_333),
.B2(n_319),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_389),
.A2(n_354),
.B(n_357),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_350),
.A2(n_309),
.B1(n_319),
.B2(n_333),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_393),
.A2(n_410),
.B1(n_387),
.B2(n_408),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_317),
.B(n_315),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_394),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_321),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_336),
.C(n_314),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_400),
.C(n_351),
.Y(n_435)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_406),
.Y(n_423)
);

FAx1_ASAP7_75t_SL g401 ( 
.A(n_377),
.B(n_342),
.CI(n_343),
.CON(n_401),
.SN(n_401)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_369),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_327),
.C(n_348),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_383),
.C(n_384),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_370),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_403),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_358),
.B(n_335),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_407),
.B(n_393),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_350),
.A2(n_365),
.B1(n_356),
.B2(n_372),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_409),
.A2(n_399),
.B1(n_405),
.B2(n_389),
.Y(n_414)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_356),
.B1(n_373),
.B2(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_428),
.B1(n_433),
.B2(n_429),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_405),
.A2(n_363),
.B1(n_376),
.B2(n_362),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_430),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_404),
.A2(n_357),
.B(n_380),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_421),
.B(n_349),
.Y(n_457)
);

AOI21xp33_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_292),
.B(n_289),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_401),
.B(n_410),
.C(n_392),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_404),
.A2(n_354),
.B(n_378),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_353),
.Y(n_422)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_422),
.Y(n_441)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_436),
.C(n_437),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_427),
.B(n_310),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_387),
.A2(n_371),
.B1(n_374),
.B2(n_359),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_429),
.A2(n_411),
.B1(n_401),
.B2(n_407),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_391),
.A2(n_342),
.B1(n_366),
.B2(n_361),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_359),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_411),
.A2(n_353),
.B1(n_351),
.B2(n_337),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_297),
.C(n_223),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_322),
.C(n_310),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_400),
.C(n_397),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_438),
.A2(n_450),
.B1(n_417),
.B2(n_415),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_406),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_446),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_434),
.B(n_398),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_440),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_395),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_445),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_412),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_388),
.C(n_322),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_455),
.C(n_436),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_451),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_382),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_454),
.C(n_431),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_223),
.C(n_237),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_457),
.A2(n_418),
.B(n_419),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_237),
.Y(n_458)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_438),
.A2(n_416),
.B1(n_428),
.B2(n_414),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_470),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_467),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_435),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

OA22x2_ASAP7_75t_L g464 ( 
.A1(n_442),
.A2(n_416),
.B1(n_420),
.B2(n_421),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_464),
.A2(n_471),
.B1(n_449),
.B2(n_423),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_423),
.Y(n_484)
);

INVx11_ASAP7_75t_L g468 ( 
.A(n_445),
.Y(n_468)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_427),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_SL g472 ( 
.A(n_444),
.B(n_422),
.C(n_423),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_472),
.Y(n_480)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_456),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_474),
.B(n_426),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_468),
.A2(n_441),
.B1(n_433),
.B2(n_449),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_475),
.A2(n_471),
.B1(n_448),
.B2(n_453),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_444),
.C(n_451),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_477),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_455),
.C(n_446),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_466),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_456),
.Y(n_479)
);

AOI21x1_ASAP7_75t_L g491 ( 
.A1(n_479),
.A2(n_458),
.B(n_464),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_486),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_484),
.A2(n_467),
.B1(n_470),
.B2(n_473),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_439),
.C(n_457),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_465),
.B(n_426),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_487),
.B(n_479),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_490),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_475),
.B(n_478),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_494),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_432),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_493),
.B(n_482),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_464),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_462),
.C(n_459),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_498),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_485),
.A2(n_459),
.B(n_454),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_499),
.A2(n_486),
.B1(n_481),
.B2(n_477),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_504),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_501),
.A2(n_497),
.B(n_490),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_488),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_484),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_495),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_507),
.A2(n_502),
.B(n_500),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_508),
.B(n_510),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_503),
.C(n_502),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_424),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_504),
.C(n_499),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_514),
.A2(n_515),
.B1(n_511),
.B2(n_247),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_247),
.B(n_15),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_517),
.A2(n_15),
.B(n_16),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_518),
.B(n_16),
.Y(n_519)
);


endmodule