module fake_jpeg_3127_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_57),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx2_ASAP7_75t_SL g85 ( 
.A(n_78),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_56),
.B1(n_70),
.B2(n_50),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_78),
.B1(n_73),
.B2(n_77),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_56),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_58),
.B(n_61),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_51),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_52),
.B1(n_62),
.B2(n_54),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_71),
.B1(n_68),
.B2(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_28),
.B1(n_42),
.B2(n_41),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_70),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_27),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_71),
.B1(n_68),
.B2(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_67),
.B1(n_58),
.B2(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_67),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_129),
.B1(n_131),
.B2(n_9),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_66),
.B1(n_61),
.B2(n_6),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_61),
.C(n_3),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_102),
.B1(n_114),
.B2(n_9),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_2),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_26),
.Y(n_138)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_138),
.Y(n_163)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_7),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_146),
.Y(n_167)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_117),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_7),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_150),
.B(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_14),
.B1(n_45),
.B2(n_17),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_10),
.B(n_12),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_29),
.B(n_40),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_25),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_13),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_10),
.B(n_12),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_132),
.B(n_13),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_155),
.C(n_145),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_149),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_174),
.A2(n_148),
.B1(n_22),
.B2(n_23),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_152),
.C(n_147),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_155),
.C(n_151),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_14),
.B(n_38),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_180),
.B(n_151),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_37),
.B(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_187),
.B(n_189),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_179),
.B1(n_173),
.B2(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_187),
.B1(n_185),
.B2(n_167),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_168),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_191),
.C(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

NAND2x1_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_197),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_207),
.A2(n_208),
.B(n_187),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_206),
.A2(n_203),
.B1(n_204),
.B2(n_199),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_208),
.B(n_201),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_175),
.A3(n_195),
.B1(n_198),
.B2(n_164),
.C1(n_178),
.C2(n_165),
.Y(n_211)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_163),
.B(n_180),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_16),
.Y(n_213)
);


endmodule