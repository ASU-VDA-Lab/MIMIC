module fake_jpeg_20181_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_1),
.C(n_2),
.Y(n_12)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_3),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_10),
.B1(n_6),
.B2(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_17),
.Y(n_26)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_9),
.B(n_17),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_26),
.B1(n_18),
.B2(n_7),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_12),
.B(n_9),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_16),
.C(n_7),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_19),
.C(n_18),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_30),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_32),
.Y(n_37)
);

AOI221xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B1(n_18),
.B2(n_34),
.C(n_36),
.Y(n_39)
);

NOR4xp25_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_30),
.C(n_3),
.D(n_2),
.Y(n_38)
);


endmodule