module fake_jpeg_4241_n_314 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_37),
.B(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_52),
.Y(n_101)
);

CKINVDCx9p33_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_61),
.Y(n_123)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_33),
.B1(n_17),
.B2(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_69),
.B1(n_83),
.B2(n_18),
.Y(n_105)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_74),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_17),
.B1(n_32),
.B2(n_14),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_26),
.B1(n_19),
.B2(n_20),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_84),
.B1(n_89),
.B2(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_78),
.Y(n_118)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_19),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_81),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_20),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_16),
.B1(n_29),
.B2(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_94),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NAND2xp67_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_22),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_34),
.B(n_18),
.C(n_24),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_99),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_98),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_18),
.B1(n_34),
.B2(n_29),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_18),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_34),
.B1(n_24),
.B2(n_31),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_49),
.A2(n_29),
.B1(n_27),
.B2(n_16),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_16),
.B1(n_27),
.B2(n_18),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_129),
.B(n_145),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_69),
.B1(n_64),
.B2(n_49),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_131),
.B1(n_139),
.B2(n_141),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_66),
.B1(n_58),
.B2(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_135),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_52),
.Y(n_133)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_51),
.B1(n_66),
.B2(n_72),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_83),
.B1(n_61),
.B2(n_65),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_97),
.B(n_55),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_161),
.B(n_128),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_58),
.B1(n_91),
.B2(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_98),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_68),
.B1(n_88),
.B2(n_80),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_148),
.B1(n_150),
.B2(n_156),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_68),
.CI(n_88),
.CON(n_146),
.SN(n_146)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_146),
.B(n_151),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_152),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_31),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_13),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_76),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_74),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_154),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_60),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_96),
.B1(n_90),
.B2(n_87),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_60),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_24),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_141),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_110),
.B1(n_117),
.B2(n_127),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_24),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_0),
.C(n_1),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_104),
.C(n_12),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_167),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_143),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_168),
.A2(n_186),
.B(n_132),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_114),
.Y(n_173)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_195),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_198),
.B(n_199),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_181),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_146),
.Y(n_216)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_187),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_112),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_130),
.A2(n_127),
.B1(n_117),
.B2(n_110),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_131),
.B1(n_144),
.B2(n_129),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_128),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_122),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_104),
.B(n_122),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_153),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_204),
.B(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_175),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_194),
.B1(n_189),
.B2(n_176),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_139),
.B1(n_137),
.B2(n_150),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_223),
.B1(n_171),
.B2(n_174),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_222),
.B1(n_174),
.B2(n_194),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_146),
.B(n_149),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_224),
.B(n_227),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_170),
.B(n_185),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_172),
.A2(n_136),
.B1(n_151),
.B2(n_164),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_163),
.B(n_2),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_177),
.B1(n_170),
.B2(n_171),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_106),
.B(n_2),
.C(n_3),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_198),
.B(n_182),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_212),
.B1(n_225),
.B2(n_216),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_245),
.B(n_202),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_195),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_239),
.C(n_240),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_196),
.B(n_179),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_236),
.B(n_248),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_231),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_226),
.B(n_207),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_241),
.B1(n_250),
.B2(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_189),
.C(n_169),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_167),
.C(n_178),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_178),
.B1(n_167),
.B2(n_100),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_165),
.B(n_2),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_208),
.A2(n_165),
.B1(n_9),
.B2(n_10),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_218),
.B(n_225),
.C(n_206),
.D(n_205),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_223),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_208),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_255),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_219),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_257),
.B(n_259),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_211),
.B1(n_220),
.B2(n_202),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_217),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_264),
.Y(n_274)
);

BUFx12f_ASAP7_75t_SL g263 ( 
.A(n_236),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_209),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_240),
.C(n_239),
.Y(n_272)
);

AOI321xp33_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_233),
.A3(n_245),
.B1(n_249),
.B2(n_225),
.C(n_246),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_236),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_230),
.C(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_258),
.C(n_259),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_232),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_238),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_210),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_288),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_284),
.C(n_286),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_267),
.B(n_258),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_279),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_261),
.C(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_267),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_268),
.A2(n_251),
.B(n_250),
.C(n_248),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_273),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_280),
.B1(n_277),
.B2(n_255),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_253),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_294),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_278),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_299),
.C(n_270),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_209),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_291),
.B(n_290),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_304),
.B(n_305),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_275),
.B1(n_289),
.B2(n_243),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_297),
.B(n_220),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_298),
.C(n_289),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.C(n_8),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_289),
.B(n_250),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_250),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_106),
.Y(n_314)
);


endmodule