module fake_jpeg_24500_n_186 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_15),
.B1(n_28),
.B2(n_18),
.Y(n_51)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_20),
.B1(n_18),
.B2(n_15),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_49),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_17),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_21),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_22),
.B1(n_21),
.B2(n_15),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_29),
.B1(n_28),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_26),
.B1(n_23),
.B2(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_21),
.B1(n_22),
.B2(n_28),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_60),
.B1(n_70),
.B2(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_67),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_65),
.B1(n_73),
.B2(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_34),
.B1(n_31),
.B2(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_38),
.B1(n_16),
.B2(n_25),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_25),
.B1(n_17),
.B2(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_50),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_94),
.B(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_40),
.B1(n_47),
.B2(n_49),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_89),
.B1(n_93),
.B2(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_47),
.B1(n_40),
.B2(n_46),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_40),
.B1(n_46),
.B2(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_56),
.B1(n_16),
.B2(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_102),
.B1(n_88),
.B2(n_92),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_100),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_90),
.B1(n_83),
.B2(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_64),
.B(n_74),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_76),
.B(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_61),
.B1(n_63),
.B2(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_73),
.B1(n_72),
.B2(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_110),
.B1(n_111),
.B2(n_78),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_32),
.C(n_45),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_75),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_45),
.B1(n_71),
.B2(n_16),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_45),
.B1(n_71),
.B2(n_24),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_8),
.B1(n_12),
.B2(n_2),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_82),
.B1(n_76),
.B2(n_2),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_117),
.B1(n_75),
.B2(n_4),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_82),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_75),
.C(n_1),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_97),
.B1(n_100),
.B2(n_106),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_99),
.B1(n_103),
.B2(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_139),
.B1(n_142),
.B2(n_6),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_105),
.B(n_98),
.C(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_6),
.Y(n_151)
);

OAI322xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_101),
.A3(n_109),
.B1(n_104),
.B2(n_102),
.C1(n_111),
.C2(n_75),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_135),
.C(n_138),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_137),
.Y(n_146)
);

NAND2x1_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_0),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_113),
.C(n_7),
.Y(n_149)
);

AO22x1_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_128),
.B1(n_125),
.B2(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_122),
.B1(n_117),
.B2(n_123),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_150),
.B(n_151),
.Y(n_161)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.C(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_142),
.C(n_135),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_153),
.C(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_156),
.C(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_147),
.C(n_145),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_142),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_166),
.C(n_169),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_152),
.B1(n_131),
.B2(n_144),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_168),
.B1(n_160),
.B2(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_148),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_161),
.A2(n_140),
.B1(n_130),
.B2(n_148),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_8),
.B(n_9),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_7),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_7),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_170),
.B(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_178),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_10),
.B(n_11),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_177),
.B(n_175),
.C(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_10),
.B(n_11),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_12),
.B(n_13),
.Y(n_186)
);


endmodule