module real_aes_17824_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AND2x4_ASAP7_75t_L g822 ( .A(n_0), .B(n_823), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_1), .A2(n_4), .B1(n_251), .B2(n_252), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_2), .A2(n_42), .B1(n_152), .B2(n_200), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_3), .A2(n_24), .B1(n_200), .B2(n_234), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_5), .A2(n_16), .B1(n_502), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_6), .A2(n_60), .B1(n_137), .B2(n_138), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_7), .A2(n_17), .B1(n_152), .B2(n_153), .Y(n_151) );
INVx1_ASAP7_75t_L g823 ( .A(n_8), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_9), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_10), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_11), .A2(n_18), .B1(n_503), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_12), .A2(n_113), .B1(n_778), .B2(n_779), .Y(n_112) );
INVx1_ASAP7_75t_L g778 ( .A(n_12), .Y(n_778) );
OR2x2_ASAP7_75t_L g111 ( .A(n_13), .B(n_37), .Y(n_111) );
BUFx2_ASAP7_75t_L g817 ( .A(n_13), .Y(n_817) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_14), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_15), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_19), .A2(n_96), .B1(n_252), .B2(n_502), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_20), .A2(n_38), .B1(n_130), .B2(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_21), .B(n_128), .Y(n_563) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_22), .A2(n_58), .B(n_143), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_23), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_25), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_26), .B(n_125), .Y(n_192) );
INVx4_ASAP7_75t_R g176 ( .A(n_27), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_28), .A2(n_46), .B1(n_156), .B2(n_249), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_29), .A2(n_54), .B1(n_156), .B2(n_502), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_30), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_31), .B(n_527), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_32), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_33), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g256 ( .A(n_34), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_SL g231 ( .A1(n_35), .A2(n_124), .B(n_152), .C(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_36), .A2(n_55), .B1(n_152), .B2(n_156), .Y(n_240) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_37), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_39), .A2(n_84), .B1(n_152), .B2(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_40), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_40), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_41), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_43), .A2(n_45), .B1(n_152), .B2(n_153), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_44), .A2(n_59), .B1(n_502), .B2(n_519), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_47), .Y(n_825) );
INVx1_ASAP7_75t_L g196 ( .A(n_48), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_49), .B(n_152), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_50), .Y(n_210) );
INVx2_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
BUFx3_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g788 ( .A(n_52), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_53), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_56), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_57), .A2(n_85), .B1(n_152), .B2(n_156), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_61), .A2(n_73), .B1(n_249), .B2(n_519), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_62), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_63), .A2(n_76), .B1(n_152), .B2(n_153), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_64), .A2(n_95), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g143 ( .A(n_65), .Y(n_143) );
AND2x4_ASAP7_75t_L g146 ( .A(n_66), .B(n_147), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_67), .A2(n_87), .B1(n_156), .B2(n_249), .Y(n_248) );
AO22x1_ASAP7_75t_L g126 ( .A1(n_68), .A2(n_74), .B1(n_127), .B2(n_130), .Y(n_126) );
INVx1_ASAP7_75t_L g147 ( .A(n_69), .Y(n_147) );
AND2x2_ASAP7_75t_L g235 ( .A(n_70), .B(n_188), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_71), .B(n_137), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_72), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_75), .B(n_200), .Y(n_211) );
INVx2_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_78), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_79), .B(n_188), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_80), .A2(n_94), .B1(n_137), .B2(n_156), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_81), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_82), .B(n_141), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_83), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_86), .B(n_188), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_88), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_89), .B(n_188), .Y(n_207) );
INVx1_ASAP7_75t_L g474 ( .A(n_90), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_90), .B(n_787), .Y(n_786) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_91), .B(n_128), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_92), .A2(n_137), .B(n_158), .C(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g181 ( .A(n_93), .B(n_182), .Y(n_181) );
NAND2xp33_ASAP7_75t_L g215 ( .A(n_97), .B(n_177), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_98), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_813), .B(n_824), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_789), .Y(n_100) );
OAI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_112), .B(n_780), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x6_ASAP7_75t_SL g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_L g792 ( .A(n_106), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_106), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x1_ASAP7_75t_L g812 ( .A(n_109), .B(n_111), .Y(n_812) );
NOR3x1_ASAP7_75t_L g820 ( .A(n_109), .B(n_804), .C(n_821), .Y(n_820) );
AND2x6_ASAP7_75t_SL g785 ( .A(n_110), .B(n_786), .Y(n_785) );
AND3x2_ASAP7_75t_L g802 ( .A(n_110), .B(n_803), .C(n_804), .Y(n_802) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g779 ( .A(n_113), .Y(n_779) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_471), .B1(n_475), .B2(n_777), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_381), .Y(n_115) );
NOR3xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_310), .C(n_352), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_284), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_183), .B1(n_259), .B2(n_270), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_164), .Y(n_120) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_121), .A2(n_304), .B(n_306), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_121), .A2(n_377), .B(n_378), .Y(n_376) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_148), .Y(n_121) );
INVx2_ASAP7_75t_L g296 ( .A(n_122), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_122), .B(n_149), .Y(n_326) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B(n_132), .C(n_144), .Y(n_123) );
INVx6_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_124), .A2(n_215), .B(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_124), .B(n_126), .Y(n_268) );
O2A1O1Ixp5_ASAP7_75t_L g561 ( .A1(n_124), .A2(n_153), .B(n_562), .C(n_563), .Y(n_561) );
BUFx8_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g135 ( .A(n_125), .Y(n_135) );
INVx1_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
INVx1_ASAP7_75t_L g195 ( .A(n_125), .Y(n_195) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g502 ( .A(n_128), .Y(n_502) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_129), .Y(n_131) );
INVx1_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_129), .Y(n_139) );
INVx3_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_129), .Y(n_200) );
INVx1_ASAP7_75t_L g228 ( .A(n_129), .Y(n_228) );
INVx2_ASAP7_75t_L g234 ( .A(n_129), .Y(n_234) );
OAI21xp33_ASAP7_75t_SL g191 ( .A1(n_130), .A2(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g267 ( .A(n_132), .Y(n_267) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_136), .B(n_140), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_133), .A2(n_198), .B(n_199), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_133), .A2(n_154), .B1(n_239), .B2(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g485 ( .A(n_134), .Y(n_485) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
INVx1_ASAP7_75t_L g547 ( .A(n_138), .Y(n_547) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_139), .B(n_173), .Y(n_172) );
OAI21xp33_ASAP7_75t_L g144 ( .A1(n_140), .A2(n_141), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
INVx2_ASAP7_75t_L g163 ( .A(n_141), .Y(n_163) );
INVx2_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g269 ( .A(n_144), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_145), .A2(n_224), .B(n_231), .Y(n_223) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx10_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
BUFx10_ASAP7_75t_L g202 ( .A(n_146), .Y(n_202) );
INVx1_ASAP7_75t_L g254 ( .A(n_146), .Y(n_254) );
AND2x2_ASAP7_75t_L g366 ( .A(n_148), .B(n_205), .Y(n_366) );
INVx1_ASAP7_75t_L g399 ( .A(n_148), .Y(n_399) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g261 ( .A(n_149), .B(n_206), .Y(n_261) );
AND2x2_ASAP7_75t_L g292 ( .A(n_149), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g301 ( .A(n_149), .Y(n_301) );
OR2x2_ASAP7_75t_L g320 ( .A(n_149), .B(n_166), .Y(n_320) );
AND2x2_ASAP7_75t_L g335 ( .A(n_149), .B(n_166), .Y(n_335) );
AO31x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_159), .A3(n_160), .B(n_161), .Y(n_149) );
OAI22x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B1(n_155), .B2(n_157), .Y(n_150) );
INVx4_ASAP7_75t_L g153 ( .A(n_152), .Y(n_153) );
INVx1_ASAP7_75t_L g503 ( .A(n_152), .Y(n_503) );
INVx1_ASAP7_75t_L g519 ( .A(n_152), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_153), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_154), .A2(n_157), .B1(n_248), .B2(n_250), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_154), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_154), .A2(n_157), .B1(n_493), .B2(n_495), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_154), .A2(n_501), .B1(n_504), .B2(n_505), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_154), .A2(n_485), .B1(n_517), .B2(n_518), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_154), .A2(n_485), .B1(n_526), .B2(n_528), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_154), .A2(n_485), .B1(n_536), .B2(n_537), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_154), .A2(n_505), .B1(n_546), .B2(n_548), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_154), .A2(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_156), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g251 ( .A(n_156), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_157), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_SL g505 ( .A(n_158), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_159), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_159), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g180 ( .A(n_160), .Y(n_180) );
AO31x2_ASAP7_75t_L g482 ( .A1(n_160), .A2(n_241), .A3(n_483), .B(n_487), .Y(n_482) );
AO31x2_ASAP7_75t_L g524 ( .A1(n_160), .A2(n_491), .A3(n_525), .B(n_530), .Y(n_524) );
AO31x2_ASAP7_75t_L g544 ( .A1(n_160), .A2(n_222), .A3(n_545), .B(n_549), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx2_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
BUFx2_ASAP7_75t_L g222 ( .A(n_163), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_163), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_163), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_165), .B(n_334), .Y(n_377) );
OR2x2_ASAP7_75t_L g465 ( .A(n_165), .B(n_326), .Y(n_465) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g293 ( .A(n_166), .Y(n_293) );
AND2x2_ASAP7_75t_L g302 ( .A(n_166), .B(n_265), .Y(n_302) );
AND2x2_ASAP7_75t_L g305 ( .A(n_166), .B(n_206), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_166), .B(n_205), .Y(n_324) );
AND2x4_ASAP7_75t_L g343 ( .A(n_166), .B(n_266), .Y(n_343) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_181), .Y(n_166) );
AO31x2_ASAP7_75t_L g515 ( .A1(n_167), .A2(n_506), .A3(n_516), .B(n_520), .Y(n_515) );
AO31x2_ASAP7_75t_L g534 ( .A1(n_167), .A2(n_253), .A3(n_535), .B(n_538), .Y(n_534) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_169), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_SL g549 ( .A(n_169), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_180), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_175) );
INVx2_ASAP7_75t_L g249 ( .A(n_177), .Y(n_249) );
INVx1_ASAP7_75t_L g527 ( .A(n_177), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_178), .Y(n_529) );
INVx1_ASAP7_75t_L g506 ( .A(n_180), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_203), .B(n_244), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_184), .B(n_338), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_186), .B(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g274 ( .A(n_186), .Y(n_274) );
OR2x2_ASAP7_75t_L g282 ( .A(n_186), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_186), .B(n_275), .Y(n_307) );
AND2x2_ASAP7_75t_L g332 ( .A(n_186), .B(n_246), .Y(n_332) );
AND2x2_ASAP7_75t_L g350 ( .A(n_186), .B(n_280), .Y(n_350) );
INVx1_ASAP7_75t_L g389 ( .A(n_186), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_186), .B(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_SL g410 ( .A(n_186), .B(n_331), .Y(n_410) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_190), .Y(n_186) );
NOR2x1_ASAP7_75t_L g217 ( .A(n_188), .B(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g241 ( .A(n_188), .Y(n_241) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g201 ( .A(n_189), .B(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_189), .B(n_488), .Y(n_487) );
BUFx3_ASAP7_75t_L g491 ( .A(n_189), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_189), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_189), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g559 ( .A(n_189), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_197), .B(n_201), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_195), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_200), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g218 ( .A(n_202), .Y(n_218) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_202), .A2(n_238), .A3(n_241), .B(n_242), .Y(n_237) );
OAI32xp33_ASAP7_75t_L g294 ( .A1(n_203), .A2(n_286), .A3(n_295), .B1(n_297), .B2(n_299), .Y(n_294) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_219), .Y(n_203) );
INVx1_ASAP7_75t_L g334 ( .A(n_204), .Y(n_334) );
AND2x2_ASAP7_75t_L g342 ( .A(n_204), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g341 ( .A(n_205), .B(n_265), .Y(n_341) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx3_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
AND2x2_ASAP7_75t_L g300 ( .A(n_206), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g406 ( .A(n_206), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_214), .B(n_217), .Y(n_208) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
OR2x2_ASAP7_75t_L g286 ( .A(n_219), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g408 ( .A(n_219), .Y(n_408) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_236), .Y(n_219) );
AND2x2_ASAP7_75t_L g309 ( .A(n_220), .B(n_237), .Y(n_309) );
INVx2_ASAP7_75t_L g331 ( .A(n_220), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_220), .B(n_246), .Y(n_351) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
AOI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_235), .Y(n_221) );
AO31x2_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_247), .A3(n_253), .B(n_255), .Y(n_246) );
AO31x2_ASAP7_75t_L g499 ( .A1(n_222), .A2(n_500), .A3(n_506), .B(n_507), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B(n_230), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_SL g494 ( .A(n_234), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_236), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g340 ( .A(n_236), .Y(n_340) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
BUFx2_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
OR2x2_ASAP7_75t_L g346 ( .A(n_237), .B(n_246), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_237), .B(n_246), .Y(n_379) );
INVx2_ASAP7_75t_L g327 ( .A(n_244), .Y(n_327) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_257), .Y(n_244) );
OR2x2_ASAP7_75t_L g314 ( .A(n_245), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g392 ( .A(n_245), .Y(n_392) );
INVx1_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
INVx1_ASAP7_75t_L g283 ( .A(n_246), .Y(n_283) );
INVx1_ASAP7_75t_L g298 ( .A(n_246), .Y(n_298) );
AO31x2_ASAP7_75t_L g490 ( .A1(n_253), .A2(n_491), .A3(n_492), .B(n_496), .Y(n_490) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_SL g567 ( .A(n_254), .Y(n_567) );
OR2x2_ASAP7_75t_L g402 ( .A(n_257), .B(n_379), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_258), .B(n_274), .Y(n_315) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
OR2x2_ASAP7_75t_L g416 ( .A(n_258), .B(n_340), .Y(n_416) );
INVxp67_ASAP7_75t_L g440 ( .A(n_258), .Y(n_440) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NAND2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_261), .B(n_302), .Y(n_369) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g318 ( .A(n_263), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g431 ( .A(n_264), .Y(n_431) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g460 ( .A(n_265), .B(n_293), .Y(n_460) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g386 ( .A(n_266), .B(n_293), .Y(n_386) );
AOI21x1_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_277), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_273), .B(n_309), .Y(n_423) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g287 ( .A(n_274), .Y(n_287) );
AND2x2_ASAP7_75t_L g337 ( .A(n_274), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_274), .B(n_331), .Y(n_380) );
OR2x2_ASAP7_75t_L g452 ( .A(n_274), .B(n_339), .Y(n_452) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g372 ( .A(n_278), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g363 ( .A(n_279), .Y(n_363) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g353 ( .A(n_282), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_282), .Y(n_364) );
OR2x2_ASAP7_75t_L g415 ( .A(n_282), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g470 ( .A(n_282), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B(n_294), .C(n_303), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g359 ( .A(n_287), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_287), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g432 ( .A(n_287), .B(n_309), .Y(n_432) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_290), .B(n_335), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_290), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g442 ( .A(n_290), .B(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g385 ( .A(n_291), .Y(n_385) );
AND2x2_ASAP7_75t_L g413 ( .A(n_292), .B(n_341), .Y(n_413) );
INVx2_ASAP7_75t_L g436 ( .A(n_292), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_292), .B(n_334), .Y(n_468) );
AND2x4_ASAP7_75t_SL g422 ( .A(n_295), .B(n_300), .Y(n_422) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g375 ( .A(n_296), .B(n_301), .Y(n_375) );
OR2x2_ASAP7_75t_L g427 ( .A(n_296), .B(n_320), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_297), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_297), .B(n_309), .Y(n_463) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g411 ( .A(n_298), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g394 ( .A(n_300), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_300), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g444 ( .A(n_301), .Y(n_444) );
BUFx2_ASAP7_75t_L g312 ( .A(n_302), .Y(n_312) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g430 ( .A(n_305), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g354 ( .A(n_309), .Y(n_354) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_309), .Y(n_371) );
NAND3xp33_ASAP7_75t_SL g310 ( .A(n_311), .B(n_321), .C(n_336), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_313), .B1(n_316), .B2(n_318), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_318), .A2(n_344), .B1(n_425), .B2(n_428), .C1(n_430), .C2(n_432), .Y(n_424) );
AND2x2_ASAP7_75t_L g456 ( .A(n_319), .B(n_405), .Y(n_456) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g404 ( .A(n_320), .B(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_327), .B1(n_328), .B2(n_333), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_SL g400 ( .A(n_324), .Y(n_400) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AND2x2_ASAP7_75t_L g387 ( .A(n_329), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g345 ( .A(n_330), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g339 ( .A(n_331), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g454 ( .A(n_332), .Y(n_454) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_335), .B(n_431), .Y(n_450) );
INVx1_ASAP7_75t_L g467 ( .A(n_335), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B1(n_342), .B2(n_344), .C1(n_347), .C2(n_348), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_343), .Y(n_347) );
AND2x2_ASAP7_75t_L g365 ( .A(n_343), .B(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g396 ( .A(n_343), .Y(n_396) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g360 ( .A(n_346), .Y(n_360) );
OR2x2_ASAP7_75t_L g429 ( .A(n_346), .B(n_410), .Y(n_429) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_358), .C(n_367), .Y(n_352) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_365), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_359), .A2(n_397), .B1(n_446), .B2(n_449), .C(n_451), .Y(n_445) );
AND2x4_ASAP7_75t_L g388 ( .A(n_360), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g419 ( .A(n_366), .Y(n_419) );
AOI211x1_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B(n_372), .C(n_376), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g437 ( .A(n_375), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_378), .B(n_426), .C(n_427), .Y(n_425) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g461 ( .A(n_379), .Y(n_461) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_433), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .C(n_412), .D(n_424), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g443 ( .A(n_386), .B(n_444), .Y(n_443) );
AOI221x1_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_413), .B1(n_414), .B2(n_417), .C(n_420), .Y(n_412) );
AND2x2_ASAP7_75t_L g438 ( .A(n_388), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_397), .B2(n_401), .C(n_403), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_395), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_400), .A2(n_404), .B1(n_407), .B2(n_409), .Y(n_403) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_404), .A2(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g426 ( .A(n_406), .Y(n_426) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g447 ( .A(n_416), .Y(n_447) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_429), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_445), .C(n_457), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B1(n_441), .B2(n_442), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g453 ( .A(n_440), .B(n_454), .Y(n_453) );
NAND2x1_ASAP7_75t_L g469 ( .A(n_440), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_455), .Y(n_451) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B1(n_462), .B2(n_464), .C(n_466), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g777 ( .A(n_471), .Y(n_777) );
BUFx12f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g811 ( .A(n_473), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g804 ( .A(n_474), .Y(n_804) );
INVx2_ASAP7_75t_L g796 ( .A(n_475), .Y(n_796) );
NOR2x1p5_ASAP7_75t_L g475 ( .A(n_476), .B(n_687), .Y(n_475) );
NAND4xp75_ASAP7_75t_L g476 ( .A(n_477), .B(n_632), .C(n_652), .D(n_668), .Y(n_476) );
NOR2x1p5_ASAP7_75t_SL g477 ( .A(n_478), .B(n_602), .Y(n_477) );
NAND4xp75_ASAP7_75t_L g478 ( .A(n_479), .B(n_540), .C(n_579), .D(n_588), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_509), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
AND2x4_ASAP7_75t_L g712 ( .A(n_481), .B(n_639), .Y(n_712) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_482), .Y(n_555) );
INVx2_ASAP7_75t_L g573 ( .A(n_482), .Y(n_573) );
AND2x2_ASAP7_75t_L g596 ( .A(n_482), .B(n_558), .Y(n_596) );
OR2x2_ASAP7_75t_L g651 ( .A(n_482), .B(n_490), .Y(n_651) );
AND2x2_ASAP7_75t_L g569 ( .A(n_489), .B(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g719 ( .A(n_489), .B(n_596), .Y(n_719) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
OR2x2_ASAP7_75t_L g556 ( .A(n_490), .B(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
AND2x2_ASAP7_75t_L g593 ( .A(n_490), .B(n_499), .Y(n_593) );
INVx1_ASAP7_75t_L g611 ( .A(n_490), .Y(n_611) );
INVx2_ASAP7_75t_L g640 ( .A(n_490), .Y(n_640) );
INVx3_ASAP7_75t_L g616 ( .A(n_498), .Y(n_616) );
INVx2_ASAP7_75t_L g621 ( .A(n_498), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_498), .B(n_572), .Y(n_626) );
AND2x2_ASAP7_75t_L g649 ( .A(n_498), .B(n_628), .Y(n_649) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_498), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_498), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g638 ( .A(n_499), .Y(n_638) );
AND2x2_ASAP7_75t_L g686 ( .A(n_499), .B(n_640), .Y(n_686) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_511), .B(n_630), .Y(n_677) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_512), .B(n_630), .Y(n_674) );
INVx1_ASAP7_75t_L g775 ( .A(n_512), .Y(n_775) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g725 ( .A(n_513), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g578 ( .A(n_514), .Y(n_578) );
OR2x2_ASAP7_75t_L g659 ( .A(n_514), .B(n_533), .Y(n_659) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g601 ( .A(n_515), .Y(n_601) );
AND2x4_ASAP7_75t_L g607 ( .A(n_515), .B(n_608), .Y(n_607) );
AOI32xp33_ASAP7_75t_L g745 ( .A1(n_522), .A2(n_648), .A3(n_746), .B1(n_748), .B2(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g694 ( .A(n_523), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_532), .Y(n_523) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_524), .Y(n_542) );
OR2x2_ASAP7_75t_L g576 ( .A(n_524), .B(n_534), .Y(n_576) );
INVx1_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
AND2x2_ASAP7_75t_L g600 ( .A(n_524), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g606 ( .A(n_524), .Y(n_606) );
INVx2_ASAP7_75t_L g631 ( .A(n_524), .Y(n_631) );
AND2x2_ASAP7_75t_L g750 ( .A(n_524), .B(n_544), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_532), .B(n_583), .Y(n_670) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g543 ( .A(n_534), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g599 ( .A(n_534), .Y(n_599) );
INVx2_ASAP7_75t_L g608 ( .A(n_534), .Y(n_608) );
AND2x4_ASAP7_75t_L g630 ( .A(n_534), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_534), .Y(n_722) );
AOI22x1_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_551), .B1(n_569), .B2(n_574), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_543), .B(n_700), .C(n_701), .D(n_702), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_543), .B(n_600), .Y(n_730) );
INVx4_ASAP7_75t_SL g583 ( .A(n_544), .Y(n_583) );
BUFx2_ASAP7_75t_L g646 ( .A(n_544), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_544), .B(n_591), .Y(n_709) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g671 ( .A(n_553), .B(n_620), .Y(n_671) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g594 ( .A(n_557), .B(n_572), .Y(n_594) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_558), .B(n_573), .Y(n_618) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_568), .Y(n_558) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_559), .A2(n_560), .B(n_568), .Y(n_613) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B(n_567), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_570), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g636 ( .A(n_570), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g675 ( .A(n_571), .B(n_593), .Y(n_675) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g718 ( .A(n_573), .B(n_628), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_574), .A2(n_691), .B1(n_693), .B2(n_696), .C(n_698), .Y(n_690) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g584 ( .A(n_576), .Y(n_584) );
OR2x2_ASAP7_75t_L g684 ( .A(n_576), .B(n_623), .Y(n_684) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_580), .A2(n_706), .B1(n_710), .B2(n_713), .Y(n_705) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
AND2x4_ASAP7_75t_L g629 ( .A(n_581), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g741 ( .A(n_581), .B(n_659), .Y(n_741) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g589 ( .A(n_583), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g605 ( .A(n_583), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g664 ( .A(n_583), .B(n_601), .Y(n_664) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_583), .Y(n_681) );
INVx1_ASAP7_75t_L g695 ( .A(n_583), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_583), .B(n_608), .Y(n_738) );
AND2x4_ASAP7_75t_L g645 ( .A(n_584), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g643 ( .A(n_586), .Y(n_643) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_587), .B(n_628), .Y(n_627) );
NAND2x1_ASAP7_75t_L g747 ( .A(n_587), .B(n_649), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B1(n_595), .B2(n_597), .Y(n_588) );
AND2x2_ASAP7_75t_L g614 ( .A(n_589), .B(n_607), .Y(n_614) );
INVx1_ASAP7_75t_L g655 ( .A(n_589), .Y(n_655) );
AND2x2_ASAP7_75t_L g762 ( .A(n_589), .B(n_623), .Y(n_762) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g595 ( .A(n_593), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g735 ( .A(n_593), .Y(n_735) );
AND2x2_ASAP7_75t_L g752 ( .A(n_593), .B(n_612), .Y(n_752) );
AND2x2_ASAP7_75t_L g768 ( .A(n_593), .B(n_718), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_594), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g691 ( .A(n_594), .B(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_594), .A2(n_684), .B1(n_699), .B2(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g654 ( .A(n_596), .Y(n_654) );
AND2x2_ASAP7_75t_L g685 ( .A(n_596), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_596), .B(n_692), .Y(n_714) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g720 ( .A(n_600), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_600), .A2(n_624), .B1(n_729), .B2(n_731), .Y(n_728) );
INVx3_ASAP7_75t_L g623 ( .A(n_601), .Y(n_623) );
AND2x2_ASAP7_75t_L g755 ( .A(n_601), .B(n_608), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_619), .Y(n_602) );
AOI32xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_609), .A3(n_612), .B1(n_614), .B2(n_615), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_606), .Y(n_701) );
INVx1_ASAP7_75t_L g726 ( .A(n_606), .Y(n_726) );
INVx3_ASAP7_75t_L g682 ( .A(n_607), .Y(n_682) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_610), .A2(n_758), .B1(n_759), .B2(n_760), .C(n_761), .Y(n_757) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g734 ( .A(n_612), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g770 ( .A(n_612), .B(n_731), .Y(n_770) );
BUFx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g628 ( .A(n_613), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_615), .B(n_643), .Y(n_642) );
AO22x1_ASAP7_75t_L g672 ( .A1(n_615), .A2(n_673), .B1(n_675), .B2(n_676), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g776 ( .A(n_615), .B(n_643), .Y(n_776) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g692 ( .A(n_616), .Y(n_692) );
INVx1_ASAP7_75t_L g702 ( .A(n_616), .Y(n_702) );
AND2x2_ASAP7_75t_L g622 ( .A(n_617), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_618), .Y(n_704) );
INVx1_ASAP7_75t_L g744 ( .A(n_618), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B(n_624), .C(n_629), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2x1p5_ASAP7_75t_L g731 ( .A(n_621), .B(n_651), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_622), .B(n_681), .Y(n_758) );
AOI31xp33_ASAP7_75t_L g641 ( .A1(n_623), .A2(n_642), .A3(n_644), .B(n_647), .Y(n_641) );
INVx4_ASAP7_75t_L g700 ( .A(n_623), .Y(n_700) );
OR2x2_ASAP7_75t_L g737 ( .A(n_623), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x4_ASAP7_75t_L g639 ( .A(n_628), .B(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_630), .Y(n_635) );
AND2x2_ASAP7_75t_L g666 ( .A(n_630), .B(n_664), .Y(n_666) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_633), .B(n_641), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g759 ( .A(n_636), .Y(n_759) );
INVx1_ASAP7_75t_L g667 ( .A(n_637), .Y(n_667) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g697 ( .A(n_638), .Y(n_697) );
AND2x2_ASAP7_75t_L g696 ( .A(n_639), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI322xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .A3(n_656), .B1(n_660), .B2(n_663), .C1(n_665), .C2(n_667), .Y(n_653) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI211x1_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_678), .Y(n_668) );
INVx1_ASAP7_75t_L g773 ( .A(n_669), .Y(n_773) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g727 ( .A(n_671), .Y(n_727) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OA21x2_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_683), .B(n_685), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx2_ASAP7_75t_L g748 ( .A(n_682), .Y(n_748) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp33_ASAP7_75t_L g743 ( .A(n_686), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_756), .Y(n_687) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_723), .C(n_739), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_705), .C(n_715), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_692), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_696), .A2(n_752), .B(n_753), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_700), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_700), .B(n_750), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_701), .B(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_702), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g761 ( .A1(n_712), .A2(n_762), .B(n_763), .Y(n_761) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .B(n_728), .C(n_732), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_734), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_738), .Y(n_760) );
OAI211xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_742), .B(n_745), .C(n_751), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_750), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g771 ( .A(n_750), .Y(n_771) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g767 ( .A(n_755), .Y(n_767) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_765), .C(n_772), .Y(n_756) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI21xp33_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_769), .B(n_771), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI21xp33_ASAP7_75t_R g772 ( .A1(n_773), .A2(n_774), .B(n_776), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_780), .A2(n_794), .B(n_798), .Y(n_793) );
INVxp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
BUFx12f_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx4_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_788), .Y(n_803) );
AO21x1_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_793), .B(n_805), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx4_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx10_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
BUFx3_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
BUFx12f_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx4f_ASAP7_75t_L g826 ( .A(n_815), .Y(n_826) );
AND2x6_ASAP7_75t_L g815 ( .A(n_816), .B(n_820), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVxp33_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
NOR2xp33_ASAP7_75t_SL g824 ( .A(n_825), .B(n_826), .Y(n_824) );
endmodule