module real_aes_8563_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_22;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
AOI21xp33_ASAP7_75t_SL g15 ( .A1(n_0), .A2(n_2), .B(n_4), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_0), .B(n_22), .Y(n_21) );
CKINVDCx14_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_1), .B(n_10), .Y(n_14) );
NAND3xp33_ASAP7_75t_SL g23 ( .A(n_2), .B(n_5), .C(n_13), .Y(n_23) );
O2A1O1Ixp33_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_7), .B(n_15), .C(n_16), .Y(n_6) );
INVx1_ASAP7_75t_L g22 ( .A(n_3), .Y(n_22) );
INVx1_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_4), .A2(n_12), .B(n_13), .Y(n_11) );
INVx2_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_10), .B(n_11), .Y(n_8) );
INVx1_ASAP7_75t_SL g13 ( .A(n_14), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
CKINVDCx9p33_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
CKINVDCx9p33_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_21), .B(n_23), .Y(n_20) );
endmodule