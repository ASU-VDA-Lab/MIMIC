module fake_jpeg_6090_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_18),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_28),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_19),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_16),
.B(n_25),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_16),
.B1(n_14),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_15),
.B1(n_20),
.B2(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_15),
.B1(n_20),
.B2(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_53),
.B1(n_45),
.B2(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_11),
.B1(n_23),
.B2(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_3),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_47),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_4),
.B(n_6),
.Y(n_59)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_53),
.CI(n_51),
.CON(n_65),
.SN(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_64),
.B1(n_58),
.B2(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_9),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_61),
.C(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_6),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_73),
.C(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_7),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_73),
.C(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_75),
.Y(n_77)
);


endmodule