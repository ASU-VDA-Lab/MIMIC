module fake_jpeg_23588_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_2),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_11),
.B1(n_8),
.B2(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx24_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_15),
.B1(n_16),
.B2(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

XNOR2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_30),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.C(n_43),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_42),
.C(n_30),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_46),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_27),
.Y(n_54)
);


endmodule