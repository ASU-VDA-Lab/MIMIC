module fake_netlist_6_553_n_2471 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2471);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2471;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1371;
wire n_1285;
wire n_383;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2468;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2373;
wire n_2050;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_56),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_140),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_122),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_142),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_53),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_9),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_111),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_173),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_169),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_144),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_167),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_171),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_71),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_115),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_46),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_73),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_126),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_132),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_212),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_8),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_42),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_25),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_2),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_67),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_79),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_131),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_73),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_211),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_218),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_99),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_41),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_135),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_164),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_107),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_124),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_198),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_25),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_83),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_159),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_127),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_147),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_91),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_210),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_48),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_55),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_123),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_109),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_70),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_102),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_32),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_118),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_23),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_35),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_94),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_69),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_104),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_53),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_121),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_214),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_41),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_64),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_28),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_80),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_182),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_108),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_192),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_174),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_89),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_186),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_27),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_69),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_155),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_65),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_152),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_38),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_13),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_23),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_117),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_230),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_102),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_45),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_67),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_68),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_175),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_19),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_47),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_137),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_35),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_228),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_224),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_219),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_181),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_168),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_49),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_184),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_11),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_65),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_180),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_208),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_134),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_66),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_217),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_21),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_148),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_191),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_60),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_81),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_34),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_103),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_6),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_48),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_216),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_97),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_96),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_89),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_85),
.Y(n_367)
);

INVxp33_ASAP7_75t_R g368 ( 
.A(n_103),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_98),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_170),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_177),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_225),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_59),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_204),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_68),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_10),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_178),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_20),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_86),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_54),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_24),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_72),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_18),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_133),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_30),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_18),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_113),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_119),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_213),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_166),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_55),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_176),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_146),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_220),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_149),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_187),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_100),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_3),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_74),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_172),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_90),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_207),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_44),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_70),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_163),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_24),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_17),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_153),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_203),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_66),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_202),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_75),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_99),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_141),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_9),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_165),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_190),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_11),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_51),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_120),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_72),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_82),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_19),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_114),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_74),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_93),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_0),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_16),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_17),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_194),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_13),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_1),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_199),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_79),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_50),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_38),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_85),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_75),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_22),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_52),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_110),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_221),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_128),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_112),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_40),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_57),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_139),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_54),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_154),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_91),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_47),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_197),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_22),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_6),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_94),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_33),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_130),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_238),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_257),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_257),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_238),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_415),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_316),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_234),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_401),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_259),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_235),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_236),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_237),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_243),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_241),
.B(n_0),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_244),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_356),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_294),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_236),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_249),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_440),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_440),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_249),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_440),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_245),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_315),
.B(n_1),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_338),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_441),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_441),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_338),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_424),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_248),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_R g496 ( 
.A(n_424),
.B(n_106),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_251),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_233),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_294),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_265),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_265),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_241),
.B(n_2),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_253),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_255),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_265),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_392),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_309),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_258),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_392),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_309),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_309),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_261),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_262),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_263),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_270),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_241),
.B(n_3),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_354),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_272),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_273),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_276),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_280),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_354),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_294),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_354),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_391),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_282),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_391),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_344),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_412),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_285),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_344),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_287),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_401),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_288),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_293),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_298),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_242),
.B(n_4),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_306),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_307),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g546 ( 
.A(n_277),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_426),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_313),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_321),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_323),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_L g552 ( 
.A(n_315),
.B(n_4),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_328),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_344),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_283),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_445),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_239),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_R g558 ( 
.A(n_315),
.B(n_5),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_330),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_315),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_335),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_341),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_401),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_316),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_242),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_342),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_236),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_247),
.B(n_5),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_286),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_343),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_267),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_346),
.Y(n_573)
);

INVxp33_ASAP7_75t_SL g574 ( 
.A(n_240),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_350),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_267),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_274),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_274),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_247),
.B(n_7),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_292),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_247),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_487),
.B(n_304),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_458),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_467),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_470),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_459),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_460),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_473),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_469),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_464),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

OA21x2_ASAP7_75t_L g594 ( 
.A1(n_479),
.A2(n_340),
.B(n_304),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_561),
.B(n_379),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_570),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_570),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_474),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_479),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_476),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_507),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_471),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_557),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_481),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_487),
.B(n_277),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_481),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_581),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_482),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_482),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_483),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_510),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_499),
.B(n_524),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_462),
.A2(n_297),
.B1(n_365),
.B2(n_301),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_483),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_535),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_535),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_459),
.B(n_286),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_486),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_494),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_552),
.B(n_304),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_581),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_485),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_497),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_468),
.B(n_340),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_493),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_504),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_472),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_564),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_505),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_R g636 ( 
.A(n_509),
.B(n_355),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_552),
.B(n_340),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_493),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_514),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_515),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_564),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_519),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_500),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_500),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_472),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_477),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_478),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_529),
.B(n_379),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_468),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_520),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_566),
.B(n_351),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_521),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_472),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_472),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_475),
.B(n_252),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_478),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_461),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_522),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_527),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_572),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_533),
.B(n_379),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_463),
.B(n_352),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_534),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_478),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_461),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_568),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_536),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_568),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_503),
.B(n_411),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_537),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_568),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_540),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_544),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_480),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_670),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_671),
.B(n_463),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_670),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_598),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_583),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_583),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_584),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_598),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_584),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_671),
.B(n_649),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_599),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_589),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_582),
.B(n_554),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_589),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_651),
.B(n_489),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_588),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_653),
.A2(n_582),
.B1(n_637),
.B2(n_624),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_589),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_588),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_582),
.B(n_246),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_595),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_582),
.B(n_246),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_599),
.B(n_545),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_670),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_595),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_582),
.B(n_250),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_592),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_658),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_636),
.Y(n_708)
);

INVxp67_ASAP7_75t_SL g709 ( 
.A(n_616),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_649),
.B(n_548),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_636),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_670),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_666),
.B(n_562),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_592),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_616),
.B(n_498),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_624),
.B(n_250),
.Y(n_716)
);

INVx6_ASAP7_75t_L g717 ( 
.A(n_658),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_591),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_593),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_593),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_596),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_666),
.B(n_563),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_612),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_596),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_619),
.B(n_555),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_634),
.B(n_574),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_658),
.B(n_573),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_651),
.B(n_490),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_653),
.B(n_501),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_653),
.B(n_501),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_601),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_670),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_634),
.B(n_575),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_670),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_658),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_612),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_624),
.A2(n_637),
.B1(n_517),
.B2(n_579),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_678),
.Y(n_738)
);

AND2x6_ASAP7_75t_L g739 ( 
.A(n_624),
.B(n_351),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_612),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_601),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_670),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_496),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_674),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_606),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_606),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_597),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_608),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_674),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_624),
.A2(n_569),
.B1(n_541),
.B2(n_546),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_607),
.B(n_555),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_614),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_621),
.B(n_513),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_614),
.Y(n_754)
);

AO22x2_ASAP7_75t_L g755 ( 
.A1(n_637),
.A2(n_609),
.B1(n_372),
.B2(n_433),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_607),
.B(n_516),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_614),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_637),
.A2(n_546),
.B1(n_568),
.B2(n_296),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_630),
.B(n_502),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_629),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_637),
.B(n_351),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_674),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_629),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_674),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_610),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_610),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_629),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_674),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_674),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_658),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_630),
.B(n_372),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_621),
.A2(n_558),
.B1(n_455),
.B2(n_422),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_658),
.B(n_411),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_664),
.B(n_585),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_638),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_638),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_642),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_613),
.Y(n_781)
);

INVx5_ASAP7_75t_L g782 ( 
.A(n_603),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_586),
.B(n_532),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_648),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_630),
.B(n_371),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_618),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_609),
.B(n_387),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_674),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_603),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_664),
.B(n_590),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_603),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_626),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_641),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_626),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_645),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_645),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_646),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_642),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_646),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_641),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_650),
.B(n_663),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_650),
.B(n_388),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_619),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_662),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_662),
.B(n_260),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_602),
.Y(n_807)
);

BUFx4f_ASAP7_75t_L g808 ( 
.A(n_594),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_603),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_673),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_603),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_620),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_604),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_603),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_620),
.Y(n_815)
);

AND2x6_ASAP7_75t_L g816 ( 
.A(n_663),
.B(n_372),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_603),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_622),
.B(n_549),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_673),
.A2(n_580),
.B(n_296),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_642),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_623),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_644),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_675),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_659),
.Y(n_824)
);

AND3x4_ASAP7_75t_L g825 ( 
.A(n_587),
.B(n_368),
.C(n_484),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_644),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_675),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_633),
.A2(n_433),
.B(n_565),
.C(n_466),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_594),
.Y(n_829)
);

INVx4_ASAP7_75t_SL g830 ( 
.A(n_625),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_659),
.B(n_502),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_628),
.B(n_550),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_647),
.B(n_389),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_644),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_625),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_594),
.B(n_433),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_625),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_667),
.B(n_352),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_667),
.B(n_360),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_587),
.B(n_360),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_715),
.B(n_632),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_709),
.B(n_635),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_747),
.B(n_639),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_688),
.A2(n_657),
.B(n_429),
.C(n_299),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_735),
.Y(n_845)
);

AND3x1_ASAP7_75t_L g846 ( 
.A(n_775),
.B(n_617),
.C(n_368),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_802),
.A2(n_560),
.B1(n_567),
.B2(n_553),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_729),
.A2(n_730),
.B(n_819),
.C(n_760),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_828),
.A2(n_802),
.B(n_680),
.C(n_819),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_733),
.B(n_640),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_695),
.B(n_643),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_805),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_717),
.B(n_594),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_683),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_683),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_691),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_774),
.A2(n_594),
.B1(n_278),
.B2(n_279),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_684),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_691),
.B(n_652),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_691),
.B(n_729),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_691),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_774),
.A2(n_278),
.B1(n_279),
.B2(n_260),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_808),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_808),
.B(n_654),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_726),
.B(n_660),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_739),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_730),
.B(n_661),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_SL g868 ( 
.A(n_708),
.B(n_677),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_802),
.A2(n_571),
.B1(n_669),
.B2(n_665),
.Y(n_869)
);

BUFx8_ASAP7_75t_L g870 ( 
.A(n_824),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_805),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_R g872 ( 
.A(n_807),
.B(n_672),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_686),
.B(n_676),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_693),
.B(n_617),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_743),
.B(n_256),
.C(n_254),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_808),
.B(n_290),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_679),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_836),
.B(n_290),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_802),
.B(n_647),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_810),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_836),
.B(n_290),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_829),
.A2(n_312),
.B(n_303),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_831),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_802),
.B(n_647),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_810),
.Y(n_885)
);

NOR2x1p5_ASAP7_75t_L g886 ( 
.A(n_708),
.B(n_264),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_823),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_737),
.B(n_647),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_774),
.A2(n_312),
.B1(n_314),
.B2(n_303),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_760),
.B(n_633),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_840),
.B(n_605),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_750),
.A2(n_491),
.B1(n_492),
.B2(n_488),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_774),
.A2(n_324),
.B1(n_329),
.B2(n_314),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_829),
.B(n_324),
.Y(n_894)
);

BUFx12f_ASAP7_75t_L g895 ( 
.A(n_807),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_774),
.A2(n_349),
.B1(n_353),
.B2(n_329),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_803),
.B(n_633),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_701),
.B(n_605),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_836),
.B(n_668),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_823),
.B(n_668),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_827),
.B(n_668),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_827),
.B(n_668),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_698),
.B(n_290),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_786),
.B(n_668),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_698),
.B(n_290),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_831),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_684),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_806),
.B(n_349),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_698),
.B(n_353),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_698),
.B(n_290),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_774),
.A2(n_396),
.B1(n_400),
.B2(n_390),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_685),
.B(n_633),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_700),
.B(n_317),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_685),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_774),
.A2(n_409),
.B1(n_414),
.B2(n_405),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_700),
.B(n_317),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_700),
.B(n_317),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_693),
.A2(n_417),
.B1(n_420),
.B2(n_416),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_687),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_687),
.B(n_633),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_728),
.A2(n_443),
.B1(n_449),
.B2(n_430),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_728),
.B(n_615),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_694),
.B(n_631),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_694),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_L g925 ( 
.A1(n_700),
.A2(n_374),
.B(n_377),
.C(n_370),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_697),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_679),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_697),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_801),
.B(n_615),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_682),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_705),
.B(n_317),
.Y(n_931)
);

OAI221xp5_ASAP7_75t_L g932 ( 
.A1(n_775),
.A2(n_429),
.B1(n_446),
.B2(n_450),
.C(n_425),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_706),
.B(n_631),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_706),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_714),
.B(n_631),
.Y(n_935)
);

BUFx5_ASAP7_75t_L g936 ( 
.A(n_739),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_682),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_801),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_813),
.Y(n_939)
);

CKINVDCx14_ASAP7_75t_R g940 ( 
.A(n_718),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_705),
.B(n_317),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_710),
.B(n_546),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_714),
.B(n_631),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_719),
.B(n_720),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_705),
.A2(n_374),
.B(n_377),
.C(n_370),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_719),
.B(n_631),
.Y(n_946)
);

INVxp33_ASAP7_75t_L g947 ( 
.A(n_838),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_785),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_SL g949 ( 
.A1(n_825),
.A2(n_382),
.B1(n_268),
.B2(n_269),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_720),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_721),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_721),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_724),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_724),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_731),
.B(n_631),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_713),
.B(n_546),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_705),
.A2(n_457),
.B1(n_452),
.B2(n_384),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_731),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_716),
.A2(n_384),
.B1(n_394),
.B2(n_393),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_815),
.B(n_382),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_711),
.B(n_266),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_679),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_776),
.A2(n_727),
.B(n_716),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_716),
.A2(n_393),
.B1(n_395),
.B2(n_394),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_741),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_716),
.B(n_317),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_739),
.B(n_363),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_735),
.B(n_395),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_711),
.B(n_271),
.Y(n_969)
);

AO22x1_ASAP7_75t_L g970 ( 
.A1(n_816),
.A2(n_299),
.B1(n_336),
.B2(n_292),
.Y(n_970)
);

AND2x6_ASAP7_75t_SL g971 ( 
.A(n_784),
.B(n_336),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_833),
.A2(n_656),
.B(n_655),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_722),
.B(n_275),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_759),
.B(n_788),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_741),
.B(n_631),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_745),
.B(n_402),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_745),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_824),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_689),
.B(n_283),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_746),
.B(n_402),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_751),
.B(n_281),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_702),
.B(n_363),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_804),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_806),
.B(n_408),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_813),
.B(n_277),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_746),
.B(n_408),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_689),
.B(n_284),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_739),
.A2(n_442),
.B1(n_444),
.B2(n_447),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_748),
.B(n_442),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_812),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_739),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_748),
.B(n_444),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_739),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_756),
.B(n_447),
.Y(n_994)
);

AND2x2_ASAP7_75t_SL g995 ( 
.A(n_753),
.B(n_363),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_756),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_766),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_702),
.B(n_363),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_L g999 ( 
.A(n_739),
.B(n_363),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_702),
.B(n_363),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_762),
.A2(n_418),
.B1(n_366),
.B2(n_376),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_762),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_762),
.A2(n_277),
.B1(n_318),
.B2(n_386),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_840),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_766),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_725),
.B(n_289),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_734),
.B(n_625),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_767),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_L g1009 ( 
.A(n_777),
.B(n_295),
.C(n_291),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_L g1010 ( 
.A(n_762),
.B(n_625),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_794),
.B(n_283),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_762),
.A2(n_418),
.B1(n_366),
.B2(n_376),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_762),
.A2(n_319),
.B1(n_300),
.B2(n_302),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_767),
.B(n_625),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_L g1015 ( 
.A(n_762),
.B(n_625),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_854),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_883),
.B(n_839),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_854),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_938),
.Y(n_1019)
);

AND2x6_ASAP7_75t_SL g1020 ( 
.A(n_841),
.B(n_818),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_855),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_855),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_856),
.A2(n_707),
.B(n_772),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_856),
.B(n_768),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_860),
.B(n_768),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_849),
.A2(n_791),
.B(n_806),
.C(n_783),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_858),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_858),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_938),
.Y(n_1029)
);

NAND2xp33_ASAP7_75t_L g1030 ( 
.A(n_936),
.B(n_816),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_907),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_907),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_949),
.B(n_757),
.C(n_308),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_939),
.B(n_821),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_924),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_870),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_924),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_863),
.B(n_707),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_926),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_842),
.B(n_832),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_926),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_843),
.B(n_821),
.Y(n_1042)
);

AND2x4_ASAP7_75t_SL g1043 ( 
.A(n_929),
.B(n_806),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_928),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_861),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_995),
.A2(n_816),
.B1(n_755),
.B2(n_783),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_861),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_852),
.B(n_781),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_928),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_1004),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_950),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_871),
.B(n_781),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_866),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_932),
.B(n_310),
.C(n_305),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_851),
.B(n_725),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_995),
.A2(n_816),
.B1(n_755),
.B2(n_793),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_950),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_880),
.B(n_885),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_948),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_983),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_867),
.B(n_838),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_866),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_983),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_908),
.A2(n_816),
.B1(n_755),
.B2(n_793),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_891),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_877),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_958),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_948),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_990),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_899),
.A2(n_707),
.B(n_772),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_866),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_887),
.B(n_787),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_922),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_866),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_L g1075 ( 
.A(n_859),
.B(n_864),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_883),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_864),
.A2(n_816),
.B1(n_755),
.B2(n_795),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_991),
.B(n_717),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_914),
.B(n_787),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_958),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_919),
.B(n_795),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_965),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_870),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_934),
.B(n_796),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_850),
.B(n_865),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_965),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_977),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_977),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_996),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_996),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_997),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_951),
.B(n_796),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_997),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_877),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_870),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_991),
.B(n_797),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_939),
.B(n_738),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_978),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1009),
.B(n_320),
.C(n_311),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_947),
.B(n_839),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_952),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_953),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_993),
.B(n_797),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_866),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_954),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_895),
.Y(n_1106)
);

AND3x2_ASAP7_75t_SL g1107 ( 
.A(n_846),
.B(n_825),
.C(n_348),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_895),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_993),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1002),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1005),
.Y(n_1111)
);

BUFx8_ASAP7_75t_L g1112 ( 
.A(n_873),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1008),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_906),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_906),
.B(n_882),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_872),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_978),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_947),
.B(n_825),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_890),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_908),
.A2(n_816),
.B1(n_798),
.B2(n_800),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_877),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_944),
.B(n_798),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_927),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_908),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_848),
.B(n_800),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1002),
.B(n_734),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_848),
.B(n_734),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_984),
.B(n_742),
.Y(n_1128)
);

AND3x1_ASAP7_75t_SL g1129 ( 
.A(n_886),
.B(n_399),
.C(n_397),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_984),
.B(n_742),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_900),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_978),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_901),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_930),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_902),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_845),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_888),
.A2(n_857),
.B1(n_974),
.B2(n_881),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_984),
.B(n_942),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_927),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_974),
.A2(n_717),
.B1(n_763),
.B2(n_742),
.Y(n_1140)
);

NOR2x1p5_ASAP7_75t_L g1141 ( 
.A(n_874),
.B(n_322),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_912),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_937),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_927),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_962),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_898),
.B(n_326),
.C(n_325),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_845),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_878),
.A2(n_717),
.B1(n_771),
.B2(n_763),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_863),
.B(n_744),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_961),
.B(n_744),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_894),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_962),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_969),
.B(n_744),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_SL g1154 ( 
.A(n_894),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_962),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_909),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_853),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_920),
.Y(n_1158)
);

INVx6_ASAP7_75t_L g1159 ( 
.A(n_845),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1014),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_956),
.B(n_763),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_845),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_923),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_SL g1164 ( 
.A(n_987),
.B(n_331),
.C(n_327),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_894),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1011),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_863),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_963),
.A2(n_792),
.B(n_749),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_933),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_894),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_979),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_894),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_879),
.B(n_771),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_904),
.B(n_771),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_970),
.B(n_884),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_894),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_875),
.B(n_789),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_SL g1178 ( 
.A(n_1006),
.B(n_333),
.C(n_332),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_935),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_868),
.B(n_679),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_878),
.B(n_789),
.Y(n_1181)
);

CKINVDCx8_ASAP7_75t_R g1182 ( 
.A(n_971),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_968),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_943),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_960),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_R g1186 ( 
.A(n_940),
.B(n_789),
.Y(n_1186)
);

OR2x4_ASAP7_75t_L g1187 ( 
.A(n_981),
.B(n_397),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_946),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_955),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_869),
.B(n_679),
.Y(n_1190)
);

CKINVDCx16_ASAP7_75t_R g1191 ( 
.A(n_940),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_881),
.B(n_744),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_909),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_975),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_936),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_973),
.B(n_690),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_SL g1197 ( 
.A(n_876),
.B(n_976),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1007),
.Y(n_1198)
);

CKINVDCx8_ASAP7_75t_R g1199 ( 
.A(n_847),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_980),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_968),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1007),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_985),
.B(n_681),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_897),
.B(n_749),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_986),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_989),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_936),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_892),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_992),
.B(n_749),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_918),
.B(n_749),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_994),
.B(n_765),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1028),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1017),
.B(n_903),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1207),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1085),
.B(n_1040),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1138),
.A2(n_945),
.B(n_925),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_1197),
.A2(n_876),
.B(n_844),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1053),
.A2(n_1015),
.B(n_1010),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1185),
.B(n_921),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1119),
.B(n_936),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1016),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1028),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1031),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1031),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1042),
.A2(n_1003),
.B(n_957),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1109),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1200),
.B(n_959),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1016),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1053),
.A2(n_1015),
.B(n_1010),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1205),
.B(n_964),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1119),
.B(n_1001),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1168),
.A2(n_972),
.B(n_905),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1127),
.A2(n_905),
.B(n_903),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1195),
.B(n_936),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1125),
.A2(n_913),
.B(n_910),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1206),
.B(n_1012),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1032),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1017),
.B(n_910),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1096),
.B(n_936),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1032),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1053),
.A2(n_999),
.B(n_967),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1061),
.A2(n_916),
.B(n_917),
.C(n_913),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1035),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1197),
.A2(n_917),
.B(n_916),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1018),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1115),
.A2(n_889),
.B1(n_893),
.B2(n_862),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1070),
.A2(n_941),
.B(n_931),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1149),
.A2(n_941),
.B(n_931),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1035),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1018),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1021),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1026),
.A2(n_998),
.B(n_982),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1096),
.B(n_936),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1149),
.A2(n_966),
.B(n_982),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1207),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1149),
.A2(n_966),
.B(n_998),
.Y(n_1256)
);

INVxp33_ASAP7_75t_L g1257 ( 
.A(n_1097),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1137),
.A2(n_692),
.A3(n_696),
.B(n_690),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1059),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1038),
.A2(n_1000),
.B(n_837),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1037),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1206),
.B(n_896),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1096),
.B(n_1013),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1192),
.A2(n_915),
.B(n_911),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1101),
.B(n_1000),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1109),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1100),
.A2(n_999),
.B(n_967),
.C(n_988),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1109),
.Y(n_1268)
);

CKINVDCx6p67_ASAP7_75t_R g1269 ( 
.A(n_1106),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1150),
.B(n_692),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1153),
.B(n_696),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1038),
.A2(n_837),
.B(n_809),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1101),
.B(n_699),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1122),
.B(n_699),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_SL g1275 ( 
.A(n_1116),
.B(n_283),
.Y(n_1275)
);

NAND2x1_ASAP7_75t_L g1276 ( 
.A(n_1207),
.B(n_681),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1021),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1062),
.A2(n_792),
.B(n_770),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1073),
.B(n_334),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1102),
.A2(n_404),
.B(n_410),
.C(n_399),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1102),
.B(n_703),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1105),
.B(n_703),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1105),
.B(n_704),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1140),
.A2(n_834),
.A3(n_826),
.B(n_822),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1038),
.A2(n_837),
.B(n_809),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1037),
.A2(n_834),
.A3(n_826),
.B(n_822),
.Y(n_1286)
);

INVx8_ASAP7_75t_L g1287 ( 
.A(n_1078),
.Y(n_1287)
);

INVx4_ASAP7_75t_L g1288 ( 
.A(n_1109),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1077),
.A2(n_723),
.B(n_704),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1111),
.B(n_723),
.Y(n_1290)
);

AOI221xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1055),
.A2(n_413),
.B1(n_446),
.B2(n_404),
.C(n_410),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1046),
.A2(n_809),
.B1(n_770),
.B2(n_765),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1161),
.A2(n_740),
.B(n_736),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1059),
.Y(n_1294)
);

NAND3xp33_ASAP7_75t_SL g1295 ( 
.A(n_1199),
.B(n_339),
.C(n_337),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1022),
.Y(n_1296)
);

NAND2x1_ASAP7_75t_L g1297 ( 
.A(n_1207),
.B(n_681),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1068),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1023),
.A2(n_740),
.B(n_736),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1111),
.B(n_752),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1181),
.A2(n_754),
.B(n_752),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1062),
.A2(n_792),
.B(n_770),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1062),
.A2(n_792),
.B(n_770),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1022),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1116),
.B(n_348),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1174),
.A2(n_758),
.B(n_754),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1065),
.B(n_345),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1025),
.B(n_758),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1167),
.A2(n_764),
.B(n_761),
.Y(n_1309)
);

O2A1O1Ixp5_ASAP7_75t_L g1310 ( 
.A1(n_1203),
.A2(n_761),
.B(n_764),
.C(n_820),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1071),
.A2(n_1104),
.B(n_1074),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1056),
.A2(n_773),
.B(n_769),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1109),
.A2(n_1110),
.B1(n_1120),
.B2(n_1103),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1196),
.B(n_769),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1050),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1196),
.B(n_1076),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1071),
.A2(n_765),
.B(n_790),
.Y(n_1317)
);

OAI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1034),
.A2(n_357),
.B(n_347),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1039),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1167),
.A2(n_778),
.B(n_773),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1047),
.B(n_765),
.Y(n_1321)
);

NAND2x1_ASAP7_75t_L g1322 ( 
.A(n_1071),
.B(n_1074),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1210),
.A2(n_1064),
.B(n_1131),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1167),
.A2(n_779),
.B(n_778),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1076),
.B(n_779),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1074),
.A2(n_811),
.B(n_790),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1051),
.Y(n_1327)
);

O2A1O1Ixp5_ASAP7_75t_L g1328 ( 
.A1(n_1190),
.A2(n_820),
.B(n_780),
.C(n_799),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1195),
.A2(n_799),
.B(n_780),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_SL g1330 ( 
.A(n_1199),
.B(n_359),
.C(n_358),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1104),
.A2(n_811),
.B(n_790),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1039),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1114),
.B(n_681),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1195),
.A2(n_508),
.B(n_506),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1051),
.A2(n_413),
.A3(n_425),
.B(n_450),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1103),
.B(n_1156),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1131),
.A2(n_1135),
.B(n_1133),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1204),
.A2(n_508),
.B(n_506),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1114),
.B(n_681),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1043),
.B(n_576),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1104),
.A2(n_811),
.B(n_790),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1058),
.B(n_712),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1176),
.A2(n_512),
.B(n_511),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1106),
.B(n_348),
.Y(n_1344)
);

AOI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1075),
.A2(n_1086),
.B(n_1057),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1133),
.A2(n_656),
.B(n_655),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1176),
.A2(n_512),
.B(n_511),
.Y(n_1347)
);

AOI221x1_ASAP7_75t_L g1348 ( 
.A1(n_1163),
.A2(n_577),
.B1(n_578),
.B2(n_518),
.C(n_556),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1057),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1124),
.A2(n_578),
.B(n_577),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1135),
.A2(n_656),
.B(n_655),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1050),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1156),
.A2(n_439),
.B(n_361),
.C(n_362),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1030),
.A2(n_811),
.B(n_790),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1118),
.A2(n_712),
.B1(n_732),
.B2(n_817),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1110),
.A2(n_712),
.B1(n_732),
.B2(n_817),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1177),
.A2(n_830),
.B(n_373),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1030),
.A2(n_1211),
.B(n_1209),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1086),
.A2(n_518),
.A3(n_523),
.B(n_525),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1103),
.B(n_712),
.Y(n_1360)
);

AOI31xp67_ASAP7_75t_L g1361 ( 
.A1(n_1044),
.A2(n_830),
.A3(n_835),
.B(n_817),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1113),
.B(n_712),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1176),
.A2(n_525),
.B(n_523),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1142),
.B(n_732),
.Y(n_1364)
);

AOI221x1_ASAP7_75t_L g1365 ( 
.A1(n_1163),
.A2(n_556),
.B1(n_528),
.B2(n_530),
.C(n_531),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1166),
.B(n_367),
.C(n_364),
.Y(n_1366)
);

AOI211x1_ASAP7_75t_L g1367 ( 
.A1(n_1048),
.A2(n_559),
.B(n_551),
.C(n_547),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1088),
.A2(n_1091),
.B(n_1089),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1088),
.A2(n_1091),
.B(n_1089),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1148),
.A2(n_528),
.B(n_526),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1157),
.A2(n_1049),
.B(n_1044),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1110),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1179),
.A2(n_526),
.A3(n_530),
.B(n_531),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1110),
.B(n_732),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1049),
.Y(n_1375)
);

AOI211x1_ASAP7_75t_L g1376 ( 
.A1(n_1052),
.A2(n_559),
.B(n_551),
.C(n_547),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1142),
.B(n_732),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1047),
.B(n_830),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1158),
.A2(n_600),
.B(n_611),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1158),
.A2(n_1173),
.B(n_1179),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1067),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1371),
.A2(n_1320),
.B(n_1309),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1371),
.A2(n_1157),
.B(n_1087),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1358),
.A2(n_1156),
.B(n_1157),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1215),
.A2(n_1024),
.B(n_1180),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1269),
.Y(n_1386)
);

OAI22x1_ASAP7_75t_L g1387 ( 
.A1(n_1345),
.A2(n_1141),
.B1(n_1208),
.B2(n_1171),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1217),
.A2(n_1194),
.A3(n_1087),
.B(n_1090),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1368),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1352),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1275),
.A2(n_1208),
.B1(n_1187),
.B2(n_1063),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1259),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1267),
.A2(n_1079),
.B(n_1072),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1221),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1369),
.Y(n_1395)
);

AO22x1_ASAP7_75t_L g1396 ( 
.A1(n_1323),
.A2(n_1112),
.B1(n_1201),
.B2(n_1193),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1309),
.A2(n_1090),
.B(n_1067),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1306),
.A2(n_1244),
.B(n_1293),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1225),
.A2(n_1146),
.B(n_1178),
.C(n_1134),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1226),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1348),
.A2(n_1194),
.A3(n_1093),
.B(n_1041),
.Y(n_1401)
);

AOI21xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1219),
.A2(n_1191),
.B(n_1069),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1306),
.A2(n_1080),
.B(n_1027),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1259),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1221),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1268),
.B(n_1047),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1228),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1316),
.B(n_1043),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1270),
.A2(n_1165),
.B(n_1151),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1320),
.A2(n_1324),
.B(n_1285),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1267),
.A2(n_1084),
.B(n_1081),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1228),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1315),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1336),
.B(n_1124),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_SL g1416 ( 
.A1(n_1380),
.A2(n_1092),
.B(n_1093),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1336),
.B(n_1128),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1245),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1324),
.A2(n_1160),
.B(n_1082),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1213),
.B(n_1169),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1337),
.A2(n_1264),
.B(n_1233),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1245),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1250),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_SL g1424 ( 
.A1(n_1220),
.A2(n_1198),
.B(n_1019),
.C(n_1029),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1272),
.A2(n_1160),
.B(n_1169),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1365),
.A2(n_1188),
.B(n_1184),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_SL g1427 ( 
.A1(n_1220),
.A2(n_1263),
.B(n_1353),
.C(n_1231),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1250),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1233),
.A2(n_1262),
.B(n_1235),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1370),
.A2(n_1188),
.B(n_1184),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1272),
.A2(n_1189),
.B(n_1094),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1251),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1213),
.B(n_1019),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1293),
.A2(n_1289),
.B(n_1232),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1238),
.B(n_1029),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1287),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1277),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1235),
.A2(n_1175),
.B(n_1173),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1294),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1295),
.A2(n_1107),
.B(n_1095),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1277),
.Y(n_1442)
);

AO31x2_ASAP7_75t_L g1443 ( 
.A1(n_1280),
.A2(n_1189),
.A3(n_1151),
.B(n_1165),
.Y(n_1443)
);

AOI221x1_ASAP7_75t_L g1444 ( 
.A1(n_1353),
.A2(n_1177),
.B1(n_1173),
.B2(n_1198),
.C(n_1172),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1214),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1296),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1285),
.A2(n_1094),
.B(n_1066),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1296),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1329),
.A2(n_1094),
.B(n_1066),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1242),
.A2(n_1054),
.B(n_1033),
.C(n_1099),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1304),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1304),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1319),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1238),
.B(n_1128),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1214),
.B(n_1128),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1313),
.A2(n_1110),
.B1(n_1045),
.B2(n_1170),
.Y(n_1456)
);

NAND2x1_ASAP7_75t_L g1457 ( 
.A(n_1234),
.B(n_1147),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1319),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1329),
.A2(n_1123),
.B(n_1066),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1260),
.A2(n_1144),
.B(n_1123),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1293),
.A2(n_1177),
.B(n_1139),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1260),
.A2(n_1144),
.B(n_1123),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1287),
.B(n_1183),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1334),
.A2(n_1152),
.B(n_1144),
.Y(n_1464)
);

OAI21xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1312),
.A2(n_1202),
.B(n_1078),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1257),
.B(n_1020),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1307),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1298),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1232),
.A2(n_1338),
.B(n_1271),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1332),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1332),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1330),
.A2(n_1164),
.B1(n_1143),
.B2(n_431),
.C(n_436),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1273),
.B(n_1340),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1307),
.B(n_1305),
.C(n_1279),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1334),
.A2(n_1155),
.B(n_1152),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1357),
.A2(n_1155),
.B(n_1152),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1314),
.B(n_1175),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1381),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1236),
.A2(n_1175),
.B(n_1130),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1370),
.A2(n_1202),
.B(n_1139),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1273),
.B(n_1340),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1227),
.A2(n_1045),
.B1(n_1170),
.B2(n_1063),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1265),
.B(n_1130),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1287),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1269),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1298),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1291),
.A2(n_1145),
.B(n_1121),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1214),
.B(n_1130),
.Y(n_1488)
);

AOI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1354),
.A2(n_1175),
.B(n_1145),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_SL g1490 ( 
.A(n_1263),
.B(n_1183),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1343),
.A2(n_1155),
.B(n_1121),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1343),
.A2(n_539),
.B(n_538),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1381),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1280),
.A2(n_1147),
.A3(n_1187),
.B(n_539),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1375),
.Y(n_1495)
);

AO32x2_ASAP7_75t_L g1496 ( 
.A1(n_1246),
.A2(n_1147),
.A3(n_1187),
.B1(n_1129),
.B2(n_1069),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1347),
.A2(n_1363),
.B(n_1247),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1212),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1255),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_SL g1500 ( 
.A1(n_1218),
.A2(n_1154),
.B(n_1172),
.Y(n_1500)
);

AO221x2_ASAP7_75t_L g1501 ( 
.A1(n_1366),
.A2(n_1107),
.B1(n_421),
.B2(n_373),
.C(n_348),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1279),
.A2(n_1045),
.B1(n_1060),
.B2(n_1068),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1347),
.A2(n_542),
.B(n_538),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1287),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1344),
.A2(n_1112),
.B1(n_1117),
.B2(n_1083),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1363),
.A2(n_543),
.B(n_542),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1230),
.A2(n_1112),
.B1(n_1117),
.B2(n_1083),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1257),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1255),
.Y(n_1509)
);

AO32x2_ASAP7_75t_L g1510 ( 
.A1(n_1258),
.A2(n_1107),
.A3(n_1154),
.B1(n_1183),
.B2(n_1201),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1222),
.A2(n_1060),
.B1(n_1143),
.B2(n_1108),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1223),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1265),
.B(n_1224),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1346),
.A2(n_543),
.B(n_1126),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1237),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1240),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1243),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1249),
.B(n_1126),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1255),
.B(n_1045),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1268),
.B(n_1288),
.Y(n_1520)
);

AO21x2_ASAP7_75t_L g1521 ( 
.A1(n_1338),
.A2(n_1126),
.B(n_1186),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1338),
.A2(n_1154),
.B(n_1183),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1241),
.A2(n_1183),
.B(n_1172),
.C(n_1045),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1261),
.B(n_1078),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1318),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1367),
.B(n_1078),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1247),
.A2(n_600),
.B(n_611),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1299),
.A2(n_600),
.B(n_611),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1274),
.B(n_1136),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1299),
.A2(n_600),
.B(n_611),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1226),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_SL g1532 ( 
.A1(n_1229),
.A2(n_1172),
.B(n_1159),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1308),
.A2(n_1162),
.B(n_1136),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1355),
.A2(n_1182),
.B1(n_1108),
.B2(n_1098),
.C(n_1095),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1327),
.Y(n_1535)
);

BUFx2_ASAP7_75t_R g1536 ( 
.A(n_1360),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1349),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1226),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1281),
.Y(n_1539)
);

AND2x4_ASAP7_75t_SL g1540 ( 
.A(n_1268),
.B(n_1172),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1282),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1283),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_SL g1543 ( 
.A1(n_1239),
.A2(n_1159),
.B(n_1162),
.C(n_129),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1335),
.B(n_1325),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1290),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1254),
.A2(n_600),
.B(n_611),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1351),
.A2(n_423),
.B(n_419),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1335),
.B(n_1372),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1226),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1300),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1254),
.A2(n_1256),
.B(n_1248),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1359),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1288),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1266),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1239),
.A2(n_1159),
.B1(n_1098),
.B2(n_1182),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1256),
.A2(n_1159),
.B(n_830),
.Y(n_1556)
);

AOI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1362),
.A2(n_1132),
.B(n_1036),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1253),
.A2(n_1036),
.B1(n_1132),
.B2(n_1360),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1248),
.A2(n_432),
.B(n_375),
.C(n_378),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1328),
.A2(n_381),
.B(n_369),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1253),
.A2(n_373),
.B1(n_421),
.B2(n_437),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1359),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1288),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1321),
.A2(n_435),
.B1(n_380),
.B2(n_383),
.Y(n_1564)
);

AO21x2_ASAP7_75t_L g1565 ( 
.A1(n_1379),
.A2(n_835),
.B(n_817),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1216),
.A2(n_835),
.B(n_817),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1335),
.B(n_373),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1301),
.A2(n_835),
.B(n_814),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1474),
.A2(n_1350),
.B1(n_421),
.B2(n_437),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1390),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1384),
.A2(n_1252),
.B(n_1342),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1421),
.A2(n_1252),
.B(n_1311),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1534),
.A2(n_428),
.B1(n_427),
.B2(n_456),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1437),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1523),
.A2(n_1252),
.B(n_1292),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1536),
.A2(n_1376),
.B1(n_1266),
.B2(n_1377),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1404),
.Y(n_1577)
);

OAI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1467),
.A2(n_438),
.B1(n_403),
.B2(n_406),
.C(n_454),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1525),
.A2(n_1321),
.B1(n_398),
.B2(n_407),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1404),
.B(n_1266),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1437),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1502),
.A2(n_1266),
.B1(n_1364),
.B2(n_1374),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1382),
.A2(n_1530),
.B(n_1528),
.Y(n_1583)
);

AOI22x1_ASAP7_75t_L g1584 ( 
.A1(n_1387),
.A2(n_1374),
.B1(n_1321),
.B2(n_1378),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1486),
.B(n_1378),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_SL g1586 ( 
.A1(n_1450),
.A2(n_1339),
.B(n_1333),
.C(n_1322),
.Y(n_1586)
);

AOI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1477),
.A2(n_1310),
.B(n_1356),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_L g1588 ( 
.A(n_1525),
.B(n_1234),
.Y(n_1588)
);

AOI222xp33_ASAP7_75t_L g1589 ( 
.A1(n_1391),
.A2(n_437),
.B1(n_421),
.B2(n_448),
.C1(n_453),
.C2(n_434),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1386),
.B(n_1378),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1413),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1498),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1390),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1473),
.B(n_1335),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_SL g1595 ( 
.A1(n_1559),
.A2(n_1297),
.B(n_1276),
.C(n_1341),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1508),
.A2(n_385),
.B1(n_451),
.B2(n_1278),
.Y(n_1596)
);

NOR2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1504),
.B(n_437),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1437),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1515),
.Y(n_1599)
);

INVx4_ASAP7_75t_SL g1600 ( 
.A(n_1437),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1434),
.B(n_1373),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1399),
.A2(n_1331),
.B(n_1326),
.C(n_1317),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1486),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1386),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1501),
.A2(n_1234),
.B1(n_1303),
.B2(n_1302),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1437),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1515),
.A2(n_1234),
.B1(n_1361),
.B2(n_12),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1535),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1444),
.A2(n_1258),
.B(n_1284),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1501),
.A2(n_1234),
.B1(n_10),
.B2(n_12),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1501),
.A2(n_1234),
.B1(n_811),
.B2(n_814),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1512),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1501),
.A2(n_7),
.B1(n_14),
.B2(n_15),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1463),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1466),
.A2(n_814),
.B1(n_835),
.B2(n_627),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1535),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1473),
.B(n_1359),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1455),
.B(n_1488),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1516),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1485),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1481),
.B(n_1359),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1387),
.A2(n_814),
.B1(n_627),
.B2(n_1373),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1441),
.A2(n_814),
.B1(n_627),
.B2(n_782),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1382),
.A2(n_1284),
.B(n_1258),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1537),
.A2(n_15),
.B1(n_16),
.B2(n_20),
.Y(n_1625)
);

BUFx12f_ASAP7_75t_L g1626 ( 
.A(n_1415),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1504),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1537),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1561),
.A2(n_1373),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1517),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1472),
.A2(n_627),
.B1(n_1373),
.B2(n_782),
.Y(n_1631)
);

AND2x2_ASAP7_75t_SL g1632 ( 
.A(n_1484),
.B(n_21),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1415),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1490),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1481),
.B(n_1286),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1454),
.A2(n_627),
.B1(n_782),
.B2(n_1258),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1517),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1392),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1528),
.A2(n_1284),
.B(n_1286),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1436),
.B(n_116),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1413),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1440),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1454),
.B(n_1286),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1507),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_1644)
);

AO31x2_ASAP7_75t_L g1645 ( 
.A1(n_1444),
.A2(n_1284),
.A3(n_1286),
.B(n_36),
.Y(n_1645)
);

INVx5_ASAP7_75t_L g1646 ( 
.A(n_1463),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1483),
.B(n_31),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1420),
.B(n_33),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1468),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1484),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1495),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1402),
.B(n_125),
.Y(n_1652)
);

INVx4_ASAP7_75t_SL g1653 ( 
.A(n_1484),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1558),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1463),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1479),
.A2(n_627),
.B1(n_782),
.B2(n_42),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1484),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1414),
.A2(n_627),
.B1(n_782),
.B2(n_43),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1539),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1393),
.A2(n_782),
.B(n_229),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1455),
.B(n_223),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1411),
.A2(n_222),
.B(n_209),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1495),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1429),
.A2(n_200),
.B(n_196),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1539),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1665)
);

BUFx8_ASAP7_75t_L g1666 ( 
.A(n_1484),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1455),
.B(n_193),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1483),
.B(n_49),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1455),
.B(n_189),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1402),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1531),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1420),
.B(n_56),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1505),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1465),
.A2(n_188),
.B(n_185),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1488),
.B(n_1417),
.Y(n_1675)
);

NAND4xp25_ASAP7_75t_L g1676 ( 
.A(n_1564),
.B(n_57),
.C(n_58),
.D(n_59),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1519),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1488),
.B(n_183),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1477),
.B(n_58),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1518),
.Y(n_1680)
);

BUFx8_ASAP7_75t_L g1681 ( 
.A(n_1549),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1520),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1414),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1683)
);

AOI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1567),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.C1(n_64),
.C2(n_71),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1541),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_1685)
);

AOI21xp33_ASAP7_75t_L g1686 ( 
.A1(n_1385),
.A2(n_76),
.B(n_77),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1488),
.B(n_179),
.Y(n_1687)
);

AND2x2_ASAP7_75t_SL g1688 ( 
.A(n_1414),
.B(n_78),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1414),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1412),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1520),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1409),
.A2(n_158),
.B(n_157),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1417),
.B(n_156),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1394),
.Y(n_1694)
);

AND2x6_ASAP7_75t_L g1695 ( 
.A(n_1520),
.B(n_151),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1417),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1490),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1518),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1418),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1520),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1417),
.B(n_145),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1530),
.A2(n_143),
.B(n_138),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1519),
.B(n_87),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1408),
.B(n_88),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1423),
.Y(n_1705)
);

NAND2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1555),
.B(n_88),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1549),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1567),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1526),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_1709)
);

NAND2x1p5_ASAP7_75t_L g1710 ( 
.A(n_1553),
.B(n_95),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1541),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_1711)
);

OAI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1511),
.A2(n_101),
.B1(n_1482),
.B2(n_1526),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1549),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1465),
.A2(n_1557),
.B(n_1439),
.C(n_1560),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1526),
.A2(n_101),
.B1(n_1524),
.B2(n_1513),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1423),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1463),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1553),
.B(n_1563),
.Y(n_1718)
);

AOI222xp33_ASAP7_75t_L g1719 ( 
.A1(n_1513),
.A2(n_1396),
.B1(n_1550),
.B2(n_1545),
.C1(n_1542),
.C2(n_1524),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1445),
.B(n_1499),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1446),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1519),
.B(n_1406),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1446),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1396),
.A2(n_1456),
.B1(n_1519),
.B2(n_1427),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1526),
.B(n_1500),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1544),
.A2(n_1416),
.B1(n_1550),
.B2(n_1545),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1549),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1542),
.B(n_1529),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1435),
.A2(n_1457),
.B(n_1514),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1435),
.A2(n_1457),
.B(n_1514),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1452),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1553),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1400),
.Y(n_1733)
);

BUFx2_ASAP7_75t_SL g1734 ( 
.A(n_1549),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1406),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1540),
.B(n_1445),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1400),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1544),
.A2(n_1416),
.B1(n_1547),
.B2(n_1548),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1548),
.B(n_1494),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_R g1741 ( 
.A(n_1547),
.B(n_1445),
.Y(n_1741)
);

BUFx12f_ASAP7_75t_L g1742 ( 
.A(n_1538),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1743)
);

CKINVDCx16_ASAP7_75t_R g1744 ( 
.A(n_1554),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1499),
.A2(n_1509),
.B1(n_1543),
.B2(n_1533),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1563),
.Y(n_1746)
);

NOR3xp33_ASAP7_75t_SL g1747 ( 
.A(n_1552),
.B(n_1562),
.C(n_1453),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1478),
.B(n_1493),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1509),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1494),
.B(n_1509),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1435),
.A2(n_1514),
.B(n_1469),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1478),
.B(n_1493),
.Y(n_1752)
);

AO31x2_ASAP7_75t_L g1753 ( 
.A1(n_1552),
.A2(n_1562),
.A3(n_1395),
.B(n_1389),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1394),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1547),
.A2(n_1389),
.B1(n_1395),
.B2(n_1521),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1514),
.A2(n_1438),
.B1(n_1442),
.B2(n_1433),
.Y(n_1756)
);

AO32x2_ASAP7_75t_L g1757 ( 
.A1(n_1510),
.A2(n_1496),
.A3(n_1388),
.B1(n_1401),
.B2(n_1443),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1424),
.A2(n_1442),
.B1(n_1458),
.B2(n_1451),
.C(n_1448),
.Y(n_1758)
);

BUFx12f_ASAP7_75t_L g1759 ( 
.A(n_1540),
.Y(n_1759)
);

CKINVDCx6p67_ASAP7_75t_R g1760 ( 
.A(n_1494),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1547),
.A2(n_1521),
.B1(n_1500),
.B2(n_1532),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1563),
.Y(n_1762)
);

CKINVDCx6p67_ASAP7_75t_R g1763 ( 
.A(n_1494),
.Y(n_1763)
);

OAI211xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1405),
.A2(n_1438),
.B(n_1432),
.C(n_1448),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1521),
.A2(n_1532),
.B1(n_1522),
.B2(n_1487),
.Y(n_1765)
);

OAI222xp33_ASAP7_75t_L g1766 ( 
.A1(n_1407),
.A2(n_1433),
.B1(n_1422),
.B2(n_1471),
.C1(n_1470),
.C2(n_1458),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1407),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1589),
.A2(n_1676),
.B1(n_1613),
.B2(n_1610),
.C(n_1578),
.Y(n_1768)
);

OAI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1589),
.A2(n_1496),
.B(n_1489),
.C(n_1428),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1676),
.A2(n_1487),
.B1(n_1470),
.B2(n_1432),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1578),
.A2(n_1489),
.B1(n_1428),
.B2(n_1471),
.C(n_1422),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1684),
.A2(n_1487),
.B1(n_1461),
.B2(n_1426),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1670),
.B(n_1487),
.C(n_1426),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1753),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1577),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1660),
.A2(n_1522),
.B(n_1469),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1579),
.A2(n_1426),
.B1(n_1430),
.B2(n_1480),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1608),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1688),
.B(n_1496),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1684),
.A2(n_1461),
.B1(n_1426),
.B2(n_1522),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1647),
.B(n_1496),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1706),
.A2(n_1461),
.B1(n_1469),
.B2(n_1565),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1616),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1476),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1668),
.B(n_1496),
.Y(n_1785)
);

INVx3_ASAP7_75t_SL g1786 ( 
.A(n_1604),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1675),
.B(n_1443),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1594),
.B(n_1510),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1644),
.A2(n_1565),
.B1(n_1398),
.B2(n_1403),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1709),
.A2(n_1403),
.B1(n_1430),
.B2(n_1480),
.C(n_1510),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1644),
.A2(n_1565),
.B1(n_1398),
.B2(n_1403),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1654),
.A2(n_1398),
.B1(n_1403),
.B2(n_1430),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1728),
.B(n_1388),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1569),
.A2(n_1430),
.B1(n_1480),
.B2(n_1510),
.C(n_1443),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1620),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1728),
.B(n_1388),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1626),
.Y(n_1797)
);

AOI222xp33_ASAP7_75t_L g1798 ( 
.A1(n_1654),
.A2(n_1476),
.B1(n_1419),
.B2(n_1397),
.C1(n_1425),
.C2(n_1506),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1652),
.A2(n_1480),
.B1(n_1419),
.B2(n_1425),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1686),
.A2(n_1510),
.B1(n_1443),
.B2(n_1388),
.C(n_1401),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1673),
.A2(n_1573),
.B1(n_1597),
.B2(n_1712),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1648),
.B(n_1388),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_SL g1803 ( 
.A1(n_1632),
.A2(n_1568),
.B1(n_1383),
.B2(n_1443),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1675),
.B(n_1460),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1629),
.A2(n_1568),
.B1(n_1383),
.B2(n_1431),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1648),
.B(n_1401),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1715),
.A2(n_1462),
.B1(n_1460),
.B2(n_1475),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1703),
.B(n_1401),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1656),
.A2(n_1462),
.B1(n_1464),
.B2(n_1475),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1628),
.Y(n_1810)
);

OAI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1629),
.A2(n_1401),
.B1(n_1397),
.B2(n_1464),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1625),
.A2(n_1503),
.B1(n_1506),
.B2(n_1492),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1649),
.A2(n_1556),
.B1(n_1449),
.B2(n_1459),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_L g1814 ( 
.A(n_1708),
.B(n_1679),
.C(n_1689),
.D(n_1683),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1686),
.A2(n_1503),
.B1(n_1492),
.B2(n_1566),
.Y(n_1815)
);

BUFx4f_ASAP7_75t_SL g1816 ( 
.A(n_1627),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1659),
.A2(n_1527),
.B1(n_1551),
.B2(n_1566),
.C(n_1546),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1640),
.A2(n_1556),
.B1(n_1447),
.B2(n_1449),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1641),
.Y(n_1819)
);

AOI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1659),
.A2(n_1527),
.B1(n_1551),
.B2(n_1546),
.C(n_1431),
.Y(n_1820)
);

OAI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1696),
.A2(n_1497),
.B(n_1447),
.C(n_1459),
.Y(n_1821)
);

OA21x2_ASAP7_75t_L g1822 ( 
.A1(n_1751),
.A2(n_1497),
.B(n_1410),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1623),
.A2(n_1410),
.B1(n_1491),
.B2(n_1680),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1698),
.A2(n_1491),
.B1(n_1591),
.B2(n_1638),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1634),
.A2(n_1697),
.B(n_1662),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1724),
.A2(n_1717),
.B1(n_1658),
.B2(n_1704),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1672),
.B(n_1570),
.Y(n_1827)
);

AND2x4_ASAP7_75t_SL g1828 ( 
.A(n_1603),
.B(n_1585),
.Y(n_1828)
);

AND2x6_ASAP7_75t_L g1829 ( 
.A(n_1693),
.B(n_1701),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1625),
.A2(n_1665),
.B1(n_1685),
.B2(n_1711),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1726),
.A2(n_1622),
.B1(n_1593),
.B2(n_1633),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1677),
.B(n_1600),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1584),
.A2(n_1714),
.B1(n_1672),
.B2(n_1642),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1665),
.A2(n_1711),
.B1(n_1685),
.B2(n_1662),
.C(n_1660),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1618),
.B(n_1612),
.Y(n_1835)
);

OAI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1674),
.A2(n_1692),
.B1(n_1631),
.B2(n_1605),
.C(n_1710),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1601),
.B(n_1617),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1674),
.A2(n_1695),
.B1(n_1621),
.B2(n_1703),
.Y(n_1838)
);

BUFx4f_ASAP7_75t_SL g1839 ( 
.A(n_1742),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1619),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1753),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1618),
.B(n_1643),
.Y(n_1842)
);

AOI222xp33_ASAP7_75t_L g1843 ( 
.A1(n_1588),
.A2(n_1695),
.B1(n_1576),
.B2(n_1596),
.C1(n_1635),
.C2(n_1701),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1576),
.A2(n_1611),
.B1(n_1646),
.B2(n_1738),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1671),
.B(n_1693),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1575),
.A2(n_1602),
.B(n_1590),
.C(n_1572),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1710),
.A2(n_1745),
.B1(n_1761),
.B2(n_1615),
.C(n_1719),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1695),
.A2(n_1719),
.B1(n_1661),
.B2(n_1678),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1603),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1603),
.Y(n_1850)
);

NOR2x1_ASAP7_75t_SL g1851 ( 
.A(n_1646),
.B(n_1725),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1575),
.A2(n_1587),
.B1(n_1755),
.B2(n_1572),
.C(n_1586),
.Y(n_1852)
);

AOI21xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1650),
.A2(n_1687),
.B(n_1667),
.Y(n_1853)
);

BUFx2_ASAP7_75t_R g1854 ( 
.A(n_1734),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1695),
.A2(n_1667),
.B1(n_1661),
.B2(n_1687),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1630),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1637),
.B(n_1651),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_SL g1858 ( 
.A1(n_1646),
.A2(n_1607),
.B1(n_1664),
.B2(n_1614),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1759),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1690),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1571),
.A2(n_1607),
.B(n_1595),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1571),
.A2(n_1729),
.B(n_1730),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1587),
.A2(n_1582),
.B1(n_1735),
.B2(n_1636),
.C(n_1741),
.Y(n_1863)
);

OAI211xp5_ASAP7_75t_L g1864 ( 
.A1(n_1664),
.A2(n_1663),
.B(n_1758),
.C(n_1747),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1646),
.A2(n_1614),
.B1(n_1655),
.B2(n_1725),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1580),
.B(n_1733),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1748),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1655),
.A2(n_1740),
.B1(n_1669),
.B2(n_1678),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1669),
.A2(n_1764),
.B1(n_1721),
.B2(n_1731),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1666),
.A2(n_1582),
.B1(n_1725),
.B2(n_1700),
.Y(n_1870)
);

AOI211x1_ASAP7_75t_L g1871 ( 
.A1(n_1766),
.A2(n_1739),
.B(n_1752),
.C(n_1705),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1749),
.B(n_1574),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1699),
.A2(n_1716),
.B1(n_1723),
.B2(n_1767),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1760),
.A2(n_1763),
.B1(n_1758),
.B2(n_1694),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1707),
.Y(n_1876)
);

AO31x2_ASAP7_75t_L g1877 ( 
.A1(n_1751),
.A2(n_1730),
.A3(n_1729),
.B(n_1756),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1754),
.B(n_1720),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1739),
.B(n_1752),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1574),
.B(n_1581),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1645),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1581),
.B(n_1606),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1743),
.A2(n_1750),
.B1(n_1722),
.B2(n_1691),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1756),
.Y(n_1884)
);

CKINVDCx8_ASAP7_75t_R g1885 ( 
.A(n_1600),
.Y(n_1885)
);

INVx5_ASAP7_75t_L g1886 ( 
.A(n_1746),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1645),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1645),
.Y(n_1888)
);

AOI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1624),
.A2(n_1639),
.B(n_1702),
.Y(n_1889)
);

OAI211xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1765),
.A2(n_1606),
.B(n_1598),
.C(n_1691),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1681),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1598),
.B(n_1682),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1682),
.B(n_1700),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1707),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1737),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_1657),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_SL g1897 ( 
.A1(n_1666),
.A2(n_1681),
.B1(n_1722),
.B2(n_1609),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1718),
.A2(n_1732),
.B(n_1736),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1657),
.A2(n_1736),
.B1(n_1609),
.B2(n_1732),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1657),
.A2(n_1737),
.B1(n_1762),
.B2(n_1746),
.Y(n_1900)
);

INVx8_ASAP7_75t_L g1901 ( 
.A(n_1707),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1737),
.A2(n_1762),
.B1(n_1727),
.B2(n_1713),
.C(n_1718),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1600),
.A2(n_1653),
.B1(n_1727),
.B2(n_1713),
.Y(n_1903)
);

OAI211xp5_ASAP7_75t_L g1904 ( 
.A1(n_1713),
.A2(n_1757),
.B(n_1583),
.C(n_1653),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1653),
.B(n_1757),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1757),
.A2(n_1215),
.B1(n_1676),
.B2(n_1085),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1753),
.Y(n_1907)
);

INVx6_ASAP7_75t_L g1908 ( 
.A(n_1666),
.Y(n_1908)
);

AOI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1578),
.A2(n_1085),
.B1(n_1215),
.B2(n_841),
.C(n_1676),
.Y(n_1909)
);

BUFx12f_ASAP7_75t_L g1910 ( 
.A(n_1620),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1579),
.A2(n_1085),
.B1(n_1215),
.B2(n_1474),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1626),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1589),
.A2(n_1085),
.B1(n_1215),
.B2(n_1676),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1728),
.B(n_1085),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1589),
.A2(n_1085),
.B1(n_1215),
.B2(n_1676),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1706),
.A2(n_1085),
.B1(n_841),
.B2(n_1040),
.Y(n_1916)
);

OR2x6_ASAP7_75t_L g1917 ( 
.A(n_1725),
.B(n_1674),
.Y(n_1917)
);

OAI211xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1589),
.A2(n_1085),
.B(n_1670),
.C(n_1215),
.Y(n_1918)
);

AO22x1_ASAP7_75t_L g1919 ( 
.A1(n_1644),
.A2(n_1085),
.B1(n_841),
.B2(n_850),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1675),
.B(n_1677),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1599),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1753),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1589),
.A2(n_1085),
.B1(n_841),
.B2(n_1040),
.C(n_1215),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1579),
.A2(n_1085),
.B1(n_1215),
.B2(n_1474),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1589),
.A2(n_1085),
.B1(n_1215),
.B2(n_1676),
.Y(n_1928)
);

AOI22xp33_ASAP7_75t_L g1929 ( 
.A1(n_1589),
.A2(n_1085),
.B1(n_1215),
.B2(n_1676),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_L g1930 ( 
.A(n_1670),
.B(n_1085),
.C(n_1215),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1660),
.A2(n_1085),
.B(n_1215),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1744),
.B(n_1085),
.Y(n_1933)
);

CKINVDCx11_ASAP7_75t_R g1934 ( 
.A(n_1627),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1579),
.A2(n_1085),
.B1(n_1215),
.B2(n_1474),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1592),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1589),
.A2(n_1085),
.B1(n_841),
.B2(n_1040),
.C(n_1215),
.Y(n_1937)
);

OAI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1676),
.A2(n_1215),
.B1(n_1085),
.B2(n_664),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1578),
.A2(n_1085),
.B1(n_1215),
.B2(n_841),
.C(n_1676),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1626),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1706),
.A2(n_1085),
.B1(n_841),
.B2(n_1040),
.Y(n_1941)
);

OR2x6_ASAP7_75t_L g1942 ( 
.A(n_1725),
.B(n_1674),
.Y(n_1942)
);

AND2x6_ASAP7_75t_SL g1943 ( 
.A(n_1652),
.B(n_1466),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1837),
.B(n_1887),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1867),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1841),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1913),
.A2(n_1915),
.B1(n_1928),
.B2(n_1929),
.Y(n_1947)
);

AND2x2_ASAP7_75t_SL g1948 ( 
.A(n_1848),
.B(n_1780),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1804),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1822),
.Y(n_1950)
);

AO21x2_ASAP7_75t_L g1951 ( 
.A1(n_1862),
.A2(n_1861),
.B(n_1776),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1804),
.B(n_1851),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1933),
.B(n_1943),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1787),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1888),
.B(n_1881),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1774),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1881),
.B(n_1806),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1884),
.B(n_1802),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1824),
.Y(n_1959)
);

INVx2_ASAP7_75t_R g1960 ( 
.A(n_1886),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1788),
.B(n_1779),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1793),
.B(n_1796),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1781),
.B(n_1785),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1787),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1905),
.B(n_1907),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1923),
.Y(n_1966)
);

AOI21xp33_ASAP7_75t_L g1967 ( 
.A1(n_1924),
.A2(n_1937),
.B(n_1906),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1849),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1822),
.Y(n_1969)
);

AOI33xp33_ASAP7_75t_L g1970 ( 
.A1(n_1913),
.A2(n_1915),
.A3(n_1929),
.B1(n_1928),
.B2(n_1938),
.B3(n_1906),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1917),
.Y(n_1971)
);

NOR2xp67_ASAP7_75t_L g1972 ( 
.A(n_1864),
.B(n_1799),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1942),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1808),
.B(n_1883),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1778),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1883),
.B(n_1783),
.Y(n_1976)
);

AO21x2_ASAP7_75t_L g1977 ( 
.A1(n_1846),
.A2(n_1811),
.B(n_1812),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1810),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1833),
.B(n_1773),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1827),
.Y(n_1980)
);

AO21x2_ASAP7_75t_L g1981 ( 
.A1(n_1811),
.A2(n_1812),
.B(n_1889),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1877),
.B(n_1921),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1860),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1775),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1914),
.B(n_1878),
.Y(n_1985)
);

OAI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1813),
.A2(n_1823),
.B(n_1777),
.Y(n_1986)
);

BUFx3_ASAP7_75t_L g1987 ( 
.A(n_1908),
.Y(n_1987)
);

OAI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1916),
.A2(n_1941),
.B1(n_1909),
.B2(n_1939),
.C(n_1918),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1931),
.A2(n_1930),
.B(n_1834),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1917),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1877),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1877),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1842),
.B(n_1899),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1856),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1899),
.B(n_1800),
.Y(n_1995)
);

INVx5_ASAP7_75t_L g1996 ( 
.A(n_1917),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1803),
.B(n_1874),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1879),
.B(n_1792),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1803),
.B(n_1874),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1768),
.A2(n_1938),
.B1(n_1911),
.B2(n_1935),
.Y(n_2000)
);

INVx5_ASAP7_75t_L g2001 ( 
.A(n_1942),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1857),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1792),
.B(n_1789),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1789),
.B(n_1791),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1934),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1791),
.B(n_1780),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1840),
.Y(n_2007)
);

NOR2xp67_ASAP7_75t_L g2008 ( 
.A(n_1904),
.B(n_1818),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1873),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1922),
.B(n_1926),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1942),
.B(n_1893),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1927),
.B(n_1932),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1784),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1871),
.B(n_1772),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1936),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_1769),
.B(n_1771),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1772),
.B(n_1892),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1830),
.A2(n_1848),
.B1(n_1801),
.B2(n_1825),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1782),
.B(n_1870),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1794),
.Y(n_2020)
);

NOR4xp25_ASAP7_75t_SL g2021 ( 
.A(n_1836),
.B(n_1847),
.C(n_1863),
.D(n_1890),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1790),
.Y(n_2022)
);

AO21x2_ASAP7_75t_L g2023 ( 
.A1(n_1809),
.A2(n_1821),
.B(n_1844),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1835),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1865),
.Y(n_2025)
);

INVx4_ASAP7_75t_SL g2026 ( 
.A(n_1829),
.Y(n_2026)
);

AND2x4_ASAP7_75t_SL g2027 ( 
.A(n_1838),
.B(n_1855),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1898),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1798),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1852),
.Y(n_2030)
);

AND2x4_ASAP7_75t_SL g2031 ( 
.A(n_1838),
.B(n_1855),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1770),
.B(n_1875),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1880),
.B(n_1882),
.Y(n_2033)
);

AO21x2_ASAP7_75t_L g2034 ( 
.A1(n_1831),
.A2(n_1925),
.B(n_1826),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1886),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1886),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1875),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1782),
.B(n_1866),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1886),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1845),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1870),
.B(n_1868),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1895),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1908),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1805),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1805),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1876),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1876),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1920),
.B(n_1807),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1919),
.B(n_1829),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_1876),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1868),
.B(n_1770),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1858),
.B(n_1897),
.Y(n_2052)
);

NAND5xp2_ASAP7_75t_SL g2053 ( 
.A(n_1988),
.B(n_1830),
.C(n_1843),
.D(n_1902),
.E(n_1869),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1987),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1975),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1949),
.Y(n_2056)
);

NOR2x1p5_ASAP7_75t_L g2057 ( 
.A(n_2049),
.B(n_1814),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1965),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1963),
.B(n_1858),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1975),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1953),
.B(n_1819),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1948),
.A2(n_1829),
.B1(n_1920),
.B2(n_1940),
.Y(n_2062)
);

OAI211xp5_ASAP7_75t_L g2063 ( 
.A1(n_2000),
.A2(n_1869),
.B(n_1853),
.C(n_1885),
.Y(n_2063)
);

AOI33xp33_ASAP7_75t_L g2064 ( 
.A1(n_2030),
.A2(n_1897),
.A3(n_1900),
.B1(n_1903),
.B2(n_1815),
.B3(n_1872),
.Y(n_2064)
);

OAI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_1989),
.A2(n_1912),
.B1(n_1797),
.B2(n_1900),
.C(n_1903),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2018),
.A2(n_1829),
.B1(n_1908),
.B2(n_1816),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1963),
.B(n_1815),
.Y(n_2067)
);

AOI221xp5_ASAP7_75t_L g2068 ( 
.A1(n_1967),
.A2(n_1850),
.B1(n_1891),
.B2(n_1859),
.C(n_1828),
.Y(n_2068)
);

OAI21xp33_ASAP7_75t_L g2069 ( 
.A1(n_1970),
.A2(n_1989),
.B(n_1967),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1947),
.A2(n_1829),
.B1(n_1839),
.B2(n_1910),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1968),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1975),
.Y(n_2072)
);

AOI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_1947),
.A2(n_1795),
.B1(n_1820),
.B2(n_1786),
.C(n_1817),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1978),
.Y(n_2074)
);

OAI21x1_ASAP7_75t_L g2075 ( 
.A1(n_1950),
.A2(n_1901),
.B(n_1854),
.Y(n_2075)
);

OAI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1979),
.A2(n_1832),
.B(n_1896),
.Y(n_2076)
);

NOR2x1_ASAP7_75t_L g2077 ( 
.A(n_1979),
.B(n_1896),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1978),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1987),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1948),
.A2(n_1839),
.B1(n_1816),
.B2(n_1786),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1980),
.B(n_1876),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1961),
.B(n_1894),
.Y(n_2082)
);

AOI33xp33_ASAP7_75t_L g2083 ( 
.A1(n_2030),
.A2(n_1832),
.A3(n_1894),
.B1(n_1901),
.B2(n_2020),
.B3(n_2045),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1961),
.B(n_1894),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2024),
.B(n_2013),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_1985),
.B(n_1894),
.Y(n_2086)
);

NOR2x1_ASAP7_75t_L g2087 ( 
.A(n_2016),
.B(n_1901),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1974),
.B(n_1954),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1962),
.B(n_2002),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_SL g2090 ( 
.A1(n_2018),
.A2(n_1948),
.B1(n_2005),
.B2(n_1987),
.Y(n_2090)
);

OAI31xp33_ASAP7_75t_L g2091 ( 
.A1(n_2027),
.A2(n_2031),
.A3(n_2006),
.B(n_2032),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2021),
.A2(n_1972),
.B1(n_2032),
.B2(n_2037),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1974),
.B(n_1954),
.Y(n_2093)
);

AND2x4_ASAP7_75t_SL g2094 ( 
.A(n_2033),
.B(n_1971),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_SL g2095 ( 
.A(n_1984),
.B(n_2043),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1983),
.Y(n_2096)
);

OAI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_1972),
.A2(n_2037),
.B1(n_2014),
.B2(n_2008),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_1952),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1983),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_1965),
.Y(n_2100)
);

BUFx3_ASAP7_75t_L g2101 ( 
.A(n_2043),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1983),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1994),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1964),
.B(n_2017),
.Y(n_2104)
);

OAI33xp33_ASAP7_75t_L g2105 ( 
.A1(n_2044),
.A2(n_2045),
.A3(n_2020),
.B1(n_2014),
.B2(n_1957),
.B3(n_1955),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_1944),
.Y(n_2106)
);

AOI211xp5_ASAP7_75t_L g2107 ( 
.A1(n_2008),
.A2(n_2006),
.B(n_2052),
.C(n_2029),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1994),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1962),
.B(n_2002),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_2042),
.Y(n_2110)
);

AOI22x1_ASAP7_75t_L g2111 ( 
.A1(n_2022),
.A2(n_2052),
.B1(n_2019),
.B2(n_2051),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_2010),
.B(n_2012),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1964),
.B(n_2017),
.Y(n_2113)
);

OAI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2021),
.A2(n_2016),
.B(n_2044),
.C(n_2022),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2034),
.A2(n_2027),
.B1(n_2031),
.B2(n_2041),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2027),
.A2(n_2031),
.B1(n_2041),
.B2(n_2051),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_1957),
.B(n_1944),
.Y(n_2117)
);

OAI221xp5_ASAP7_75t_L g2118 ( 
.A1(n_2029),
.A2(n_2022),
.B1(n_2028),
.B2(n_1959),
.C(n_2025),
.Y(n_2118)
);

NAND2xp33_ASAP7_75t_R g2119 ( 
.A(n_2040),
.B(n_2033),
.Y(n_2119)
);

INVx3_ASAP7_75t_L g2120 ( 
.A(n_1949),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1976),
.B(n_1997),
.Y(n_2121)
);

INVxp67_ASAP7_75t_L g2122 ( 
.A(n_2009),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1976),
.B(n_1997),
.Y(n_2123)
);

INVxp33_ASAP7_75t_L g2124 ( 
.A(n_2010),
.Y(n_2124)
);

AO21x2_ASAP7_75t_L g2125 ( 
.A1(n_1951),
.A2(n_1981),
.B(n_1969),
.Y(n_2125)
);

NAND3xp33_ASAP7_75t_L g2126 ( 
.A(n_2028),
.B(n_2025),
.C(n_1995),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_2012),
.B(n_2043),
.Y(n_2127)
);

AOI222xp33_ASAP7_75t_L g2128 ( 
.A1(n_2004),
.A2(n_2003),
.B1(n_1999),
.B2(n_1995),
.C1(n_2019),
.C2(n_2034),
.Y(n_2128)
);

OA222x2_ASAP7_75t_L g2129 ( 
.A1(n_1998),
.A2(n_2038),
.B1(n_1958),
.B2(n_2039),
.C1(n_1968),
.C2(n_1955),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1999),
.B(n_1993),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1946),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2034),
.A2(n_2004),
.B1(n_2003),
.B2(n_1977),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1946),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_2056),
.Y(n_2134)
);

INVx5_ASAP7_75t_L g2135 ( 
.A(n_2079),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2121),
.B(n_1958),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2098),
.B(n_2040),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2055),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2055),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_2069),
.B(n_2034),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2098),
.B(n_1973),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2056),
.B(n_1952),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2088),
.B(n_1973),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2088),
.B(n_1949),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2093),
.B(n_1949),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2093),
.B(n_1949),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2121),
.B(n_1982),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_2118),
.B(n_2033),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2104),
.B(n_1949),
.Y(n_2149)
);

AND2x4_ASAP7_75t_SL g2150 ( 
.A(n_2079),
.B(n_1971),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2123),
.B(n_1982),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2123),
.B(n_1966),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2060),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2104),
.B(n_1977),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_2092),
.B(n_2033),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_2131),
.Y(n_2156)
);

AND2x4_ASAP7_75t_L g2157 ( 
.A(n_2056),
.B(n_1952),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2060),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2113),
.B(n_2129),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2117),
.B(n_1977),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2113),
.B(n_1977),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2072),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2130),
.B(n_2011),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2058),
.B(n_1966),
.Y(n_2164)
);

AND2x4_ASAP7_75t_SL g2165 ( 
.A(n_2079),
.B(n_1971),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2072),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2130),
.B(n_2011),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2074),
.Y(n_2168)
);

INVxp67_ASAP7_75t_SL g2169 ( 
.A(n_2133),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2100),
.B(n_2011),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2074),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2089),
.B(n_2109),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2059),
.B(n_2124),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_2120),
.B(n_1952),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_2120),
.B(n_2001),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2117),
.B(n_1998),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2106),
.B(n_2038),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2085),
.B(n_1992),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2122),
.B(n_1992),
.Y(n_2179)
);

BUFx2_ASAP7_75t_L g2180 ( 
.A(n_2120),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2059),
.B(n_2011),
.Y(n_2181)
);

NAND3xp33_ASAP7_75t_L g2182 ( 
.A(n_2128),
.B(n_2007),
.C(n_2015),
.Y(n_2182)
);

NAND3xp33_ASAP7_75t_L g2183 ( 
.A(n_2114),
.B(n_2007),
.C(n_2015),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2132),
.B(n_1956),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2067),
.B(n_1990),
.Y(n_2185)
);

AO21x2_ASAP7_75t_L g2186 ( 
.A1(n_2125),
.A2(n_1950),
.B(n_1969),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2082),
.B(n_1990),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2096),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_2094),
.B(n_2001),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2082),
.B(n_1990),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_2078),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2084),
.B(n_1990),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2099),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_2094),
.B(n_2001),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2084),
.B(n_1990),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2099),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2071),
.B(n_1990),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2102),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2110),
.B(n_1991),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_2177),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2138),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2159),
.B(n_2112),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_2140),
.A2(n_2090),
.B(n_2053),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2138),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2159),
.B(n_2071),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2135),
.B(n_2189),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2142),
.B(n_2054),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2140),
.A2(n_2053),
.B1(n_2111),
.B2(n_2057),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2172),
.B(n_2126),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_2182),
.B(n_2107),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2172),
.B(n_2081),
.Y(n_2211)
);

OR2x6_ASAP7_75t_L g2212 ( 
.A(n_2182),
.B(n_1971),
.Y(n_2212)
);

NOR2x1_ASAP7_75t_L g2213 ( 
.A(n_2183),
.B(n_2077),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2139),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2139),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2142),
.B(n_2054),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2160),
.B(n_2102),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2153),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2160),
.B(n_2108),
.Y(n_2219)
);

NAND2x1p5_ASAP7_75t_L g2220 ( 
.A(n_2135),
.B(n_1996),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2136),
.B(n_2086),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2136),
.B(n_2115),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2142),
.B(n_2101),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2191),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2191),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2153),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2158),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2158),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_2135),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_2142),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2157),
.B(n_2101),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_2148),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2176),
.B(n_2108),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2157),
.B(n_2127),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2186),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2162),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2162),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2166),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2186),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2176),
.B(n_2147),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2191),
.Y(n_2241)
);

INVxp67_ASAP7_75t_L g2242 ( 
.A(n_2148),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2155),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2173),
.B(n_2111),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2166),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2168),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2168),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_2135),
.B(n_1996),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2191),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2157),
.B(n_1971),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2173),
.B(n_1945),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2171),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2147),
.B(n_2103),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2157),
.B(n_1971),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2171),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2201),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2206),
.B(n_2154),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2201),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2204),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2204),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2205),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2214),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2214),
.Y(n_2263)
);

NOR3xp33_ASAP7_75t_L g2264 ( 
.A(n_2210),
.B(n_2073),
.C(n_2097),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2215),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2206),
.B(n_2154),
.Y(n_2266)
);

INVx2_ASAP7_75t_SL g2267 ( 
.A(n_2206),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2209),
.B(n_2151),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2215),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2240),
.B(n_2151),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2206),
.B(n_2161),
.Y(n_2271)
);

OR2x6_ASAP7_75t_L g2272 ( 
.A(n_2213),
.B(n_2183),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2218),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_2240),
.B(n_2184),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2250),
.B(n_2161),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2218),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2232),
.B(n_2155),
.Y(n_2277)
);

NOR3xp33_ASAP7_75t_L g2278 ( 
.A(n_2203),
.B(n_2065),
.C(n_2068),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2226),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2250),
.B(n_2185),
.Y(n_2280)
);

AND2x2_ASAP7_75t_SL g2281 ( 
.A(n_2208),
.B(n_2080),
.Y(n_2281)
);

OAI32xp33_ASAP7_75t_L g2282 ( 
.A1(n_2244),
.A2(n_2184),
.A3(n_2116),
.B1(n_2119),
.B2(n_2177),
.Y(n_2282)
);

NOR2x1_ASAP7_75t_L g2283 ( 
.A(n_2213),
.B(n_2087),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2242),
.B(n_2185),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2202),
.B(n_2152),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2222),
.B(n_2061),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2226),
.Y(n_2287)
);

NOR2xp67_ASAP7_75t_SL g2288 ( 
.A(n_2229),
.B(n_2135),
.Y(n_2288)
);

OR2x2_ASAP7_75t_L g2289 ( 
.A(n_2200),
.B(n_2178),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2224),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2205),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2202),
.B(n_2152),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2227),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2243),
.B(n_2163),
.Y(n_2294)
);

HB1xp67_ASAP7_75t_L g2295 ( 
.A(n_2212),
.Y(n_2295)
);

NOR3xp33_ASAP7_75t_L g2296 ( 
.A(n_2229),
.B(n_2063),
.C(n_2105),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2212),
.A2(n_2070),
.B1(n_2095),
.B2(n_2076),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2254),
.B(n_2174),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2227),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2228),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2221),
.B(n_2163),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2254),
.B(n_2174),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2248),
.B(n_2091),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2207),
.B(n_2174),
.Y(n_2304)
);

HB1xp67_ASAP7_75t_L g2305 ( 
.A(n_2212),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2211),
.B(n_2167),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_R g2307 ( 
.A(n_2251),
.B(n_2079),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2212),
.B(n_2167),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2212),
.B(n_2057),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2248),
.B(n_2189),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2228),
.Y(n_2311)
);

AOI222xp33_ASAP7_75t_L g2312 ( 
.A1(n_2281),
.A2(n_2248),
.B1(n_2062),
.B2(n_2181),
.C1(n_2143),
.C2(n_1986),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2280),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2264),
.B(n_2181),
.Y(n_2314)
);

AOI21xp33_ASAP7_75t_L g2315 ( 
.A1(n_2272),
.A2(n_2282),
.B(n_2309),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_2272),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2283),
.B(n_2248),
.Y(n_2317)
);

OAI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2278),
.A2(n_2220),
.B(n_2087),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2282),
.A2(n_2255),
.B1(n_2238),
.B2(n_2252),
.C(n_2237),
.Y(n_2319)
);

AOI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2281),
.A2(n_2066),
.B1(n_2023),
.B2(n_2194),
.Y(n_2320)
);

AOI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2272),
.A2(n_2023),
.B1(n_2194),
.B2(n_2189),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2272),
.A2(n_2023),
.B1(n_2194),
.B2(n_2189),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2297),
.B(n_2220),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2256),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2256),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2296),
.B(n_2234),
.Y(n_2326)
);

OAI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2303),
.A2(n_2220),
.B1(n_2230),
.B2(n_2178),
.C(n_2077),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2286),
.A2(n_2310),
.B1(n_2261),
.B2(n_2277),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2280),
.Y(n_2329)
);

OAI221xp5_ASAP7_75t_L g2330 ( 
.A1(n_2284),
.A2(n_2230),
.B1(n_2164),
.B2(n_2253),
.C(n_2233),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2258),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2258),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2274),
.B(n_2233),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2265),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2265),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2269),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2291),
.A2(n_2268),
.B1(n_2308),
.B2(n_2294),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2304),
.B(n_2207),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2269),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2273),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2273),
.Y(n_2341)
);

OAI222xp33_ASAP7_75t_L g2342 ( 
.A1(n_2288),
.A2(n_2230),
.B1(n_2135),
.B2(n_2141),
.C1(n_2231),
.C2(n_2223),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2301),
.B(n_2234),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2276),
.Y(n_2344)
);

NAND4xp25_ASAP7_75t_SL g2345 ( 
.A(n_2257),
.B(n_2064),
.C(n_2083),
.D(n_2231),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2276),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2285),
.B(n_2143),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2290),
.Y(n_2348)
);

OAI21xp33_ASAP7_75t_L g2349 ( 
.A1(n_2274),
.A2(n_1993),
.B(n_2253),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2304),
.B(n_2216),
.Y(n_2350)
);

OAI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2292),
.A2(n_2267),
.B1(n_2305),
.B2(n_2295),
.Y(n_2351)
);

AOI21xp33_ASAP7_75t_SL g2352 ( 
.A1(n_2267),
.A2(n_2075),
.B(n_2194),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2290),
.Y(n_2353)
);

AOI322xp5_ASAP7_75t_L g2354 ( 
.A1(n_2315),
.A2(n_2257),
.A3(n_2266),
.B1(n_2271),
.B2(n_2275),
.C1(n_2302),
.C2(n_2298),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2317),
.B(n_2266),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2319),
.B(n_2320),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2314),
.B(n_2275),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2313),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2341),
.Y(n_2359)
);

AOI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2316),
.A2(n_2288),
.B1(n_2271),
.B2(n_2262),
.C(n_2293),
.Y(n_2360)
);

AO21x1_ASAP7_75t_L g2361 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2259),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2326),
.B(n_2270),
.Y(n_2362)
);

AOI221x1_ASAP7_75t_L g2363 ( 
.A1(n_2351),
.A2(n_2287),
.B1(n_2279),
.B2(n_2260),
.C(n_2263),
.Y(n_2363)
);

OAI221xp5_ASAP7_75t_L g2364 ( 
.A1(n_2318),
.A2(n_2270),
.B1(n_2289),
.B2(n_2300),
.C(n_2299),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2313),
.B(n_2289),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2341),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2324),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2328),
.B(n_2306),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2338),
.B(n_2298),
.Y(n_2369)
);

AOI21xp33_ASAP7_75t_SL g2370 ( 
.A1(n_2323),
.A2(n_2075),
.B(n_2302),
.Y(n_2370)
);

INVx2_ASAP7_75t_SL g2371 ( 
.A(n_2329),
.Y(n_2371)
);

A2O1A1Ixp33_ASAP7_75t_L g2372 ( 
.A1(n_2323),
.A2(n_1986),
.B(n_2135),
.C(n_2150),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2325),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2331),
.Y(n_2374)
);

NAND2xp33_ASAP7_75t_L g2375 ( 
.A(n_2321),
.B(n_2307),
.Y(n_2375)
);

AOI31xp33_ASAP7_75t_L g2376 ( 
.A1(n_2352),
.A2(n_2223),
.A3(n_2216),
.B(n_2175),
.Y(n_2376)
);

OAI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2322),
.A2(n_2175),
.B(n_2164),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2329),
.B(n_2217),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2337),
.B(n_2170),
.Y(n_2379)
);

A2O1A1Ixp33_ASAP7_75t_L g2380 ( 
.A1(n_2327),
.A2(n_2165),
.B(n_2150),
.C(n_1996),
.Y(n_2380)
);

AOI211xp5_ASAP7_75t_L g2381 ( 
.A1(n_2342),
.A2(n_2239),
.B(n_2235),
.C(n_2175),
.Y(n_2381)
);

O2A1O1Ixp33_ASAP7_75t_L g2382 ( 
.A1(n_2312),
.A2(n_2239),
.B(n_2235),
.C(n_2023),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2332),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2338),
.B(n_2170),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2358),
.Y(n_2385)
);

OAI321xp33_ASAP7_75t_L g2386 ( 
.A1(n_2356),
.A2(n_2330),
.A3(n_2349),
.B1(n_2333),
.B2(n_2335),
.C(n_2334),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2358),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2359),
.Y(n_2388)
);

INVx4_ASAP7_75t_L g2389 ( 
.A(n_2371),
.Y(n_2389)
);

O2A1O1Ixp33_ASAP7_75t_L g2390 ( 
.A1(n_2356),
.A2(n_2339),
.B(n_2340),
.C(n_2346),
.Y(n_2390)
);

A2O1A1Ixp33_ASAP7_75t_L g2391 ( 
.A1(n_2382),
.A2(n_2370),
.B(n_2381),
.C(n_2360),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2354),
.B(n_2350),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2368),
.B(n_2362),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2366),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2357),
.B(n_2345),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2355),
.B(n_2350),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2355),
.Y(n_2397)
);

INVx1_ASAP7_75t_SL g2398 ( 
.A(n_2355),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2369),
.B(n_2343),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2365),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2367),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2373),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2379),
.B(n_2384),
.Y(n_2403)
);

OAI21xp33_ASAP7_75t_SL g2404 ( 
.A1(n_2376),
.A2(n_2333),
.B(n_2344),
.Y(n_2404)
);

NOR2xp67_ASAP7_75t_L g2405 ( 
.A(n_2364),
.B(n_2348),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2383),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2374),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2361),
.B(n_2347),
.Y(n_2408)
);

INVxp67_ASAP7_75t_L g2409 ( 
.A(n_2363),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2398),
.B(n_2380),
.Y(n_2410)
);

NOR4xp75_ASAP7_75t_L g2411 ( 
.A(n_2392),
.B(n_2377),
.C(n_2375),
.D(n_2372),
.Y(n_2411)
);

NOR4xp25_ASAP7_75t_L g2412 ( 
.A(n_2409),
.B(n_2375),
.C(n_2372),
.D(n_2380),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_SL g2413 ( 
.A(n_2409),
.B(n_2336),
.C(n_2378),
.Y(n_2413)
);

NAND5xp2_ASAP7_75t_L g2414 ( 
.A(n_2386),
.B(n_2197),
.C(n_2187),
.D(n_2190),
.E(n_2192),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_L g2415 ( 
.A(n_2391),
.B(n_2353),
.C(n_2348),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2393),
.B(n_2353),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2397),
.Y(n_2417)
);

NAND3x1_ASAP7_75t_L g2418 ( 
.A(n_2397),
.B(n_2230),
.C(n_2252),
.Y(n_2418)
);

OAI21xp33_ASAP7_75t_SL g2419 ( 
.A1(n_2408),
.A2(n_2195),
.B(n_2192),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2385),
.Y(n_2420)
);

AOI322xp5_ASAP7_75t_L g2421 ( 
.A1(n_2395),
.A2(n_2239),
.A3(n_2235),
.B1(n_2137),
.B2(n_2141),
.C1(n_2146),
.C2(n_2144),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2400),
.B(n_2187),
.Y(n_2422)
);

NOR3xp33_ASAP7_75t_SL g2423 ( 
.A(n_2402),
.B(n_2255),
.C(n_2247),
.Y(n_2423)
);

O2A1O1Ixp33_ASAP7_75t_L g2424 ( 
.A1(n_2413),
.A2(n_2390),
.B(n_2395),
.C(n_2408),
.Y(n_2424)
);

OAI221xp5_ASAP7_75t_L g2425 ( 
.A1(n_2412),
.A2(n_2404),
.B1(n_2405),
.B2(n_2393),
.C(n_2416),
.Y(n_2425)
);

NAND4xp25_ASAP7_75t_L g2426 ( 
.A(n_2414),
.B(n_2396),
.C(n_2389),
.D(n_2403),
.Y(n_2426)
);

AOI211xp5_ASAP7_75t_SL g2427 ( 
.A1(n_2413),
.A2(n_2387),
.B(n_2406),
.C(n_2401),
.Y(n_2427)
);

OAI321xp33_ASAP7_75t_L g2428 ( 
.A1(n_2415),
.A2(n_2407),
.A3(n_2399),
.B1(n_2394),
.B2(n_2388),
.C(n_2389),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2417),
.B(n_2217),
.Y(n_2429)
);

OAI211xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2423),
.A2(n_2236),
.B(n_2247),
.C(n_2246),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2422),
.B(n_2190),
.Y(n_2431)
);

AOI221xp5_ASAP7_75t_L g2432 ( 
.A1(n_2410),
.A2(n_2237),
.B1(n_2246),
.B2(n_2245),
.C(n_2238),
.Y(n_2432)
);

OAI222xp33_ASAP7_75t_L g2433 ( 
.A1(n_2411),
.A2(n_2175),
.B1(n_2197),
.B2(n_2180),
.C1(n_2219),
.C2(n_2134),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2419),
.A2(n_2150),
.B1(n_2165),
.B2(n_2079),
.Y(n_2434)
);

NOR3xp33_ASAP7_75t_L g2435 ( 
.A(n_2420),
.B(n_2423),
.C(n_2421),
.Y(n_2435)
);

AOI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2425),
.A2(n_2418),
.B(n_2195),
.C(n_2174),
.Y(n_2436)
);

AOI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2435),
.A2(n_2165),
.B1(n_2245),
.B2(n_2236),
.Y(n_2437)
);

AOI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2424),
.A2(n_2249),
.B(n_2241),
.Y(n_2438)
);

NOR3xp33_ASAP7_75t_L g2439 ( 
.A(n_2428),
.B(n_2134),
.C(n_2180),
.Y(n_2439)
);

INVx5_ASAP7_75t_L g2440 ( 
.A(n_2427),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2429),
.Y(n_2441)
);

XNOR2xp5_ASAP7_75t_L g2442 ( 
.A(n_2426),
.B(n_2048),
.Y(n_2442)
);

NAND2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2440),
.B(n_2431),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2440),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_2441),
.Y(n_2445)
);

NAND4xp25_ASAP7_75t_L g2446 ( 
.A(n_2437),
.B(n_2432),
.C(n_2434),
.D(n_2430),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2442),
.B(n_2219),
.Y(n_2447)
);

NOR2x1_ASAP7_75t_L g2448 ( 
.A(n_2438),
.B(n_2433),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2436),
.B(n_2144),
.Y(n_2449)
);

HB1xp67_ASAP7_75t_L g2450 ( 
.A(n_2439),
.Y(n_2450)
);

AOI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2445),
.A2(n_2134),
.B1(n_2137),
.B2(n_2225),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2448),
.A2(n_2224),
.B(n_2241),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2444),
.B(n_2134),
.Y(n_2453)
);

AOI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2450),
.A2(n_2249),
.B1(n_2225),
.B2(n_2149),
.Y(n_2454)
);

NAND4xp25_ASAP7_75t_L g2455 ( 
.A(n_2446),
.B(n_1968),
.C(n_2145),
.D(n_2149),
.Y(n_2455)
);

OAI321xp33_ASAP7_75t_L g2456 ( 
.A1(n_2443),
.A2(n_2444),
.A3(n_2447),
.B1(n_2449),
.B2(n_2035),
.C(n_2036),
.Y(n_2456)
);

AOI211xp5_ASAP7_75t_L g2457 ( 
.A1(n_2456),
.A2(n_2146),
.B(n_2145),
.C(n_2199),
.Y(n_2457)
);

NOR3xp33_ASAP7_75t_L g2458 ( 
.A(n_2455),
.B(n_2039),
.C(n_2047),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2454),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2453),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2460),
.B(n_2452),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2461),
.Y(n_2462)
);

HB1xp67_ASAP7_75t_L g2463 ( 
.A(n_2462),
.Y(n_2463)
);

INVxp67_ASAP7_75t_L g2464 ( 
.A(n_2462),
.Y(n_2464)
);

AO21x2_ASAP7_75t_L g2465 ( 
.A1(n_2463),
.A2(n_2459),
.B(n_2458),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2464),
.B(n_2451),
.Y(n_2466)
);

AOI222xp33_ASAP7_75t_L g2467 ( 
.A1(n_2466),
.A2(n_2457),
.B1(n_2169),
.B2(n_2196),
.C1(n_2193),
.C2(n_2188),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2465),
.A2(n_2169),
.B(n_2198),
.Y(n_2468)
);

AOI322xp5_ASAP7_75t_L g2469 ( 
.A1(n_2468),
.A2(n_2467),
.A3(n_2156),
.B1(n_2198),
.B2(n_2047),
.C1(n_2046),
.C2(n_2050),
.Y(n_2469)
);

OAI221xp5_ASAP7_75t_R g2470 ( 
.A1(n_2469),
.A2(n_1960),
.B1(n_2156),
.B2(n_2026),
.C(n_2199),
.Y(n_2470)
);

AOI211xp5_ASAP7_75t_L g2471 ( 
.A1(n_2470),
.A2(n_2179),
.B(n_2193),
.C(n_2188),
.Y(n_2471)
);


endmodule