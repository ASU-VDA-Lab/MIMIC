module real_jpeg_3343_n_23 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_23);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_23;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_47;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_0),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_1),
.B(n_48),
.C(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_2),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_5),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_6),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_7),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_9),
.B(n_73),
.C(n_78),
.Y(n_72)
);

AOI221xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_60),
.B2(n_63),
.C(n_64),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_11),
.B(n_71),
.C(n_79),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_12),
.B(n_36),
.C(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_14),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_13),
.A2(n_14),
.B(n_20),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_13),
.A2(n_41),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_69),
.C(n_80),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_17),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_20),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_53),
.C(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_57),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_55),
.B(n_56),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_51),
.B(n_54),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B(n_50),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_46),
.B(n_49),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_44),
.B(n_45),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B(n_43),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_67),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_65),
.B(n_81),
.C(n_82),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);


endmodule