module fake_jpeg_478_n_165 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx2_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_35),
.B(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_15),
.B(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_45),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx2_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_25),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_42),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_30),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_76),
.B1(n_55),
.B2(n_60),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_71),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_31),
.A2(n_21),
.B1(n_27),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_65),
.B1(n_57),
.B2(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_26),
.B1(n_27),
.B2(n_7),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_73),
.B1(n_80),
.B2(n_56),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_29),
.B(n_5),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_5),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_10),
.B(n_38),
.C(n_40),
.Y(n_80)
);

INVxp33_ASAP7_75t_SL g118 ( 
.A(n_84),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_93),
.B1(n_97),
.B2(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_68),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_81),
.C(n_77),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_85),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_71),
.B1(n_64),
.B2(n_69),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_66),
.B1(n_63),
.B2(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_104),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_68),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_53),
.Y(n_104)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_79),
.B1(n_54),
.B2(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_92),
.Y(n_132)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_94),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_86),
.B1(n_85),
.B2(n_99),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_95),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_123),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_89),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_105),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_121),
.C(n_116),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_103),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_117),
.B(n_105),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_99),
.B1(n_104),
.B2(n_91),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_107),
.B1(n_117),
.B2(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_133),
.B(n_114),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_129),
.C(n_130),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_115),
.B1(n_109),
.B2(n_106),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_141),
.B(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_149),
.C(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_148),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_126),
.B(n_133),
.C(n_124),
.D(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_154),
.C(n_153),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_141),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_146),
.B(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_126),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

OAI21x1_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_137),
.B(n_114),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_160),
.B(n_137),
.C(n_107),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_162),
.Y(n_165)
);


endmodule