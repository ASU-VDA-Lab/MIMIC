module fake_jpeg_25514_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx9p33_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_17),
.B1(n_30),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_53),
.B1(n_54),
.B2(n_26),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_39),
.B1(n_42),
.B2(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_60),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_41),
.B(n_21),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_62),
.Y(n_118)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_39),
.B1(n_41),
.B2(n_36),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_76),
.B1(n_80),
.B2(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_39),
.B1(n_42),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_28),
.B1(n_24),
.B2(n_47),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_82),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_33),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_26),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_22),
.Y(n_87)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_25),
.B(n_21),
.C(n_24),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_26),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_93),
.B1(n_56),
.B2(n_25),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_43),
.A2(n_38),
.B1(n_35),
.B2(n_24),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_57),
.C(n_52),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_112),
.C(n_35),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_30),
.B1(n_17),
.B2(n_61),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_108),
.B(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_115),
.B1(n_80),
.B2(n_72),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_47),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_38),
.C(n_35),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_76),
.B1(n_88),
.B2(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_65),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_86),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_47),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_84),
.B1(n_74),
.B2(n_66),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_144),
.B1(n_113),
.B2(n_103),
.Y(n_167)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_109),
.B1(n_108),
.B2(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_129),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_47),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_130),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_16),
.A3(n_23),
.B1(n_35),
.B2(n_38),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_133),
.B(n_134),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_28),
.B1(n_66),
.B2(n_89),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_28),
.CON(n_133),
.SN(n_133)
);

AO21x2_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_38),
.B(n_73),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_148),
.B1(n_116),
.B2(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_23),
.B(n_17),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_150),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_30),
.B1(n_61),
.B2(n_0),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_147),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_30),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_114),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_6),
.B1(n_14),
.B2(n_2),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_6),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_97),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_8),
.B(n_14),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_95),
.B(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_175),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_157),
.B(n_173),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_165),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_169),
.B1(n_181),
.B2(n_184),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_95),
.C(n_117),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_168),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_171),
.B1(n_177),
.B2(n_179),
.Y(n_202)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_116),
.B1(n_113),
.B2(n_103),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_102),
.B1(n_5),
.B2(n_2),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_102),
.B(n_1),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_5),
.C(n_13),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_10),
.B1(n_13),
.B2(n_3),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_3),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_4),
.B1(n_10),
.B2(n_12),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_152),
.B(n_148),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_15),
.B1(n_4),
.B2(n_1),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_125),
.A2(n_15),
.B1(n_4),
.B2(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_205),
.B(n_128),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_197),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_132),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_211),
.B(n_210),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_129),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_149),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_171),
.B1(n_160),
.B2(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_153),
.C(n_165),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_223),
.C(n_189),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_157),
.B(n_162),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_220),
.B(n_225),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_153),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_15),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_157),
.B(n_160),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_156),
.C(n_176),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_188),
.B(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_230),
.B(n_186),
.Y(n_236)
);

XOR2x1_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_133),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_144),
.B(n_151),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_227),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_237),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_193),
.A3(n_199),
.B1(n_191),
.B2(n_195),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_225),
.C(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_189),
.C(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_243),
.C(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_207),
.C(n_192),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_197),
.B1(n_204),
.B2(n_202),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_219),
.B1(n_221),
.B2(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_194),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_215),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_198),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_202),
.B(n_136),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_251),
.B(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_141),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_249),
.B(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_221),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_259),
.B(n_265),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_268),
.Y(n_280)
);

BUFx4f_ASAP7_75t_SL g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_243),
.C(n_242),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_278),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_247),
.B1(n_244),
.B2(n_219),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_254),
.B1(n_257),
.B2(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_254),
.C(n_253),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_261),
.C(n_265),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_284),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_261),
.B1(n_240),
.B2(n_220),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_236),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_288),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_290),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_265),
.B1(n_264),
.B2(n_256),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_234),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_272),
.B(n_275),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_288),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_286),
.B1(n_272),
.B2(n_287),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_280),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_291),
.B(n_217),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_279),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.C(n_299),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_298),
.B(n_293),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_305),
.B(n_301),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_295),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_215),
.Y(n_310)
);


endmodule