module fake_netlist_1_11300_n_689 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_689);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_689;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_30), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_34), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_76), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_57), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_65), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_75), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_48), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_42), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_12), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_63), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_28), .Y(n_93) );
OR2x2_ASAP7_75t_L g94 ( .A(n_45), .B(n_61), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_19), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_67), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_59), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_36), .Y(n_98) );
CKINVDCx14_ASAP7_75t_R g99 ( .A(n_54), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_0), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_10), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_52), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_23), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_10), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_43), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_15), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_39), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_26), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_33), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_3), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
BUFx10_ASAP7_75t_L g119 ( .A(n_5), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_6), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_46), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_24), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_35), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_12), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_103), .A2(n_38), .B(n_78), .Y(n_125) );
NOR2x1_ASAP7_75t_L g126 ( .A(n_110), .B(n_37), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
OA22x2_ASAP7_75t_SL g128 ( .A1(n_109), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_100), .B(n_1), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_103), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_102), .A2(n_2), .B1(n_4), .B2(n_6), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
OR2x2_ASAP7_75t_L g135 ( .A(n_124), .B(n_7), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_104), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_84), .B(n_44), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_115), .B(n_7), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_96), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_99), .B(n_8), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_116), .B(n_8), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_96), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_116), .A2(n_9), .B1(n_11), .B2(n_13), .Y(n_151) );
NAND2x1p5_ASAP7_75t_L g152 ( .A(n_94), .B(n_49), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_118), .B(n_9), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_97), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_98), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_105), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_91), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_120), .B(n_13), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_106), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_136), .A2(n_88), .B1(n_113), .B2(n_112), .Y(n_165) );
NOR3xp33_ASAP7_75t_L g166 ( .A(n_130), .B(n_101), .C(n_90), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_136), .B(n_99), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_132), .B(n_108), .Y(n_172) );
NOR2x1p5_ASAP7_75t_L g173 ( .A(n_135), .B(n_83), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_138), .B(n_119), .Y(n_174) );
NAND3xp33_ASAP7_75t_L g175 ( .A(n_143), .B(n_83), .C(n_86), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_132), .B(n_111), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
OR2x6_ASAP7_75t_L g178 ( .A(n_152), .B(n_107), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_138), .B(n_119), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_128), .A2(n_114), .B1(n_113), .B2(n_112), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_162), .B(n_119), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_158), .B(n_87), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_158), .B(n_87), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_158), .B(n_86), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_162), .B(n_88), .Y(n_187) );
INVxp33_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_134), .B(n_107), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_134), .B(n_50), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_155), .B(n_14), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
BUFx8_ASAP7_75t_SL g196 ( .A(n_146), .Y(n_196) );
INVxp33_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_135), .B(n_14), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_127), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_139), .B(n_15), .C(n_17), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_155), .B(n_17), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_133), .A2(n_18), .B1(n_21), .B2(n_22), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_129), .A2(n_25), .B1(n_27), .B2(n_29), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_164), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_164), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
NAND2xp33_ASAP7_75t_SL g208 ( .A(n_139), .B(n_31), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_140), .B(n_32), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_127), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_140), .B(n_40), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_157), .B(n_161), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_205), .B(n_161), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_206), .B(n_129), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_205), .B(n_157), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_167), .B(n_137), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_183), .B(n_152), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_178), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_191), .Y(n_224) );
BUFx8_ASAP7_75t_L g225 ( .A(n_174), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_184), .B(n_129), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_183), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_173), .A2(n_151), .B1(n_147), .B2(n_163), .Y(n_228) );
OAI21xp33_ASAP7_75t_SL g229 ( .A1(n_170), .A2(n_137), .B(n_131), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_178), .B(n_137), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g232 ( .A1(n_181), .A2(n_141), .B1(n_125), .B2(n_156), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_186), .B(n_142), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_178), .A2(n_131), .B1(n_142), .B2(n_156), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_165), .A2(n_125), .B1(n_126), .B2(n_156), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_169), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_169), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_182), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_185), .B(n_160), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_180), .B(n_159), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_196), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_192), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_204), .B(n_160), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_179), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_196), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_175), .B(n_160), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_183), .B(n_209), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_166), .B(n_160), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_193), .Y(n_254) );
BUFx6f_ASAP7_75t_SL g255 ( .A(n_195), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_209), .B(n_160), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_194), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_209), .B(n_159), .Y(n_260) );
AND2x6_ASAP7_75t_SL g261 ( .A(n_187), .B(n_159), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_207), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_198), .B(n_159), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_188), .B(n_159), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_211), .B(n_156), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_188), .B(n_156), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_179), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_208), .A2(n_154), .B1(n_125), .B2(n_150), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_197), .B(n_154), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_191), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_211), .B(n_154), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_189), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_197), .B(n_125), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_211), .B(n_150), .Y(n_276) );
NOR2xp67_ASAP7_75t_L g277 ( .A(n_245), .B(n_200), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_269), .A2(n_214), .B(n_172), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_232), .A2(n_181), .B1(n_176), .B2(n_208), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_275), .A2(n_212), .B(n_176), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_234), .B(n_202), .C(n_181), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_241), .A2(n_212), .B1(n_210), .B2(n_190), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_250), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_222), .A2(n_212), .B(n_207), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_225), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_224), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_222), .A2(n_177), .B(n_168), .Y(n_289) );
CKINVDCx10_ASAP7_75t_R g290 ( .A(n_255), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_225), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_231), .B(n_41), .Y(n_292) );
NOR2x1_ASAP7_75t_L g293 ( .A(n_231), .B(n_177), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_218), .B(n_203), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_221), .B(n_150), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_225), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_239), .B(n_150), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_221), .B(n_150), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_274), .A2(n_149), .B1(n_148), .B2(n_144), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_SL g300 ( .A1(n_256), .A2(n_168), .B(n_55), .C(n_56), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_271), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_252), .A2(n_149), .B(n_148), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_223), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_227), .B(n_149), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_252), .A2(n_149), .B(n_148), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g307 ( .A(n_228), .B(n_263), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_218), .B(n_47), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_227), .B(n_149), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_220), .A2(n_148), .B1(n_144), .B2(n_62), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_256), .A2(n_148), .B(n_144), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
O2A1O1Ixp5_ASAP7_75t_L g314 ( .A1(n_251), .A2(n_58), .B(n_60), .C(n_64), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_216), .A2(n_66), .B1(n_68), .B2(n_69), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g316 ( .A(n_218), .B(n_229), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_255), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_257), .B(n_79), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_221), .B(n_71), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_260), .A2(n_72), .B(n_74), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_219), .B(n_77), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_244), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_260), .A2(n_265), .B(n_272), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_258), .B(n_262), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_243), .A2(n_247), .B1(n_254), .B2(n_237), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_251), .A2(n_267), .B(n_273), .C(n_226), .Y(n_326) );
NOR2xp33_ASAP7_75t_SL g327 ( .A(n_235), .B(n_253), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_253), .Y(n_328) );
NOR3xp33_ASAP7_75t_SL g329 ( .A(n_267), .B(n_264), .C(n_233), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_244), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_217), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_326), .A2(n_269), .B(n_272), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_290), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_279), .A2(n_253), .B(n_240), .C(n_242), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_304), .B(n_261), .Y(n_337) );
AO31x2_ASAP7_75t_L g338 ( .A1(n_315), .A2(n_248), .A3(n_259), .B(n_238), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_313), .B(n_270), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_279), .A2(n_265), .B1(n_276), .B2(n_262), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_280), .A2(n_276), .B(n_262), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_324), .A2(n_262), .B(n_244), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_329), .B(n_217), .C(n_236), .Y(n_343) );
NOR2xp33_ASAP7_75t_SL g344 ( .A(n_291), .B(n_244), .Y(n_344) );
BUFx4_ASAP7_75t_R g345 ( .A(n_296), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_307), .B(n_236), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_292), .Y(n_347) );
AOI21x1_ASAP7_75t_L g348 ( .A1(n_318), .A2(n_238), .B(n_249), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_282), .A2(n_268), .B(n_249), .C(n_266), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_SL g350 ( .A1(n_318), .A2(n_266), .B(n_268), .C(n_321), .Y(n_350) );
OAI22xp5_ASAP7_75t_SL g351 ( .A1(n_286), .A2(n_284), .B1(n_294), .B2(n_281), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_294), .A2(n_292), .B1(n_327), .B2(n_316), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_325), .A2(n_309), .B(n_323), .C(n_283), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_317), .A2(n_309), .B1(n_319), .B2(n_297), .C(n_298), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_287), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_303), .A2(n_306), .A3(n_301), .B(n_288), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_324), .A2(n_285), .B(n_310), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_277), .A2(n_293), .B1(n_301), .B2(n_288), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_295), .B(n_331), .Y(n_361) );
AOI221x1_ASAP7_75t_L g362 ( .A1(n_299), .A2(n_320), .B1(n_312), .B2(n_289), .C(n_287), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_SL g363 ( .A1(n_305), .A2(n_310), .B(n_311), .C(n_330), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_287), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_287), .A2(n_302), .B1(n_283), .B2(n_305), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_300), .A2(n_314), .B1(n_302), .B2(n_322), .C(n_278), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_302), .A2(n_279), .B1(n_307), .B2(n_231), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_354), .A2(n_302), .B(n_333), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_355), .A2(n_351), .B1(n_353), .B2(n_347), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_332), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_334), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_345), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_366), .A2(n_362), .B(n_336), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_352), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_348), .A2(n_358), .B(n_341), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_360), .B(n_339), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_350), .A2(n_363), .B(n_349), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_351), .A2(n_367), .B1(n_337), .B2(n_344), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_359), .A2(n_346), .B(n_340), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_361), .A2(n_365), .B1(n_343), .B2(n_364), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_342), .A2(n_356), .B(n_364), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_338), .A2(n_357), .B(n_356), .Y(n_382) );
OA21x2_ASAP7_75t_L g383 ( .A1(n_338), .A2(n_357), .B(n_356), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_335), .A2(n_347), .B1(n_187), .B2(n_189), .Y(n_384) );
INVx4_ASAP7_75t_SL g385 ( .A(n_357), .Y(n_385) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_338), .Y(n_386) );
AO21x2_ASAP7_75t_L g387 ( .A1(n_354), .A2(n_333), .B(n_336), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_350), .A2(n_354), .B(n_363), .Y(n_388) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_337), .B(n_231), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g390 ( .A1(n_353), .A2(n_274), .B(n_279), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_332), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_332), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_332), .Y(n_394) );
AOI21x1_ASAP7_75t_L g395 ( .A1(n_348), .A2(n_362), .B(n_318), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_332), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_396), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_388), .A2(n_375), .B(n_377), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_383), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_370), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_383), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_385), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_390), .A2(n_378), .B1(n_369), .B2(n_376), .Y(n_405) );
BUFx2_ASAP7_75t_SL g406 ( .A(n_391), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_371), .B(n_396), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_394), .B(n_392), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_384), .A2(n_389), .B(n_372), .C(n_376), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_391), .Y(n_411) );
CKINVDCx6p67_ASAP7_75t_R g412 ( .A(n_386), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_394), .B(n_392), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_393), .B(n_387), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_393), .B(n_387), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
OAI21x1_ASAP7_75t_L g419 ( .A1(n_395), .A2(n_375), .B(n_368), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_395), .A2(n_387), .B(n_379), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_374), .B(n_373), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_385), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_372), .A2(n_380), .B1(n_373), .B2(n_381), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_373), .A2(n_279), .B(n_390), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_368), .A2(n_336), .B(n_354), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_386), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_414), .B(n_422), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_414), .B(n_422), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_422), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_400), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_414), .B(n_398), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_420), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_398), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_402), .B(n_417), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_420), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_424), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_402), .B(n_417), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_401), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_402), .B(n_417), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_397), .B(n_401), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_397), .B(n_416), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
INVx5_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
NOR2x1_ASAP7_75t_SL g449 ( .A(n_406), .B(n_429), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_429), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_428), .B(n_408), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_407), .B(n_416), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_429), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_408), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_404), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_409), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_428), .B(n_415), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_418), .B(n_409), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_423), .B(n_415), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_409), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_418), .B(n_413), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_423), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_430), .B(n_421), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_443), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_468), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_433), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_454), .B(n_413), .Y(n_476) );
OR2x6_ASAP7_75t_L g477 ( .A(n_438), .B(n_415), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_430), .B(n_421), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_443), .Y(n_479) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_468), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_430), .B(n_421), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_448), .B(n_415), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_451), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_455), .A2(n_405), .B1(n_415), .B2(n_412), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_451), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_454), .B(n_413), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_421), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_453), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_453), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_431), .B(n_421), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_460), .B(n_411), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_431), .B(n_427), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_432), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_434), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_446), .B(n_412), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_467), .B(n_419), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_446), .B(n_427), .Y(n_499) );
AND2x4_ASAP7_75t_SL g500 ( .A(n_436), .B(n_412), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_446), .B(n_419), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_448), .Y(n_502) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_438), .B(n_405), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_435), .B(n_419), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_435), .B(n_411), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_435), .B(n_399), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_445), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_466), .B(n_399), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_448), .B(n_399), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_469), .B(n_399), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_463), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_466), .B(n_399), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_437), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_466), .B(n_399), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_470), .B(n_426), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_425), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_439), .B(n_425), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_467), .B(n_426), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_439), .B(n_410), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_439), .B(n_410), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_477), .B(n_467), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_486), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_483), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_472), .B(n_444), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_508), .B(n_458), .Y(n_530) );
NOR2xp33_ASAP7_75t_SL g531 ( .A(n_500), .B(n_450), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_480), .B(n_463), .Y(n_532) );
BUFx3_ASAP7_75t_L g533 ( .A(n_500), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_496), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_516), .B(n_458), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_518), .B(n_440), .Y(n_536) );
AND3x2_ASAP7_75t_L g537 ( .A(n_524), .B(n_450), .C(n_440), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_512), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_483), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g540 ( .A(n_502), .B(n_448), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_518), .B(n_459), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_497), .B(n_459), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_506), .B(n_434), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_493), .B(n_442), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_475), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_493), .B(n_442), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_506), .B(n_447), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_499), .B(n_442), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_497), .B(n_447), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_499), .B(n_459), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_505), .B(n_444), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_505), .B(n_444), .Y(n_553) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_482), .A2(n_465), .B(n_436), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_477), .B(n_467), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_485), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_515), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_522), .B(n_436), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_513), .B(n_456), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_477), .B(n_467), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_513), .B(n_456), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_477), .B(n_448), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_474), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_524), .B(n_461), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_522), .B(n_465), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_472), .B(n_464), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_494), .B(n_461), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_476), .B(n_464), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_490), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_525), .B(n_452), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_494), .B(n_457), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_498), .B(n_448), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_502), .B(n_448), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_487), .B(n_457), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_490), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_525), .B(n_452), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_507), .B(n_452), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_473), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_527), .B(n_491), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_534), .B(n_491), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_529), .B(n_478), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_534), .B(n_481), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_533), .A2(n_484), .B1(n_503), .B2(n_482), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_580), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_529), .B(n_478), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_531), .A2(n_503), .B1(n_521), .B2(n_520), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_549), .B(n_507), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_538), .B(n_532), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_545), .B(n_517), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_568), .B(n_481), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_528), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_546), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_562), .B(n_498), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_539), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_556), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_568), .B(n_488), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_533), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_551), .B(n_488), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_538), .B(n_492), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g603 ( .A1(n_536), .A2(n_521), .B1(n_520), .B2(n_514), .C1(n_509), .C2(n_504), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_566), .B(n_509), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_547), .B(n_517), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_544), .B(n_495), .Y(n_607) );
NAND3xp33_ASAP7_75t_SL g608 ( .A(n_554), .B(n_482), .C(n_510), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_557), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_565), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_548), .B(n_514), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_541), .B(n_504), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_575), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_543), .A2(n_523), .B1(n_498), .B2(n_474), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_572), .B(n_501), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_540), .A2(n_510), .B(n_448), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_552), .B(n_553), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_559), .B(n_501), .Y(n_619) );
OAI32xp33_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_510), .A3(n_462), .B1(n_519), .B2(n_511), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_561), .B(n_479), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_608), .A2(n_449), .B(n_562), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_609), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_590), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_585), .A2(n_578), .B1(n_560), .B2(n_555), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_594), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_594), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_582), .B(n_570), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_613), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_583), .B(n_523), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_595), .B(n_562), .Y(n_632) );
AOI21xp33_ASAP7_75t_SL g633 ( .A1(n_590), .A2(n_564), .B(n_550), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_617), .A2(n_620), .B(n_614), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_583), .B(n_523), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_613), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_593), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_603), .B(n_567), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g639 ( .A1(n_600), .A2(n_564), .A3(n_574), .B(n_560), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_602), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_584), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_602), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_587), .B(n_579), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_596), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_586), .Y(n_645) );
NAND4xp25_ASAP7_75t_SL g646 ( .A(n_588), .B(n_576), .C(n_558), .D(n_537), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_597), .Y(n_647) );
AOI21xp33_ASAP7_75t_L g648 ( .A1(n_614), .A2(n_530), .B(n_535), .Y(n_648) );
AO21x1_ASAP7_75t_L g649 ( .A1(n_639), .A2(n_595), .B(n_621), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_633), .A2(n_581), .B(n_607), .C(n_618), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_640), .B(n_642), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_644), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_646), .A2(n_595), .B(n_574), .C(n_555), .Y(n_653) );
OAI311xp33_ASAP7_75t_L g654 ( .A1(n_626), .A2(n_615), .A3(n_519), .B1(n_605), .C1(n_591), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_625), .A2(n_615), .B1(n_589), .B2(n_611), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_632), .B(n_587), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_638), .A2(n_619), .B(n_592), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_644), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_641), .A2(n_592), .B1(n_599), .B2(n_560), .Y(n_659) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_634), .A2(n_555), .A3(n_526), .B(n_599), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_632), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_637), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_623), .A2(n_462), .B1(n_526), .B2(n_574), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_641), .A2(n_526), .B1(n_601), .B2(n_622), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_657), .A2(n_648), .B1(n_645), .B2(n_624), .C(n_647), .Y(n_665) );
AOI211x1_ASAP7_75t_SL g666 ( .A1(n_655), .A2(n_637), .B(n_630), .C(n_628), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_661), .A2(n_632), .B1(n_629), .B2(n_643), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_654), .A2(n_635), .B1(n_631), .B2(n_643), .C(n_606), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_649), .A2(n_635), .B1(n_631), .B2(n_610), .C(n_598), .Y(n_669) );
OA22x2_ASAP7_75t_L g670 ( .A1(n_659), .A2(n_537), .B1(n_604), .B2(n_616), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_651), .A2(n_653), .B1(n_663), .B2(n_664), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_653), .B(n_660), .C(n_650), .D(n_656), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_652), .B(n_658), .Y(n_673) );
NOR2x1p5_ASAP7_75t_L g674 ( .A(n_672), .B(n_662), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_671), .A2(n_629), .B1(n_636), .B2(n_627), .C(n_628), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_669), .B(n_636), .C(n_627), .Y(n_677) );
NAND3xp33_ASAP7_75t_SL g678 ( .A(n_666), .B(n_630), .C(n_604), .Y(n_678) );
BUFx3_ASAP7_75t_L g679 ( .A(n_675), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_674), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_677), .B(n_668), .Y(n_681) );
OR3x1_ASAP7_75t_L g682 ( .A(n_680), .B(n_678), .C(n_676), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_679), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_682), .A2(n_681), .B1(n_679), .B2(n_670), .Y(n_684) );
AOI22x1_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_683), .B1(n_667), .B2(n_665), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_601), .B(n_616), .C(n_612), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_569), .B1(n_462), .B2(n_511), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_573), .B1(n_557), .B2(n_612), .C(n_441), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_688), .A2(n_577), .B1(n_441), .B2(n_471), .Y(n_689) );
endmodule