module fake_jpeg_3416_n_63 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_0),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx6p67_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_9),
.B1(n_10),
.B2(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.C(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_28),
.B(n_29),
.C(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AOI211xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_30),
.B(n_28),
.C(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_39),
.B1(n_33),
.B2(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_44),
.B1(n_43),
.B2(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_16),
.B(n_10),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_53),
.B(n_22),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_47),
.C(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_56),
.B(n_52),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_22),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_22),
.B(n_20),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_60),
.Y(n_63)
);


endmodule