module fake_jpeg_416_n_202 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_80),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_76),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_70),
.B1(n_58),
.B2(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_53),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_70),
.B1(n_76),
.B2(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_76),
.B1(n_64),
.B2(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_66),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_52),
.B1(n_55),
.B2(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_72),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_72),
.B1(n_69),
.B2(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_116),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_111),
.B(n_31),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_75),
.B1(n_74),
.B2(n_65),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_75),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_28),
.Y(n_127)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_2),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_88),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_65),
.C(n_29),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_127),
.C(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_134),
.Y(n_152)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_23),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_3),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_138),
.B1(n_142),
.B2(n_9),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_103),
.B1(n_14),
.B2(n_16),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_159),
.B1(n_131),
.B2(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_162),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_24),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_25),
.Y(n_151)
);

CKINVDCx12_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_139),
.C(n_130),
.Y(n_157)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_158),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_163),
.Y(n_175)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_35),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_36),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_165),
.B(n_39),
.C(n_40),
.D(n_43),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_38),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_152),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_182),
.B(n_172),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_148),
.C(n_155),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_186),
.C(n_187),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_159),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_171),
.B1(n_168),
.B2(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_185),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_158),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_48),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_192),
.Y(n_195)
);

XOR2x1_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_176),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_182),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_179),
.B1(n_178),
.B2(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_190),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_197),
.A2(n_195),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_167),
.C(n_50),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_49),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_51),
.Y(n_202)
);


endmodule