module fake_jpeg_11297_n_290 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_55),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_52),
.Y(n_111)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_21),
.B(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_21),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_58),
.B(n_63),
.Y(n_125)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_64),
.Y(n_104)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_68),
.Y(n_108)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_2),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_76),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_81),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_4),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_25),
.B1(n_16),
.B2(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_42),
.C(n_22),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_130),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_119),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_25),
.B1(n_16),
.B2(n_23),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_95),
.A2(n_106),
.B1(n_107),
.B2(n_115),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_22),
.B1(n_39),
.B2(n_30),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_116),
.B1(n_118),
.B2(n_123),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_46),
.A2(n_23),
.B1(n_25),
.B2(n_40),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_39),
.B1(n_30),
.B2(n_29),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_26),
.B1(n_20),
.B2(n_29),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_26),
.B1(n_20),
.B2(n_6),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_65),
.A2(n_11),
.B1(n_12),
.B2(n_52),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_101),
.B(n_103),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_57),
.A2(n_11),
.B1(n_12),
.B2(n_72),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_60),
.B1(n_70),
.B2(n_67),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_132),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_80),
.B1(n_87),
.B2(n_56),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_131),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_85),
.B1(n_79),
.B2(n_87),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_94),
.B1(n_126),
.B2(n_99),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_73),
.A2(n_47),
.B1(n_49),
.B2(n_85),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_47),
.B1(n_49),
.B2(n_85),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_125),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_114),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_99),
.Y(n_142)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_89),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_131),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_151),
.B(n_90),
.Y(n_182)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

CKINVDCx9p33_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_157),
.Y(n_185)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_93),
.B(n_94),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_161),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_93),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_101),
.B(n_122),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_129),
.B1(n_90),
.B2(n_88),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_120),
.B1(n_105),
.B2(n_128),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_105),
.B1(n_120),
.B2(n_109),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_130),
.B1(n_118),
.B2(n_128),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_175),
.B1(n_183),
.B2(n_159),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_97),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_158),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_159),
.B1(n_162),
.B2(n_175),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_151),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_180),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_105),
.B1(n_120),
.B2(n_112),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_112),
.C(n_129),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_142),
.B1(n_155),
.B2(n_156),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_184),
.B(n_162),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_160),
.B1(n_163),
.B2(n_141),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_141),
.A3(n_145),
.B1(n_157),
.B2(n_137),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_136),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_159),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_149),
.B(n_154),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_149),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_208),
.B1(n_171),
.B2(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_138),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_150),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_142),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_199),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_201),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_176),
.B(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_179),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_210),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_184),
.B1(n_189),
.B2(n_169),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_180),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_168),
.C(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_219),
.C(n_205),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_205),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_224),
.A2(n_191),
.B1(n_168),
.B2(n_173),
.Y(n_241)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_219),
.C(n_212),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

AOI22x1_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_208),
.B1(n_206),
.B2(n_190),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_243),
.B1(n_244),
.B2(n_224),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_198),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_209),
.B1(n_207),
.B2(n_199),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_240),
.B1(n_241),
.B2(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_192),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_239),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_202),
.B(n_210),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_248),
.C(n_249),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_226),
.C(n_218),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_252),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_254),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_217),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_228),
.C(n_213),
.Y(n_256)
);

AO221x1_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_239),
.B1(n_228),
.B2(n_233),
.C(n_230),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_253),
.B1(n_250),
.B2(n_248),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_255),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_263),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_221),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_244),
.B(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_254),
.B(n_235),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_272),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_243),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_273),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_259),
.B1(n_260),
.B2(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_273),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_282),
.A2(n_270),
.B(n_259),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_263),
.A3(n_272),
.B1(n_281),
.B2(n_282),
.C1(n_261),
.C2(n_274),
.Y(n_286)
);

AOI31xp33_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_263),
.A3(n_274),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_223),
.Y(n_290)
);


endmodule