module fake_jpeg_29942_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_15),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_28),
.C(n_23),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_14),
.C(n_31),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_31),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_67),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_24),
.B1(n_17),
.B2(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_71),
.B1(n_14),
.B2(n_2),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_31),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_14),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_36),
.A2(n_29),
.B1(n_28),
.B2(n_16),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_47),
.B(n_29),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_81),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_31),
.Y(n_107)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_54),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_13),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_10),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_93),
.B1(n_48),
.B2(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_9),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_68),
.B(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_103),
.B1(n_51),
.B2(n_89),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_107),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_110),
.B1(n_100),
.B2(n_85),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_106),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_51),
.B1(n_55),
.B2(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_12),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_13),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_1),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_119),
.B1(n_94),
.B2(n_103),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_75),
.C(n_80),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_76),
.C(n_62),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_62),
.C(n_61),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_100),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_133),
.B(n_134),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_108),
.B(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_114),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_120),
.C(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_102),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_134),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_101),
.A3(n_95),
.B1(n_108),
.B2(n_99),
.C1(n_97),
.C2(n_94),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_135),
.A3(n_131),
.B1(n_128),
.B2(n_97),
.C1(n_123),
.C2(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_150),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_144),
.A2(n_127),
.B(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_90),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_106),
.C(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_138),
.B(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_154),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_109),
.C(n_104),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_148),
.B(n_150),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_159),
.C(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_152),
.A3(n_109),
.B1(n_87),
.B2(n_90),
.C1(n_56),
.C2(n_59),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_161),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_5),
.C(n_87),
.Y(n_164)
);


endmodule