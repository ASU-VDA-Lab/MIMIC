module fake_netlist_6_3603_n_1807 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1807);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1807;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx8_ASAP7_75t_SL g158 ( 
.A(n_107),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_40),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_53),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_6),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_5),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_93),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_54),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_7),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_21),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_90),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_48),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_119),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_82),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_58),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_44),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_18),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_88),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_65),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_5),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_20),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_43),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_49),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_30),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_72),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_68),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_66),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_8),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_28),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_86),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_73),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_59),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_124),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_95),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_128),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_31),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_40),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_139),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_157),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_39),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_74),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_67),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_137),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_8),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_27),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_11),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_87),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_24),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_104),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_45),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_76),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_127),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_113),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_30),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_120),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_81),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_35),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_43),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_57),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_55),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_62),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_126),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_50),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_112),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_24),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_70),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_34),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_37),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_20),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_55),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_46),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_152),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_49),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_17),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_56),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_60),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_11),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_141),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_94),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_150),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_18),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_47),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_34),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_156),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_46),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_109),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_147),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_33),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_41),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_48),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_2),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_14),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_54),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_35),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_101),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_121),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_130),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_22),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_98),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_89),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_99),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_186),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_199),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_197),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_199),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_203),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_203),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_160),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_221),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_221),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_213),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_213),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_223),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_223),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_190),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_230),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_262),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_295),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_230),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_219),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_234),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_234),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_235),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_226),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_180),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_189),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_219),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_242),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_224),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_162),
.Y(n_348)
);

BUFx2_ASAP7_75t_SL g349 ( 
.A(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_242),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_249),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_165),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_249),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_265),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_265),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_164),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_170),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_274),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_274),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_189),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_161),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_278),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_278),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_171),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_226),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_172),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_168),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_293),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_303),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_173),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_267),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_189),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_178),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_280),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_174),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_267),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_181),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_166),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_182),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_183),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_192),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_193),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_166),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_167),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_194),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_180),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_323),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_206),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_159),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_206),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_159),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_218),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_343),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_294),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_286),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_326),
.A2(n_240),
.B1(n_301),
.B2(n_254),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_362),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_334),
.B(n_304),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_309),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_321),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_334),
.B(n_304),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_315),
.B(n_195),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_376),
.Y(n_423)
);

BUFx12f_ASAP7_75t_L g424 ( 
.A(n_317),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_366),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_324),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_328),
.B(n_204),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_314),
.B(n_163),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_328),
.B(n_205),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_324),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_325),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_357),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_318),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_325),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_318),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_332),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_341),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_319),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_319),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_341),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_326),
.B(n_304),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_332),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_329),
.B(n_207),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_335),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_335),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_337),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_331),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_340),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_327),
.A2(n_281),
.B1(n_310),
.B2(n_208),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_451),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_L g460 ( 
.A1(n_448),
.A2(n_316),
.B1(n_327),
.B2(n_339),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

BUFx6f_ASAP7_75t_SL g462 ( 
.A(n_393),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_451),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_416),
.B(n_373),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_410),
.B(n_381),
.Y(n_467)
);

BUFx8_ASAP7_75t_SL g468 ( 
.A(n_455),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_410),
.B(n_383),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_384),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_396),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_396),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_414),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_424),
.B(n_167),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_440),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_444),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_440),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_434),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_431),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

BUFx6f_ASAP7_75t_SL g492 ( 
.A(n_393),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

BUFx6f_ASAP7_75t_SL g495 ( 
.A(n_393),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_434),
.B(n_385),
.Y(n_498)
);

BUFx8_ASAP7_75t_SL g499 ( 
.A(n_455),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_394),
.B(n_386),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_436),
.B(n_389),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_390),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_420),
.B(n_329),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_169),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_439),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_446),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_420),
.B(n_338),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_416),
.B(n_369),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_436),
.B(n_348),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_394),
.B(n_431),
.C(n_450),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_424),
.B(n_169),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_448),
.B(n_377),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_390),
.B(n_347),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_450),
.B(n_392),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_431),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_SL g530 ( 
.A1(n_392),
.A2(n_351),
.B(n_338),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

NOR2x1p5_ASAP7_75t_L g532 ( 
.A(n_391),
.B(n_351),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_433),
.Y(n_533)
);

AOI21x1_ASAP7_75t_L g534 ( 
.A1(n_408),
.A2(n_184),
.B(n_175),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_433),
.B(n_360),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_407),
.A2(n_280),
.B1(n_360),
.B2(n_286),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_395),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_402),
.B(n_352),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_408),
.B(n_184),
.C(n_175),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_409),
.A2(n_415),
.B1(n_419),
.B2(n_458),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_402),
.A2(n_370),
.B1(n_239),
.B2(n_257),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_398),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_399),
.B(n_380),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

OAI21xp33_ASAP7_75t_SL g545 ( 
.A1(n_399),
.A2(n_458),
.B(n_378),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_393),
.B(n_210),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_439),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_399),
.B(n_380),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_395),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_407),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_407),
.B(n_211),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_400),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_400),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_401),
.Y(n_557)
);

INVx4_ASAP7_75t_SL g558 ( 
.A(n_423),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_407),
.B(n_212),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_407),
.B(n_185),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_447),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_400),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_425),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_408),
.Y(n_565)
);

BUFx6f_ASAP7_75t_SL g566 ( 
.A(n_408),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_404),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_413),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_404),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_404),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_415),
.B(n_419),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_435),
.B(n_333),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_417),
.B(n_217),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_447),
.B(n_247),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_417),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_422),
.B(n_222),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_447),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_447),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_405),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_405),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_447),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_405),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_423),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_423),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_409),
.B(n_247),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_423),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_397),
.B(n_368),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_397),
.B(n_368),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_422),
.Y(n_592)
);

AND2x2_ASAP7_75t_SL g593 ( 
.A(n_397),
.B(n_189),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_429),
.B(n_228),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_429),
.A2(n_276),
.B1(n_201),
.B2(n_200),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_432),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_432),
.B(n_378),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_437),
.B(n_247),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_437),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_411),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_438),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_411),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_438),
.B(n_176),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_441),
.B(n_247),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_441),
.B(n_177),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_403),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_443),
.Y(n_607)
);

CKINVDCx6p67_ASAP7_75t_R g608 ( 
.A(n_428),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_525),
.A2(n_246),
.B(n_313),
.C(n_307),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_487),
.B(n_445),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_518),
.A2(n_246),
.B1(n_313),
.B2(n_307),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_490),
.B(n_515),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_518),
.B(n_228),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_481),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_552),
.B(n_445),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_551),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_472),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_552),
.B(n_445),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_503),
.B(n_445),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_561),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_475),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_503),
.B(n_228),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_555),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_530),
.A2(n_185),
.B(n_188),
.C(n_198),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_428),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_L g629 ( 
.A1(n_540),
.A2(n_251),
.B1(n_198),
.B2(n_202),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_557),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_488),
.A2(n_285),
.B1(n_255),
.B2(n_251),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_601),
.B(n_445),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_488),
.A2(n_188),
.B1(n_202),
.B2(n_209),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_SL g635 ( 
.A(n_540),
.B(n_428),
.C(n_187),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_593),
.B(n_228),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_475),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_561),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_463),
.Y(n_639)
);

AND2x2_ASAP7_75t_SL g640 ( 
.A(n_593),
.B(n_209),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_593),
.B(n_228),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_569),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_471),
.A2(n_214),
.B1(n_216),
.B2(n_220),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_601),
.B(n_449),
.Y(n_644)
);

NOR3xp33_ASAP7_75t_L g645 ( 
.A(n_574),
.B(n_191),
.C(n_179),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_475),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_565),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_531),
.A2(n_412),
.B(n_411),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_449),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_463),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_501),
.B(n_449),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_484),
.B(n_472),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_531),
.B(n_225),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_490),
.B(n_443),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_555),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_531),
.A2(n_418),
.B(n_412),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_533),
.B(n_452),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_510),
.B(n_452),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_590),
.B(n_435),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_476),
.Y(n_662)
);

O2A1O1Ixp5_ASAP7_75t_L g663 ( 
.A1(n_510),
.A2(n_214),
.B(n_216),
.C(n_297),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_523),
.B(n_229),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_466),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_523),
.B(n_231),
.Y(n_666)
);

AND2x6_ASAP7_75t_SL g667 ( 
.A(n_465),
.B(n_346),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_570),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_526),
.B(n_452),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_526),
.B(n_454),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_571),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_539),
.A2(n_220),
.B1(n_236),
.B2(n_241),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_466),
.B(n_232),
.Y(n_673)
);

AOI22x1_ASAP7_75t_L g674 ( 
.A1(n_560),
.A2(n_255),
.B1(n_297),
.B2(n_285),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_571),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_517),
.B(n_196),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_477),
.B(n_233),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_592),
.B(n_454),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_500),
.A2(n_277),
.B1(n_237),
.B2(n_248),
.Y(n_679)
);

INVx4_ASAP7_75t_SL g680 ( 
.A(n_475),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_477),
.B(n_264),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_484),
.B(n_453),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_591),
.B(n_453),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_557),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_592),
.B(n_504),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_578),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_539),
.A2(n_560),
.B1(n_588),
.B2(n_536),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_556),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_592),
.B(n_454),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_578),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_504),
.B(n_236),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_478),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_560),
.A2(n_243),
.B1(n_244),
.B2(n_258),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_478),
.B(n_283),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_545),
.A2(n_298),
.B1(n_287),
.B2(n_299),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_476),
.B(n_456),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_596),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_562),
.B(n_456),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_SL g699 ( 
.A(n_562),
.B(n_581),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_530),
.B(n_308),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_511),
.B(n_258),
.Y(n_701)
);

INVxp33_ASAP7_75t_L g702 ( 
.A(n_575),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_467),
.B(n_215),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g704 ( 
.A(n_545),
.B(n_245),
.C(n_227),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_511),
.B(n_259),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_535),
.B(n_259),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_596),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_565),
.B(n_311),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_535),
.B(n_263),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_591),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_599),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_599),
.B(n_263),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_607),
.B(n_266),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_607),
.B(n_266),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_490),
.B(n_270),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_565),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_SL g717 ( 
.A(n_577),
.B(n_238),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_515),
.B(n_270),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_581),
.B(n_346),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_515),
.B(n_606),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_560),
.B(n_457),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_546),
.B(n_312),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_470),
.B(n_250),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_543),
.B(n_457),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_486),
.B(n_304),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_462),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_538),
.B(n_253),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_460),
.B(n_442),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_543),
.B(n_442),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_486),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_549),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_549),
.B(n_350),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_584),
.B(n_516),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_541),
.B(n_256),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_532),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_529),
.B(n_350),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_576),
.B(n_442),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_524),
.B(n_260),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_579),
.B(n_261),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_532),
.A2(n_306),
.B1(n_269),
.B2(n_272),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_556),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_563),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_529),
.B(n_353),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_598),
.B(n_353),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_563),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_496),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_597),
.B(n_354),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_584),
.B(n_354),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_568),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_572),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_462),
.A2(n_355),
.B1(n_358),
.B2(n_359),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_SL g753 ( 
.A(n_521),
.B(n_268),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_572),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_554),
.B(n_273),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_559),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_603),
.B(n_403),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_506),
.Y(n_758)
);

INVx6_ASAP7_75t_L g759 ( 
.A(n_482),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_573),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_595),
.B(n_605),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_573),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_582),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_586),
.B(n_403),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_582),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_583),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_589),
.A2(n_426),
.B(n_418),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_604),
.B(n_355),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_583),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_459),
.B(n_403),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_585),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_608),
.B(n_358),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_462),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_608),
.B(n_359),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_585),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_459),
.B(n_403),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_469),
.A2(n_361),
.B(n_364),
.C(n_365),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_469),
.B(n_412),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_473),
.B(n_418),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_473),
.B(n_479),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_600),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_464),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_731),
.B(n_482),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_639),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_640),
.A2(n_492),
.B1(n_495),
.B2(n_566),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_730),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_649),
.B(n_479),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_652),
.B(n_461),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_616),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_616),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_746),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_743),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_639),
.Y(n_794)
);

AO22x1_ASAP7_75t_L g795 ( 
.A1(n_761),
.A2(n_547),
.B1(n_275),
.B2(n_289),
.Y(n_795)
);

AND2x2_ASAP7_75t_SL g796 ( 
.A(n_640),
.B(n_594),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_653),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_710),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_732),
.B(n_482),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_736),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_685),
.B(n_461),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_732),
.B(n_482),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_610),
.B(n_461),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_761),
.A2(n_492),
.B1(n_495),
.B2(n_566),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_647),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_676),
.B(n_494),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_676),
.B(n_494),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_682),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_772),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_651),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_R g812 ( 
.A(n_630),
.B(n_547),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_739),
.B(n_747),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_647),
.B(n_464),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_651),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_665),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_647),
.B(n_464),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_612),
.B(n_482),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_739),
.B(n_494),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_774),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_635),
.B(n_505),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_SL g822 ( 
.A(n_629),
.B(n_292),
.C(n_282),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_756),
.A2(n_492),
.B1(n_495),
.B2(n_566),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_734),
.A2(n_374),
.B(n_361),
.C(n_364),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_613),
.B(n_494),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_614),
.B(n_512),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_647),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_617),
.B(n_512),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_696),
.B(n_505),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_683),
.B(n_505),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_619),
.B(n_512),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_665),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_623),
.B(n_512),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_697),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_628),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_759),
.B(n_505),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_629),
.A2(n_284),
.B1(n_288),
.B2(n_290),
.C(n_291),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_697),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_638),
.B(n_513),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_642),
.Y(n_840)
);

BUFx8_ASAP7_75t_L g841 ( 
.A(n_620),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_650),
.B(n_513),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_660),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_734),
.B(n_505),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_782),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_668),
.B(n_513),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_671),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_675),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_751),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_751),
.Y(n_850)
);

O2A1O1Ixp5_ASAP7_75t_L g851 ( 
.A1(n_615),
.A2(n_534),
.B(n_567),
.C(n_483),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_725),
.B(n_520),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_759),
.B(n_520),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_661),
.B(n_520),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_762),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_686),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_690),
.B(n_513),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_684),
.B(n_534),
.Y(n_858)
);

AO22x1_ASAP7_75t_L g859 ( 
.A1(n_727),
.A2(n_279),
.B1(n_296),
.B2(n_305),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_782),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_704),
.B(n_520),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_782),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_752),
.B(n_464),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_612),
.B(n_520),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_707),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_765),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_655),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_711),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_765),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_716),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_622),
.B(n_655),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_703),
.A2(n_580),
.B1(n_564),
.B2(n_507),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_662),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_SL g874 ( 
.A1(n_758),
.A2(n_300),
.B1(n_302),
.B2(n_499),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_727),
.B(n_480),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_755),
.A2(n_728),
.B1(n_664),
.B2(n_666),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_744),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_721),
.Y(n_878)
);

OR2x2_ASAP7_75t_SL g879 ( 
.A(n_759),
.B(n_468),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_680),
.B(n_726),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_691),
.B(n_528),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_701),
.B(n_528),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_766),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_766),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_644),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_752),
.B(n_464),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_678),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_667),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_705),
.B(n_528),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_782),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_706),
.B(n_528),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_689),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_709),
.B(n_480),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_775),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_724),
.B(n_480),
.Y(n_895)
);

INVx8_ASAP7_75t_L g896 ( 
.A(n_719),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_687),
.B(n_474),
.Y(n_897)
);

CKINVDCx14_ASAP7_75t_R g898 ( 
.A(n_717),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_775),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_687),
.B(n_474),
.Y(n_900)
);

AND2x6_ASAP7_75t_SL g901 ( 
.A(n_703),
.B(n_365),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_637),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_624),
.B(n_474),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_755),
.B(n_480),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_624),
.B(n_474),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_726),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_637),
.B(n_474),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_773),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_646),
.B(n_483),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_781),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_728),
.A2(n_509),
.B1(n_485),
.B2(n_497),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_646),
.B(n_485),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_680),
.B(n_367),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_729),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_735),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_737),
.B(n_489),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_611),
.B(n_768),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_664),
.A2(n_497),
.B1(n_489),
.B2(n_502),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_781),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_744),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_773),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_SL g922 ( 
.A1(n_702),
.A2(n_367),
.B1(n_371),
.B2(n_372),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_611),
.B(n_542),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_723),
.B(n_371),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_741),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_636),
.A2(n_641),
.B1(n_631),
.B2(n_634),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_742),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_631),
.A2(n_634),
.B1(n_641),
.B2(n_636),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_626),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_720),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_658),
.B(n_542),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_745),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_695),
.A2(n_372),
.B1(n_374),
.B2(n_602),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_738),
.B(n_491),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_693),
.B(n_542),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_748),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_750),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_SL g938 ( 
.A1(n_723),
.A2(n_527),
.B1(n_493),
.B2(n_502),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_666),
.A2(n_677),
.B1(n_681),
.B2(n_673),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_719),
.Y(n_940)
);

CKINVDCx14_ASAP7_75t_R g941 ( 
.A(n_753),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_719),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_615),
.A2(n_602),
.B1(n_600),
.B2(n_527),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_680),
.B(n_491),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_656),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_688),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_754),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_733),
.B(n_493),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_673),
.A2(n_550),
.B1(n_519),
.B2(n_508),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_677),
.A2(n_550),
.B1(n_519),
.B2(n_508),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_749),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_760),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_763),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_659),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_769),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_693),
.B(n_542),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_771),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_738),
.B(n_553),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_700),
.B(n_553),
.Y(n_959)
);

AND2x6_ASAP7_75t_L g960 ( 
.A(n_780),
.B(n_544),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_749),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_618),
.A2(n_544),
.B(n_509),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_633),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_669),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_621),
.B(n_522),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_648),
.A2(n_522),
.B(n_427),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_779),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_749),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_672),
.A2(n_426),
.B1(n_427),
.B2(n_553),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_778),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_645),
.B(n_4),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_700),
.B(n_740),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_681),
.B(n_4),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_670),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_972),
.A2(n_694),
.B(n_627),
.C(n_698),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_813),
.A2(n_643),
.B(n_609),
.C(n_627),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_832),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_835),
.B(n_694),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_914),
.B(n_712),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_914),
.B(n_713),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_844),
.A2(n_722),
.B1(n_708),
.B2(n_654),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_832),
.Y(n_982)
);

OA22x2_ASAP7_75t_L g983 ( 
.A1(n_800),
.A2(n_692),
.B1(n_625),
.B2(n_679),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_819),
.A2(n_654),
.B(n_625),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_797),
.B(n_722),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_904),
.A2(n_567),
.B(n_764),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_810),
.B(n_715),
.Y(n_987)
);

INVx5_ASAP7_75t_L g988 ( 
.A(n_860),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_954),
.A2(n_567),
.B(n_757),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_844),
.B(n_708),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_877),
.B(n_718),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_835),
.B(n_714),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_SL g993 ( 
.A1(n_872),
.A2(n_672),
.B1(n_699),
.B2(n_609),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_786),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_803),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_880),
.B(n_776),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_803),
.Y(n_997)
);

BUFx2_ASAP7_75t_SL g998 ( 
.A(n_791),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_954),
.B(n_770),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_809),
.B(n_777),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_893),
.A2(n_657),
.B(n_553),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_806),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_884),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_798),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_972),
.A2(n_674),
.B1(n_767),
.B2(n_587),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_809),
.B(n_777),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_895),
.A2(n_587),
.B(n_548),
.Y(n_1007)
);

O2A1O1Ixp5_ASAP7_75t_SL g1008 ( 
.A1(n_948),
.A2(n_663),
.B(n_7),
.C(n_10),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_799),
.B(n_587),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_928),
.A2(n_587),
.B1(n_548),
.B2(n_514),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_921),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_928),
.A2(n_587),
.B1(n_548),
.B2(n_514),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_884),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_784),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_878),
.B(n_548),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_964),
.B(n_548),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_799),
.B(n_514),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_921),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_885),
.B(n_514),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_931),
.A2(n_514),
.B(n_558),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_917),
.B(n_558),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_794),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_974),
.B(n_558),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_812),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_973),
.A2(n_427),
.B1(n_426),
.B2(n_558),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_958),
.A2(n_146),
.B(n_136),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_958),
.A2(n_134),
.B(n_133),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_792),
.B(n_6),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_811),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_881),
.A2(n_129),
.B(n_123),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_882),
.A2(n_118),
.B(n_114),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_SL g1032 ( 
.A(n_796),
.B(n_111),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_802),
.B(n_867),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_806),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_921),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_829),
.B(n_13),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_921),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_798),
.B(n_14),
.Y(n_1038)
);

INVx3_ASAP7_75t_SL g1039 ( 
.A(n_915),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_974),
.B(n_105),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_820),
.B(n_15),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_876),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_880),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_889),
.A2(n_103),
.B(n_102),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_815),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_816),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_875),
.B(n_19),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_836),
.B(n_96),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_841),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_941),
.B(n_92),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_834),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_887),
.B(n_80),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_824),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_838),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_830),
.B(n_23),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_926),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_SL g1057 ( 
.A(n_860),
.B(n_79),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_879),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_789),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_875),
.B(n_25),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_897),
.A2(n_900),
.B(n_851),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_SL g1062 ( 
.A1(n_948),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_824),
.A2(n_31),
.B(n_32),
.C(n_36),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_812),
.Y(n_1064)
);

OR2x6_ASAP7_75t_L g1065 ( 
.A(n_836),
.B(n_853),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_840),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_SL g1067 ( 
.A1(n_821),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_796),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_939),
.A2(n_42),
.B(n_45),
.C(n_50),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_843),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_860),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_806),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_790),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_891),
.A2(n_69),
.B(n_75),
.Y(n_1074)
);

CKINVDCx14_ASAP7_75t_R g1075 ( 
.A(n_874),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_830),
.B(n_51),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_793),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_SL g1078 ( 
.A1(n_897),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_933),
.A2(n_52),
.B(n_56),
.C(n_821),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_806),
.B(n_827),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_807),
.A2(n_808),
.B(n_801),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_788),
.A2(n_871),
.B(n_959),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_920),
.B(n_852),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_861),
.A2(n_959),
.B(n_822),
.C(n_847),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_848),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_SL g1086 ( 
.A(n_888),
.B(n_922),
.C(n_837),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_873),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_827),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_856),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_827),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_787),
.A2(n_804),
.B(n_923),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_802),
.B(n_867),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_827),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_783),
.B(n_920),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_795),
.B(n_854),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_935),
.A2(n_956),
.B(n_900),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_861),
.A2(n_971),
.B1(n_933),
.B2(n_930),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_836),
.B(n_853),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_841),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_860),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_892),
.B(n_963),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_822),
.A2(n_865),
.B(n_868),
.C(n_870),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_862),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_930),
.B(n_967),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_903),
.A2(n_905),
.B(n_845),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_849),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_930),
.B(n_970),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_785),
.A2(n_853),
.B1(n_863),
.B2(n_886),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_934),
.A2(n_805),
.B(n_858),
.C(n_783),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_942),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_968),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_818),
.B(n_864),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_940),
.B(n_951),
.Y(n_1113)
);

AO21x1_ASAP7_75t_L g1114 ( 
.A1(n_916),
.A2(n_863),
.B(n_886),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_850),
.Y(n_1115)
);

BUFx4f_ASAP7_75t_L g1116 ( 
.A(n_940),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_968),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_845),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_R g1119 ( 
.A(n_941),
.B(n_898),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_930),
.A2(n_864),
.B1(n_818),
.B2(n_913),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_925),
.A2(n_936),
.B(n_932),
.C(n_927),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_SL g1122 ( 
.A1(n_898),
.A2(n_947),
.B(n_785),
.C(n_902),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_947),
.B(n_937),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_859),
.B(n_908),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_862),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_953),
.B(n_869),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_1055),
.B(n_823),
.C(n_938),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1101),
.B(n_961),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_981),
.A2(n_952),
.B(n_955),
.C(n_957),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1032),
.A2(n_961),
.B1(n_913),
.B2(n_940),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1066),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_990),
.A2(n_896),
.B(n_940),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1101),
.B(n_951),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_SL g1134 ( 
.A(n_1049),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1082),
.A2(n_916),
.B(n_817),
.Y(n_1135)
);

AO22x2_ASAP7_75t_L g1136 ( 
.A1(n_1056),
.A2(n_901),
.B1(n_924),
.B2(n_953),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1097),
.A2(n_951),
.B1(n_896),
.B2(n_890),
.Y(n_1137)
);

AOI211x1_ASAP7_75t_L g1138 ( 
.A1(n_1056),
.A2(n_944),
.B(n_842),
.C(n_825),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_980),
.B(n_951),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_SL g1140 ( 
.A1(n_975),
.A2(n_1109),
.B(n_1084),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1065),
.A2(n_890),
.B(n_862),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1070),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_1087),
.B(n_908),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1114),
.A2(n_846),
.A3(n_857),
.B(n_826),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1081),
.A2(n_814),
.B(n_817),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_980),
.B(n_979),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1076),
.B(n_949),
.C(n_950),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_992),
.B(n_896),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_976),
.A2(n_906),
.B(n_902),
.C(n_918),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1096),
.A2(n_911),
.B(n_965),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1047),
.A2(n_828),
.B(n_831),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1083),
.B(n_906),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1001),
.A2(n_962),
.B(n_966),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1102),
.A2(n_945),
.B(n_839),
.C(n_833),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1036),
.B(n_945),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1108),
.A2(n_894),
.A3(n_910),
.B(n_899),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1085),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1089),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_R g1159 ( 
.A(n_1119),
.B(n_919),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1060),
.A2(n_862),
.B1(n_890),
.B2(n_943),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_978),
.B(n_1104),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_989),
.A2(n_944),
.B(n_907),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1108),
.A2(n_1010),
.A3(n_1012),
.B(n_986),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_999),
.A2(n_907),
.B(n_909),
.Y(n_1164)
);

AO32x2_ASAP7_75t_L g1165 ( 
.A1(n_1068),
.A2(n_960),
.A3(n_943),
.B1(n_866),
.B2(n_883),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1007),
.A2(n_909),
.B(n_912),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1024),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_1018),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1104),
.B(n_1107),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1039),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1086),
.B(n_929),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1079),
.B(n_929),
.C(n_946),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1105),
.A2(n_855),
.B(n_946),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1067),
.B(n_969),
.C(n_960),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_994),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_984),
.A2(n_960),
.B(n_969),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1061),
.A2(n_960),
.B(n_1010),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1120),
.A2(n_960),
.B1(n_1118),
.B2(n_1098),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1011),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_994),
.B(n_1004),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1110),
.B(n_1094),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1014),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1022),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1011),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1061),
.A2(n_1012),
.B(n_1020),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1005),
.A2(n_1040),
.B(n_1021),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_SL g1187 ( 
.A(n_1095),
.B(n_1032),
.C(n_1069),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1008),
.A2(n_983),
.B(n_1040),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1029),
.Y(n_1189)
);

INVxp67_ASAP7_75t_SL g1190 ( 
.A(n_1018),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_987),
.B(n_1116),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1052),
.A2(n_1016),
.B(n_1026),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1052),
.A2(n_1016),
.B(n_1027),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1000),
.B(n_1006),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1068),
.A2(n_1053),
.B(n_1063),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1126),
.A2(n_1015),
.B(n_1019),
.Y(n_1196)
);

AOI221x1_ASAP7_75t_L g1197 ( 
.A1(n_1042),
.A2(n_993),
.B1(n_1030),
.B2(n_1074),
.C(n_1031),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1124),
.B(n_1123),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1018),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1065),
.A2(n_1098),
.B1(n_1048),
.B2(n_1064),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1117),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_995),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1045),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_983),
.A2(n_1062),
.B(n_1015),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1122),
.A2(n_985),
.B(n_1121),
.Y(n_1205)
);

NAND3x1_ASAP7_75t_L g1206 ( 
.A(n_1038),
.B(n_1028),
.C(n_1041),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1112),
.B(n_1126),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1035),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1019),
.A2(n_1023),
.A3(n_1057),
.B(n_977),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_1113),
.A2(n_1044),
.B(n_991),
.C(n_1009),
.Y(n_1210)
);

NAND3x1_ASAP7_75t_L g1211 ( 
.A(n_1075),
.B(n_1058),
.C(n_1050),
.Y(n_1211)
);

AO32x2_ASAP7_75t_L g1212 ( 
.A1(n_1093),
.A2(n_1100),
.A3(n_1078),
.B1(n_1098),
.B2(n_1065),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_988),
.A2(n_1017),
.B(n_1033),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1112),
.B(n_1054),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1046),
.B(n_1051),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1092),
.B(n_982),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_997),
.A2(n_1003),
.B(n_1013),
.C(n_1059),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1111),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1080),
.A2(n_1034),
.B(n_1088),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_998),
.B(n_1048),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_988),
.A2(n_1025),
.B(n_1048),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1035),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_SL g1223 ( 
.A1(n_1093),
.A2(n_1100),
.B(n_1106),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1099),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1035),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1116),
.B(n_1073),
.Y(n_1226)
);

INVx3_ASAP7_75t_SL g1227 ( 
.A(n_1043),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1080),
.A2(n_1072),
.B(n_1088),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1077),
.A2(n_1115),
.A3(n_996),
.B(n_1002),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_996),
.A2(n_1002),
.A3(n_1034),
.B(n_1090),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1043),
.B(n_1072),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1043),
.B(n_1037),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1037),
.A2(n_1071),
.B(n_1103),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1090),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_988),
.A2(n_1037),
.B(n_1071),
.Y(n_1235)
);

CKINVDCx12_ASAP7_75t_R g1236 ( 
.A(n_988),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1071),
.B(n_1103),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1103),
.B(n_1125),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1125),
.B(n_996),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1125),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_996),
.A2(n_962),
.B(n_966),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1096),
.A2(n_1082),
.B(n_1061),
.Y(n_1242)
);

O2A1O1Ixp5_ASAP7_75t_L g1243 ( 
.A1(n_1047),
.A2(n_844),
.B(n_1060),
.C(n_990),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_981),
.A2(n_761),
.B(n_844),
.C(n_972),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1066),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1066),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1001),
.A2(n_962),
.B(n_966),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_994),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1066),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1096),
.A2(n_1082),
.B(n_1061),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1096),
.A2(n_1082),
.B(n_1061),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1096),
.A2(n_1082),
.B(n_1061),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_1122),
.A2(n_1084),
.B(n_975),
.C(n_990),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_981),
.A2(n_761),
.B(n_844),
.C(n_972),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1101),
.B(n_525),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1083),
.B(n_696),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1101),
.B(n_525),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1083),
.B(n_696),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_994),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1083),
.B(n_696),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_994),
.B(n_314),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1065),
.B(n_1098),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1066),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1083),
.B(n_696),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1004),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1082),
.A2(n_1081),
.B(n_1091),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_1118),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1082),
.A2(n_1081),
.B(n_1091),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1114),
.A2(n_975),
.A3(n_1084),
.B(n_1108),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_994),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1004),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_SL g1272 ( 
.A1(n_1056),
.A2(n_990),
.B(n_1068),
.C(n_615),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1082),
.A2(n_1081),
.B(n_1091),
.Y(n_1273)
);

AOI31xp67_ASAP7_75t_L g1274 ( 
.A1(n_981),
.A2(n_990),
.A3(n_983),
.B(n_876),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1180),
.B(n_1146),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1256),
.B(n_1258),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1202),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1131),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1161),
.B(n_1260),
.Y(n_1280)
);

AO32x2_ASAP7_75t_L g1281 ( 
.A1(n_1137),
.A2(n_1178),
.A3(n_1160),
.B1(n_1165),
.B2(n_1274),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1224),
.A2(n_1261),
.B1(n_1148),
.B2(n_1262),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1179),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1264),
.B(n_1194),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_SL g1285 ( 
.A(n_1184),
.B(n_1170),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1273),
.A2(n_1254),
.B(n_1244),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1142),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1230),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1157),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1158),
.Y(n_1290)
);

AOI221xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1171),
.A2(n_1200),
.B1(n_1198),
.B2(n_1137),
.C(n_1205),
.Y(n_1291)
);

BUFx5_ASAP7_75t_L g1292 ( 
.A(n_1234),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1245),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1246),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1249),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1263),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1230),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1130),
.A2(n_1187),
.B1(n_1195),
.B2(n_1128),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_SL g1299 ( 
.A1(n_1174),
.A2(n_1195),
.B(n_1149),
.C(n_1188),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_SL g1300 ( 
.A1(n_1221),
.A2(n_1130),
.B(n_1204),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_1136),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1135),
.A2(n_1162),
.B(n_1166),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1248),
.B(n_1259),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1182),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1215),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1183),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1248),
.B(n_1259),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1127),
.A2(n_1136),
.B1(n_1262),
.B2(n_1147),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1145),
.A2(n_1173),
.B(n_1176),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1133),
.B(n_1139),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1179),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1197),
.A2(n_1186),
.A3(n_1193),
.B(n_1192),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1242),
.A2(n_1251),
.B(n_1250),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1155),
.B(n_1262),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1189),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1242),
.A2(n_1252),
.B(n_1250),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1231),
.B(n_1207),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1203),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1179),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1267),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1156),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1175),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1150),
.A2(n_1196),
.B(n_1164),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1150),
.A2(n_1272),
.B(n_1210),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1237),
.B(n_1220),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1239),
.A2(n_1188),
.B(n_1160),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1204),
.A2(n_1243),
.B(n_1219),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1216),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1228),
.A2(n_1213),
.B(n_1172),
.Y(n_1330)
);

OAI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1127),
.A2(n_1147),
.B1(n_1132),
.B2(n_1181),
.C(n_1152),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1230),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1156),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1270),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1206),
.A2(n_1154),
.B(n_1129),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1214),
.Y(n_1336)
);

AOI221xp5_ASAP7_75t_L g1337 ( 
.A1(n_1253),
.A2(n_1151),
.B1(n_1138),
.B2(n_1265),
.C(n_1271),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1217),
.A2(n_1233),
.B(n_1235),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1201),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1223),
.A2(n_1191),
.B(n_1163),
.Y(n_1340)
);

NOR2xp67_ASAP7_75t_L g1341 ( 
.A(n_1167),
.B(n_1184),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1199),
.A2(n_1232),
.B(n_1226),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1199),
.A2(n_1238),
.B(n_1229),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1229),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1190),
.A2(n_1163),
.B(n_1144),
.Y(n_1345)
);

AOI221xp5_ASAP7_75t_L g1346 ( 
.A1(n_1218),
.A2(n_1134),
.B1(n_1227),
.B2(n_1269),
.C(n_1240),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1163),
.A2(n_1144),
.B(n_1269),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1144),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1209),
.A2(n_1212),
.B(n_1143),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1236),
.A2(n_1211),
.B1(n_1225),
.B2(n_1168),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1225),
.B(n_1208),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1168),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1208),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1212),
.A2(n_1165),
.B(n_1209),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1159),
.B(n_1222),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1209),
.A2(n_1212),
.B(n_1165),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1222),
.B(n_1168),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1222),
.B(n_1134),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1175),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1187),
.A2(n_844),
.B1(n_574),
.B2(n_761),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1131),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1185),
.A2(n_1273),
.B(n_1268),
.Y(n_1364)
);

AO32x2_ASAP7_75t_L g1365 ( 
.A1(n_1137),
.A2(n_1056),
.A3(n_1068),
.B1(n_1108),
.B2(n_993),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_844),
.C(n_1032),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1175),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1202),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_844),
.C(n_1032),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1266),
.A2(n_1273),
.B(n_1268),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1167),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1169),
.B(n_1161),
.Y(n_1376)
);

OAI222xp33_ASAP7_75t_L g1377 ( 
.A1(n_1130),
.A2(n_1067),
.B1(n_540),
.B2(n_1068),
.C1(n_1056),
.C2(n_410),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1131),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1224),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1266),
.A2(n_1273),
.B(n_1268),
.Y(n_1381)
);

OR2x6_ASAP7_75t_L g1382 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1131),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1206),
.A2(n_844),
.B1(n_439),
.B2(n_507),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1202),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_844),
.C(n_1032),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_465),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_465),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1255),
.A2(n_540),
.B1(n_1032),
.B2(n_419),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1168),
.B(n_1011),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1131),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1202),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1244),
.A2(n_1254),
.A3(n_1177),
.B(n_1185),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1202),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_844),
.C(n_1032),
.Y(n_1397)
);

AOI22x1_ASAP7_75t_L g1398 ( 
.A1(n_1136),
.A2(n_1193),
.B1(n_1192),
.B2(n_1027),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1168),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1175),
.Y(n_1400)
);

OAI22x1_ASAP7_75t_L g1401 ( 
.A1(n_1127),
.A2(n_844),
.B1(n_540),
.B2(n_574),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1175),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1175),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1202),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_465),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1175),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1153),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_844),
.C(n_574),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1360),
.A2(n_1385),
.B1(n_1308),
.B2(n_1397),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_R g1410 ( 
.A(n_1355),
.B(n_1285),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1376),
.B(n_1310),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1376),
.B(n_1310),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1279),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_L g1414 ( 
.A(n_1280),
.B(n_1275),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1276),
.B(n_1317),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1278),
.B(n_1361),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1380),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1317),
.B(n_1326),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1389),
.A2(n_1405),
.B(n_1390),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1290),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1284),
.B(n_1359),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1367),
.A2(n_1397),
.B1(n_1370),
.B2(n_1387),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1377),
.A2(n_1391),
.B(n_1367),
.C(n_1387),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1370),
.A2(n_1408),
.B(n_1335),
.C(n_1298),
.Y(n_1424)
);

O2A1O1Ixp5_ASAP7_75t_L g1425 ( 
.A1(n_1286),
.A2(n_1316),
.B(n_1374),
.C(n_1381),
.Y(n_1425)
);

NOR2xp67_ASAP7_75t_L g1426 ( 
.A(n_1368),
.B(n_1400),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1322),
.A2(n_1382),
.B1(n_1373),
.B2(n_1372),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1290),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1325),
.A2(n_1356),
.B(n_1324),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1291),
.A2(n_1337),
.B(n_1331),
.C(n_1365),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1322),
.A2(n_1382),
.B1(n_1282),
.B2(n_1305),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1296),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1299),
.A2(n_1402),
.B(n_1339),
.C(n_1300),
.Y(n_1433)
);

OAI31xp33_ASAP7_75t_L g1434 ( 
.A1(n_1355),
.A2(n_1299),
.A3(n_1336),
.B(n_1323),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1322),
.A2(n_1382),
.B(n_1364),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1304),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1317),
.B(n_1301),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1326),
.B(n_1314),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1325),
.A2(n_1356),
.B(n_1324),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1306),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1322),
.A2(n_1382),
.B(n_1364),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1306),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1283),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1329),
.B(n_1303),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1303),
.A2(n_1307),
.B1(n_1346),
.B2(n_1320),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1315),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1307),
.A2(n_1334),
.B(n_1403),
.C(n_1406),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1401),
.B(n_1277),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1401),
.B(n_1277),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1287),
.A2(n_1383),
.B(n_1318),
.C(n_1378),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1369),
.B(n_1386),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1392),
.A2(n_1352),
.B(n_1341),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1326),
.B(n_1358),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1350),
.A2(n_1293),
.B1(n_1294),
.B2(n_1362),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1289),
.A2(n_1393),
.B(n_1295),
.C(n_1338),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1394),
.B(n_1396),
.Y(n_1456)
);

OAI22x1_ASAP7_75t_L g1457 ( 
.A1(n_1398),
.A2(n_1315),
.B1(n_1297),
.B2(n_1332),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1311),
.B(n_1375),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1380),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1395),
.B(n_1342),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1394),
.B(n_1404),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1309),
.A2(n_1347),
.B(n_1302),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1375),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1396),
.B(n_1404),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1392),
.A2(n_1353),
.B(n_1340),
.C(n_1399),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1395),
.B(n_1342),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1351),
.B(n_1357),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1340),
.A2(n_1399),
.B(n_1333),
.C(n_1321),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1311),
.A2(n_1319),
.B1(n_1283),
.B2(n_1352),
.Y(n_1469)
);

O2A1O1Ixp5_ASAP7_75t_L g1470 ( 
.A1(n_1321),
.A2(n_1333),
.B(n_1348),
.C(n_1297),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1351),
.B(n_1357),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1348),
.A2(n_1313),
.B(n_1332),
.C(n_1297),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1309),
.A2(n_1347),
.B(n_1302),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1313),
.A2(n_1288),
.B(n_1332),
.C(n_1344),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1288),
.A2(n_1365),
.B(n_1354),
.C(n_1395),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1288),
.A2(n_1365),
.B(n_1354),
.C(n_1395),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1327),
.B(n_1343),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1365),
.A2(n_1312),
.B(n_1281),
.C(n_1330),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1319),
.B(n_1352),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1281),
.A2(n_1312),
.B1(n_1327),
.B2(n_1328),
.C(n_1345),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1343),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1345),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1281),
.A2(n_1292),
.B1(n_1312),
.B2(n_1328),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1349),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1349),
.A2(n_1281),
.B(n_1312),
.C(n_1366),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_L g1486 ( 
.A(n_1292),
.B(n_1363),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1371),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1379),
.A2(n_1384),
.B(n_1388),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1407),
.B(n_1276),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1407),
.B(n_1326),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1326),
.B(n_1262),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1276),
.B(n_1317),
.Y(n_1492)
);

INVx11_ASAP7_75t_L g1493 ( 
.A(n_1375),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1374),
.A2(n_1244),
.B(n_1254),
.Y(n_1494)
);

O2A1O1Ixp5_ASAP7_75t_L g1495 ( 
.A1(n_1389),
.A2(n_1405),
.B(n_1390),
.C(n_1335),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1376),
.B(n_1310),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1325),
.A2(n_1381),
.B(n_1374),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1279),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1279),
.Y(n_1499)
);

BUFx8_ASAP7_75t_SL g1500 ( 
.A(n_1375),
.Y(n_1500)
);

NAND3xp33_ASAP7_75t_L g1501 ( 
.A(n_1495),
.B(n_1424),
.C(n_1409),
.Y(n_1501)
);

AOI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_1495),
.B2(n_1422),
.C(n_1430),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1490),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1460),
.B(n_1466),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1481),
.B(n_1486),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1484),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1489),
.B(n_1477),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1488),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1434),
.A2(n_1427),
.B1(n_1494),
.B2(n_1414),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1485),
.B(n_1429),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1485),
.A2(n_1480),
.B(n_1425),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1430),
.A2(n_1425),
.B(n_1435),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1483),
.B(n_1429),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1441),
.A2(n_1433),
.B(n_1445),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1429),
.B(n_1439),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1439),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1448),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1410),
.B(n_1431),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1421),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1439),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1449),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1437),
.B(n_1487),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1487),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1410),
.A2(n_1454),
.B1(n_1411),
.B2(n_1412),
.Y(n_1525)
);

OAI21xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1496),
.A2(n_1436),
.B(n_1442),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1472),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1482),
.B(n_1462),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1413),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1491),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1482),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1420),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1428),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1470),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1457),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1470),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1440),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1437),
.B(n_1475),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1444),
.B(n_1498),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1476),
.B(n_1497),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1432),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1462),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1468),
.B(n_1465),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1446),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1473),
.B(n_1499),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1450),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1416),
.B(n_1461),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1418),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1517),
.B(n_1521),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1545),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1531),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1545),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1545),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1506),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1517),
.B(n_1447),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1521),
.B(n_1426),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1505),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1501),
.A2(n_1492),
.B1(n_1415),
.B2(n_1453),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1504),
.B(n_1464),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1504),
.B(n_1456),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1505),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1519),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1507),
.B(n_1438),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1501),
.A2(n_1455),
.B1(n_1459),
.B2(n_1417),
.C(n_1451),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1502),
.A2(n_1463),
.B1(n_1500),
.B2(n_1467),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1537),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1507),
.B(n_1471),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1529),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1546),
.B(n_1519),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1510),
.B(n_1443),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1521),
.B(n_1443),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1537),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1523),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1570),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1569),
.B(n_1503),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1549),
.B(n_1523),
.Y(n_1579)
);

AOI211xp5_ASAP7_75t_L g1580 ( 
.A1(n_1566),
.A2(n_1502),
.B(n_1514),
.C(n_1512),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1570),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1571),
.B(n_1564),
.Y(n_1583)
);

OAI322xp33_ASAP7_75t_L g1584 ( 
.A1(n_1556),
.A2(n_1546),
.A3(n_1547),
.B1(n_1539),
.B2(n_1513),
.C1(n_1538),
.C2(n_1518),
.Y(n_1584)
);

OAI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1556),
.A2(n_1525),
.B(n_1509),
.Y(n_1585)
);

OAI321xp33_ASAP7_75t_L g1586 ( 
.A1(n_1557),
.A2(n_1509),
.A3(n_1543),
.B1(n_1527),
.B2(n_1513),
.C(n_1540),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1558),
.B(n_1543),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1575),
.B(n_1564),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1555),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1558),
.B(n_1543),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1567),
.A2(n_1559),
.B1(n_1557),
.B2(n_1571),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1551),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1567),
.A2(n_1543),
.B1(n_1527),
.B2(n_1513),
.C(n_1526),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1559),
.A2(n_1526),
.B1(n_1510),
.B2(n_1535),
.C(n_1539),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1562),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1543),
.Y(n_1598)
);

AOI33xp33_ASAP7_75t_L g1599 ( 
.A1(n_1568),
.A2(n_1510),
.A3(n_1540),
.B1(n_1532),
.B2(n_1533),
.B3(n_1515),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1572),
.A2(n_1522),
.B1(n_1530),
.B2(n_1543),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1555),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1568),
.A2(n_1535),
.B1(n_1547),
.B2(n_1574),
.C(n_1540),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1569),
.B(n_1572),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1574),
.A2(n_1548),
.B1(n_1533),
.B2(n_1532),
.C(n_1544),
.Y(n_1604)
);

OAI332xp33_ASAP7_75t_L g1605 ( 
.A1(n_1575),
.A2(n_1524),
.A3(n_1534),
.B1(n_1536),
.B2(n_1528),
.B3(n_1542),
.C1(n_1541),
.C2(n_1544),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1572),
.A2(n_1522),
.B1(n_1530),
.B2(n_1548),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1562),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1550),
.B(n_1503),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1560),
.B(n_1522),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1565),
.A2(n_1511),
.B1(n_1527),
.B2(n_1530),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1588),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1587),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1582),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1593),
.B(n_1552),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1603),
.B(n_1552),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1608),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1581),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1587),
.B(n_1558),
.Y(n_1623)
);

OAI21xp33_ASAP7_75t_L g1624 ( 
.A1(n_1585),
.A2(n_1527),
.B(n_1561),
.Y(n_1624)
);

INVx4_ASAP7_75t_SL g1625 ( 
.A(n_1587),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1589),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1576),
.Y(n_1627)
);

NOR2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1583),
.B(n_1558),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1589),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1586),
.A2(n_1520),
.B(n_1516),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1584),
.A2(n_1527),
.B(n_1511),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1590),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1590),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1578),
.B(n_1553),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1588),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1592),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_L g1641 ( 
.A(n_1631),
.B(n_1628),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1633),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1621),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1615),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1614),
.B(n_1598),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1621),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1622),
.Y(n_1648)
);

NAND4xp25_ASAP7_75t_L g1649 ( 
.A(n_1624),
.B(n_1580),
.C(n_1596),
.D(n_1595),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1614),
.B(n_1598),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1636),
.B(n_1598),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1615),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_SL g1654 ( 
.A(n_1613),
.B(n_1591),
.C(n_1599),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1620),
.B(n_1500),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1636),
.B(n_1623),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1618),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1622),
.Y(n_1658)
);

OAI21xp33_ASAP7_75t_L g1659 ( 
.A1(n_1613),
.A2(n_1599),
.B(n_1602),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1630),
.A2(n_1600),
.B1(n_1606),
.B2(n_1604),
.C(n_1527),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1563),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1625),
.B(n_1563),
.Y(n_1663)
);

AND2x4_ASAP7_75t_SL g1664 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1616),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1607),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1605),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1625),
.B(n_1609),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1627),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1620),
.B(n_1463),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1628),
.Y(n_1671)
);

NOR2xp67_ASAP7_75t_L g1672 ( 
.A(n_1620),
.B(n_1609),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1640),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1658),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1658),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_L g1677 ( 
.A1(n_1649),
.A2(n_1634),
.B(n_1633),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1642),
.Y(n_1678)
);

OAI31xp33_ASAP7_75t_L g1679 ( 
.A1(n_1649),
.A2(n_1633),
.A3(n_1634),
.B(n_1640),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1644),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1672),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1647),
.B(n_1617),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1493),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1641),
.B(n_1625),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1644),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1659),
.B(n_1630),
.C(n_1634),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1617),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1642),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1642),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1653),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1670),
.B(n_1619),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1653),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1654),
.B(n_1612),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1641),
.B(n_1625),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1612),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1665),
.Y(n_1700)
);

INVxp67_ASAP7_75t_SL g1701 ( 
.A(n_1672),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1651),
.A2(n_1630),
.B(n_1638),
.Y(n_1702)
);

NOR5xp2_ASAP7_75t_L g1703 ( 
.A(n_1661),
.B(n_1626),
.C(n_1635),
.D(n_1632),
.E(n_1629),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1665),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1671),
.B(n_1625),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1670),
.B(n_1619),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1648),
.B(n_1638),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1671),
.B(n_1619),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1674),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1675),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1698),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1685),
.B(n_1673),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1707),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1682),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1687),
.B(n_1656),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1677),
.A2(n_1654),
.B1(n_1661),
.B2(n_1668),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1691),
.Y(n_1718)
);

AOI222xp33_ASAP7_75t_L g1719 ( 
.A1(n_1681),
.A2(n_1673),
.B1(n_1648),
.B2(n_1655),
.C1(n_1668),
.C2(n_1666),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1692),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1676),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1680),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1656),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1688),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1697),
.B(n_1643),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1705),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1707),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1698),
.B(n_1656),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1693),
.Y(n_1729)
);

CKINVDCx16_ASAP7_75t_R g1730 ( 
.A(n_1686),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1707),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1696),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1705),
.B(n_1664),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1699),
.B(n_1643),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1726),
.B(n_1689),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_1720),
.Y(n_1736)
);

BUFx12f_ASAP7_75t_L g1737 ( 
.A(n_1726),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1716),
.A2(n_1679),
.B(n_1719),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1726),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1719),
.A2(n_1702),
.B(n_1686),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1726),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1733),
.A2(n_1701),
.B1(n_1630),
.B2(n_1694),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1717),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1733),
.B(n_1708),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1712),
.A2(n_1630),
.B1(n_1706),
.B2(n_1703),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1713),
.B(n_1708),
.Y(n_1746)
);

AOI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1718),
.A2(n_1709),
.B1(n_1704),
.B2(n_1700),
.C1(n_1664),
.C2(n_1646),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1713),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1720),
.A2(n_1643),
.B(n_1646),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1730),
.A2(n_1645),
.B1(n_1652),
.B2(n_1650),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1712),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1728),
.Y(n_1752)
);

AOI321xp33_ASAP7_75t_L g1753 ( 
.A1(n_1710),
.A2(n_1646),
.A3(n_1650),
.B1(n_1645),
.B2(n_1652),
.C(n_1699),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1736),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1752),
.B(n_1711),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1738),
.B(n_1714),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1743),
.B(n_1725),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1748),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1746),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1746),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1739),
.B(n_1711),
.Y(n_1761)
);

INVxp33_ASAP7_75t_L g1762 ( 
.A(n_1735),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1740),
.A2(n_1730),
.B1(n_1744),
.B2(n_1715),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1741),
.Y(n_1764)
);

AO21x1_ASAP7_75t_L g1765 ( 
.A1(n_1762),
.A2(n_1740),
.B(n_1745),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1762),
.A2(n_1749),
.B(n_1747),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1756),
.A2(n_1728),
.B1(n_1750),
.B2(n_1737),
.Y(n_1767)
);

OAI21xp33_ASAP7_75t_L g1768 ( 
.A1(n_1763),
.A2(n_1751),
.B(n_1747),
.Y(n_1768)
);

NOR4xp25_ASAP7_75t_L g1769 ( 
.A(n_1759),
.B(n_1753),
.C(n_1749),
.D(n_1721),
.Y(n_1769)
);

AOI21xp33_ASAP7_75t_L g1770 ( 
.A1(n_1754),
.A2(n_1725),
.B(n_1713),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1758),
.A2(n_1742),
.B1(n_1760),
.B2(n_1755),
.Y(n_1771)
);

OAI21xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1755),
.A2(n_1753),
.B(n_1731),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1761),
.A2(n_1710),
.B(n_1721),
.Y(n_1773)
);

AOI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1757),
.A2(n_1731),
.B(n_1727),
.C(n_1722),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1769),
.B(n_1766),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1774),
.Y(n_1776)
);

NOR2x1_ASAP7_75t_SL g1777 ( 
.A(n_1773),
.B(n_1727),
.Y(n_1777)
);

AOI322xp5_ASAP7_75t_L g1778 ( 
.A1(n_1768),
.A2(n_1764),
.A3(n_1722),
.B1(n_1732),
.B2(n_1724),
.C1(n_1729),
.C2(n_1727),
.Y(n_1778)
);

XNOR2x2_ASAP7_75t_L g1779 ( 
.A(n_1771),
.B(n_1731),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1776),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_SL g1782 ( 
.A(n_1775),
.B(n_1770),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1778),
.B(n_1767),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1779),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1775),
.B(n_1765),
.Y(n_1785)
);

AOI321xp33_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1772),
.A3(n_1724),
.B1(n_1732),
.B2(n_1729),
.C(n_1734),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1780),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1782),
.B(n_1734),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1781),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1784),
.A2(n_1664),
.B1(n_1695),
.B2(n_1683),
.Y(n_1790)
);

OR2x6_ASAP7_75t_L g1791 ( 
.A(n_1789),
.B(n_1783),
.Y(n_1791)
);

BUFx8_ASAP7_75t_SL g1792 ( 
.A(n_1787),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1788),
.A2(n_1782),
.B(n_1645),
.Y(n_1793)
);

XNOR2xp5_ASAP7_75t_L g1794 ( 
.A(n_1791),
.B(n_1790),
.Y(n_1794)
);

AOI32xp33_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1786),
.A3(n_1792),
.B1(n_1793),
.B2(n_1650),
.Y(n_1795)
);

INVx4_ASAP7_75t_L g1796 ( 
.A(n_1795),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1795),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1797),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1796),
.B(n_1652),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1799),
.A2(n_1796),
.B1(n_1695),
.B2(n_1683),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1798),
.A2(n_1690),
.B1(n_1662),
.B2(n_1663),
.Y(n_1801)
);

O2A1O1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1800),
.A2(n_1458),
.B(n_1690),
.C(n_1669),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1801),
.B(n_1657),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1669),
.B(n_1657),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1804),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1674),
.B1(n_1657),
.B2(n_1660),
.C(n_1669),
.Y(n_1806)
);

AOI211xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1452),
.B(n_1469),
.C(n_1479),
.Y(n_1807)
);


endmodule