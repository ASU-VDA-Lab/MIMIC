module real_jpeg_7306_n_15 (n_8, n_0, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_100, n_106, n_11, n_14, n_7, n_3, n_99, n_5, n_4, n_102, n_105, n_98, n_101, n_1, n_13, n_103, n_15);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_100;
input n_106;
input n_11;
input n_14;
input n_7;
input n_3;
input n_99;
input n_5;
input n_4;
input n_102;
input n_105;
input n_98;
input n_101;
input n_1;
input n_13;
input n_103;

output n_15;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_0),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_83),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_7),
.B(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_8),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_11),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_11),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_14),
.B(n_34),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_26),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_24),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_84),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_95),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_86),
.B(n_92),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21x1_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_82),
.B(n_85),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_75),
.B(n_81),
.Y(n_40)
);

AO221x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_51),
.B1(n_72),
.B2(n_73),
.C(n_74),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_71),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_70),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_66),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_80),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_98),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_99),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_100),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_101),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_102),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_103),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_104),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_105),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_106),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_107),
.Y(n_89)
);


endmodule