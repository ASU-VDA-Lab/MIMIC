module fake_jpeg_10459_n_208 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_17),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp67_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_27),
.B1(n_33),
.B2(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_45),
.Y(n_66)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_4),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_48),
.Y(n_74)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_37),
.B(n_32),
.C(n_33),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_57),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_61),
.Y(n_95)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_27),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_41),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_36),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_78),
.B(n_84),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_89),
.B1(n_90),
.B2(n_97),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_35),
.C(n_45),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_88),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_31),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_31),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_20),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_21),
.B1(n_28),
.B2(n_6),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_18),
.B1(n_22),
.B2(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_12),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_11),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_103),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_59),
.B1(n_53),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_72),
.B1(n_83),
.B2(n_86),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_77),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_108),
.Y(n_124)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_16),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_79),
.B(n_76),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_85),
.B(n_82),
.Y(n_131)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_128),
.B1(n_86),
.B2(n_102),
.C(n_13),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_78),
.B1(n_71),
.B2(n_70),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_139),
.B1(n_110),
.B2(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_6),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_73),
.C(n_85),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_120),
.C(n_103),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_87),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_82),
.B1(n_72),
.B2(n_87),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_102),
.B1(n_113),
.B2(n_108),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.C(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_141),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_134),
.C(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_120),
.C(n_118),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_119),
.A3(n_107),
.B1(n_104),
.B2(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_114),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_15),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_139),
.Y(n_161)
);

OA22x2_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_158)
);

NOR2x1_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_7),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_150),
.C(n_156),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_126),
.B(n_131),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_167),
.B(n_169),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_168),
.C(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_142),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_136),
.B(n_129),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_173),
.A2(n_158),
.B1(n_140),
.B2(n_123),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_148),
.C(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.Y(n_186)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_180),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_168),
.C(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_135),
.C(n_152),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_155),
.C(n_122),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_171),
.B1(n_167),
.B2(n_166),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_173),
.B(n_160),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_185),
.B(n_190),
.Y(n_197)
);

NAND4xp25_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_171),
.C(n_162),
.D(n_164),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_9),
.C(n_10),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_136),
.B(n_129),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_192),
.A2(n_193),
.B(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_132),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_132),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_9),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_11),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_12),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_197),
.A2(n_190),
.B(n_185),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_195),
.B(n_197),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_200),
.B(n_14),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_202),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_188),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_187),
.C(n_10),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_206),
.Y(n_208)
);


endmodule