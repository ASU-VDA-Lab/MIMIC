module fake_jpeg_24445_n_236 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_26),
.B1(n_21),
.B2(n_19),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_44),
.B1(n_14),
.B2(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_14),
.B1(n_27),
.B2(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_17),
.B1(n_27),
.B2(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_60),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_20),
.B1(n_22),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_52),
.B1(n_43),
.B2(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_63),
.A2(n_70),
.B1(n_47),
.B2(n_49),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_20),
.B1(n_31),
.B2(n_30),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_45),
.B(n_55),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_20),
.C(n_34),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_23),
.C(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_85),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_45),
.B1(n_48),
.B2(n_47),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_88),
.B1(n_84),
.B2(n_98),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_55),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_58),
.B(n_56),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_95),
.B(n_28),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_51),
.C(n_31),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_76),
.B1(n_61),
.B2(n_28),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_111),
.B1(n_113),
.B2(n_80),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_72),
.CI(n_62),
.CON(n_105),
.SN(n_105)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_75),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_63),
.B(n_69),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_118),
.B(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_67),
.B1(n_15),
.B2(n_23),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_67),
.B1(n_15),
.B2(n_25),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_119),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_57),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_90),
.C(n_91),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_82),
.B1(n_79),
.B2(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_139),
.Y(n_151)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_83),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_133),
.B(n_136),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_137),
.B1(n_138),
.B2(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.C(n_135),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_3),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_96),
.C(n_87),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_96),
.B(n_24),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_74),
.C(n_78),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_80),
.B(n_0),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_93),
.B1(n_97),
.B2(n_1),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_1),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_8),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_6),
.C2(n_7),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_149),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_112),
.B1(n_109),
.B2(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_142),
.B1(n_136),
.B2(n_134),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_111),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_156),
.B(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_153),
.A2(n_155),
.B(n_157),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_105),
.C(n_102),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_158),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_115),
.B1(n_107),
.B2(n_114),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_105),
.C(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_4),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_131),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_123),
.B1(n_140),
.B2(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_128),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_178),
.C(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

HAxp5_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_148),
.CON(n_188),
.SN(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_159),
.C(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_169),
.C(n_159),
.Y(n_198)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_190),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_192),
.B(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_176),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_198),
.C(n_203),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_194),
.B1(n_201),
.B2(n_189),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_204),
.B(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_207),
.Y(n_217)
);

NAND4xp25_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_180),
.C(n_184),
.D(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_183),
.C(n_186),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_210),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_185),
.C(n_172),
.Y(n_210)
);

FAx1_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_188),
.CI(n_185),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_6),
.Y(n_219)
);

AND2x4_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_148),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_13),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_207),
.A2(n_201),
.B(n_165),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_148),
.B1(n_150),
.B2(n_8),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_7),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_7),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_224),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_9),
.B(n_10),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_10),
.B(n_11),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_10),
.C(n_11),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_228),
.C(n_227),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_232),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_12),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_12),
.Y(n_236)
);


endmodule