module real_jpeg_32249_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_0),
.Y(n_161)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_0),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_0),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_37),
.B1(n_102),
.B2(n_105),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_1),
.A2(n_37),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_1),
.A2(n_37),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_4),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_5),
.A2(n_186),
.B1(n_222),
.B2(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_45),
.B1(n_91),
.B2(n_95),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_154),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_45),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_6),
.A2(n_45),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_6),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_6),
.B(n_110),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_6),
.A2(n_327),
.A3(n_329),
.B1(n_330),
.B2(n_336),
.Y(n_326)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_9),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_11),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_11),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_11),
.A2(n_127),
.B1(n_162),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_127),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_11),
.A2(n_127),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_377),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_251),
.B(n_375),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_212),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_16),
.B(n_212),
.Y(n_376)
);

OAI21xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_145),
.B(n_211),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_17),
.B(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_60),
.Y(n_17)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_18),
.B(n_61),
.C(n_99),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_19),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NOR2x1p5_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_20),
.Y(n_155)
);

AO22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_22),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_22),
.Y(n_205)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_25),
.Y(n_250)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_27),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_32),
.B(n_51),
.Y(n_235)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_46),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_47),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_45),
.A2(n_261),
.A3(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_45),
.B(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_45),
.B(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_45),
.B(n_366),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_46),
.Y(n_210)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_51),
.B(n_237),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_98),
.B1(n_99),
.B2(n_144),
.Y(n_60)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_76),
.B(n_90),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_62),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_62),
.B(n_90),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_62),
.B(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_62),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_63),
.Y(n_358)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_69),
.Y(n_316)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_69),
.Y(n_319)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_76),
.B(n_90),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_76),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_76),
.B(n_221),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_112)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_87),
.Y(n_278)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_94),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_94),
.Y(n_281)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_97),
.Y(n_270)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_121),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_100),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_132),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_107),
.Y(n_263)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_110),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g401 ( 
.A1(n_111),
.A2(n_133),
.B(n_245),
.Y(n_401)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AO21x2_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_134),
.B(n_138),
.Y(n_133)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_133),
.B(n_245),
.Y(n_294)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_181),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_146),
.B(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_147),
.B(n_182),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.C(n_156),
.Y(n_147)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_149),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_257)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_154),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2x1_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_171),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_158),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_159),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_161),
.Y(n_353)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_162),
.Y(n_328)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_165),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_165),
.B(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_184),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_172),
.B(n_313),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_182),
.Y(n_408)
);

HAxp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_191),
.CON(n_182),
.SN(n_182)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_191),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_188),
.B(n_190),
.Y(n_183)
);

AO21x2_ASAP7_75t_L g271 ( 
.A1(n_188),
.A2(n_216),
.B(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_190),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_190),
.B(n_310),
.Y(n_396)
);

OAI31xp33_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.A3(n_196),
.B(n_201),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_210),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_230),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_229),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_214),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_215),
.B(n_218),
.Y(n_399)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_219),
.B(n_289),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_220),
.B(n_275),
.Y(n_305)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_224),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_224),
.Y(n_395)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_229),
.B(n_230),
.C(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_231),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_233),
.A2(n_385),
.B(n_387),
.Y(n_384)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_234),
.A2(n_386),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_242),
.Y(n_386)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_284),
.B(n_374),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_282),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_254),
.B(n_282),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_273),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_273),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_260),
.A2(n_271),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_301),
.B(n_373),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_299),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_286),
.B(n_299),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_295),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_321)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_290),
.B(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_322),
.B(n_372),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_320),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_303),
.B(n_320),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

BUFx4f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_352),
.Y(n_351)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_348),
.B(n_371),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_345),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_345),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_343),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_326),
.B1(n_343),
.B2(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_355),
.B(n_370),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_SL g370 ( 
.A(n_350),
.B(n_354),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_362),
.Y(n_361)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_360),
.B(n_369),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_359),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_405),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2x1p5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_382),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_389),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_397),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_396),
.Y(n_390)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI22x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_404),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);


endmodule