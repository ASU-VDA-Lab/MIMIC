module fake_jpeg_16117_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_31),
.B(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_27),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_60),
.B1(n_64),
.B2(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_59),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_57),
.B1(n_61),
.B2(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_23),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_62),
.B1(n_19),
.B2(n_25),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_26),
.B1(n_29),
.B2(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_22),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_16),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_82),
.B1(n_83),
.B2(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_57),
.B1(n_34),
.B2(n_56),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_37),
.C(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_45),
.B1(n_39),
.B2(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_33),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_29),
.B1(n_35),
.B2(n_39),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_58),
.B1(n_49),
.B2(n_53),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_23),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_48),
.B(n_15),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_87),
.Y(n_115)
);

FAx1_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_50),
.CI(n_60),
.CON(n_87),
.SN(n_87)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_74),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_44),
.B1(n_46),
.B2(n_21),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_63),
.Y(n_97)
);

OR2x6_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_84),
.Y(n_125)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_44),
.B1(n_46),
.B2(n_34),
.Y(n_103)
);

OAI22x1_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_105),
.B1(n_107),
.B2(n_73),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_44),
.B1(n_56),
.B2(n_16),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_16),
.B1(n_21),
.B2(n_37),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_120),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_76),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_116),
.C(n_118),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_37),
.C(n_65),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_37),
.C(n_36),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_98),
.B1(n_87),
.B2(n_95),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_107),
.B(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_85),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_129),
.CI(n_36),
.CON(n_148),
.SN(n_148)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_93),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_73),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_86),
.A3(n_87),
.B1(n_92),
.B2(n_91),
.C1(n_93),
.C2(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_54),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_87),
.B(n_98),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_137),
.B(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_98),
.B1(n_94),
.B2(n_79),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_149),
.B1(n_79),
.B2(n_89),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_73),
.B(n_105),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_66),
.B1(n_75),
.B2(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_125),
.B1(n_126),
.B2(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_66),
.B1(n_75),
.B2(n_68),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_66),
.A3(n_81),
.B1(n_37),
.B2(n_24),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_110),
.B1(n_129),
.B2(n_116),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_108),
.C(n_122),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_154),
.C(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_54),
.C(n_72),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_101),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_139),
.B1(n_151),
.B2(n_135),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_163),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_136),
.B(n_9),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_165),
.B(n_11),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_0),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_164),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_133),
.B(n_146),
.Y(n_165)
);

INVxp33_ASAP7_75t_SL g167 ( 
.A(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_170),
.B1(n_162),
.B2(n_163),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_54),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_8),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_101),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_5),
.C(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_165),
.A2(n_151),
.B1(n_144),
.B2(n_137),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_181),
.B1(n_186),
.B2(n_161),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_132),
.C(n_148),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_132),
.C(n_148),
.Y(n_177)
);

HAxp5_ASAP7_75t_SL g203 ( 
.A(n_178),
.B(n_186),
.CON(n_203),
.SN(n_203)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_147),
.C(n_141),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_182),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_89),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_54),
.C(n_30),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_89),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_30),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_5),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_166),
.B(n_156),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_198),
.B(n_203),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_184),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_164),
.B1(n_155),
.B2(n_166),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_199),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_195),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_182),
.C(n_30),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_173),
.C(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_201),
.C(n_173),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_183),
.C(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_191),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_212),
.A2(n_197),
.B1(n_193),
.B2(n_203),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_13),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_204),
.C(n_6),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_207),
.B(n_1),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_199),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_11),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.C(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_209),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_219),
.B(n_224),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_230),
.B(n_1),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_207),
.B(n_12),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_237),
.C(n_227),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_3),
.C(n_4),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_3),
.C(n_4),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_235),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_242),
.B(n_4),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_245),
.B(n_4),
.Y(n_246)
);


endmodule