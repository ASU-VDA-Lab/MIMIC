module fake_jpeg_2037_n_268 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_67),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_60),
.Y(n_96)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_1),
.Y(n_60)
);

NAND2x1_ASAP7_75t_SL g61 ( 
.A(n_23),
.B(n_1),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_66),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_19),
.B(n_2),
.CON(n_70),
.SN(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_19),
.B(n_22),
.C(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_32),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_77),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_44),
.B1(n_26),
.B2(n_18),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_44),
.B1(n_26),
.B2(n_18),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_31),
.B1(n_40),
.B2(n_29),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_85),
.A2(n_102),
.B1(n_106),
.B2(n_108),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_45),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_28),
.C(n_37),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_5),
.C(n_8),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_63),
.B1(n_57),
.B2(n_41),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_28),
.B1(n_45),
.B2(n_33),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_33),
.B1(n_37),
.B2(n_29),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_103),
.B1(n_107),
.B2(n_100),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_79),
.B(n_90),
.C(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_40),
.B1(n_22),
.B2(n_25),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_56),
.A2(n_19),
.B1(n_61),
.B2(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_40),
.B1(n_19),
.B2(n_34),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_40),
.B1(n_34),
.B2(n_4),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_53),
.A2(n_2),
.B(n_3),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_114),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_111),
.B1(n_93),
.B2(n_95),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_133),
.Y(n_152)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_129),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_132),
.Y(n_173)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_9),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_9),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_12),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_140),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_107),
.B(n_102),
.C(n_116),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_81),
.A2(n_93),
.B1(n_101),
.B2(n_104),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_104),
.B1(n_111),
.B2(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_95),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_148),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_99),
.B1(n_112),
.B2(n_116),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_140),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_147),
.B1(n_134),
.B2(n_127),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_141),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_162),
.C(n_153),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_136),
.B1(n_119),
.B2(n_131),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_139),
.B1(n_121),
.B2(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_126),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_180),
.B1(n_183),
.B2(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_162),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_181),
.B(n_156),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_191),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_139),
.B1(n_128),
.B2(n_125),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_138),
.B(n_139),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_143),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_187),
.C(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_130),
.B1(n_149),
.B2(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_164),
.B(n_171),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_157),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_202),
.C(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_204),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_163),
.B(n_164),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_207),
.B(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_210),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_180),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_165),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_158),
.C(n_166),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_175),
.C(n_176),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_222),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_158),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_217),
.Y(n_234)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_201),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_219),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_204),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_178),
.C(n_183),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_199),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_198),
.B1(n_196),
.B2(n_195),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_215),
.B(n_225),
.Y(n_243)
);

AO22x1_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_196),
.B1(n_178),
.B2(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_211),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_193),
.B(n_208),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_229),
.B(n_226),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_214),
.CI(n_213),
.CON(n_238),
.SN(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_240),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_244),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_234),
.B(n_232),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_222),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_215),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_209),
.C(n_188),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_247),
.Y(n_253)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_234),
.C(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_251),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_208),
.C(n_219),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_252),
.B(n_245),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_232),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_238),
.B(n_203),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_250),
.C(n_238),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_257),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_253),
.B1(n_218),
.B2(n_203),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_191),
.B(n_185),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_265),
.A2(n_185),
.B1(n_189),
.B2(n_161),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_264),
.B(n_172),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_267),
.Y(n_268)
);


endmodule