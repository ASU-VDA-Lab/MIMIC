module fake_jpeg_2192_n_536 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_536);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_68),
.Y(n_127)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_31),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_70),
.Y(n_210)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_33),
.B(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_83),
.Y(n_130)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_80),
.Y(n_177)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_81),
.Y(n_183)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_39),
.B(n_15),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_42),
.B(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_86),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_15),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_19),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_88),
.B(n_115),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_13),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_93),
.Y(n_173)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_35),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_35),
.B1(n_52),
.B2(n_46),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_12),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_102),
.Y(n_186)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_55),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_104),
.B(n_106),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_27),
.B(n_14),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_21),
.B(n_0),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_108),
.B(n_112),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_11),
.Y(n_112)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_43),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_117),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_37),
.B(n_0),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

CKINVDCx11_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_19),
.Y(n_120)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_25),
.B(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_36),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_122),
.B(n_6),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_126),
.A2(n_109),
.B1(n_120),
.B2(n_113),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_129),
.B(n_134),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_36),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_46),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_138),
.B(n_141),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_30),
.B(n_43),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_140),
.A2(n_174),
.B(n_152),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_52),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_63),
.B(n_37),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_143),
.B(n_157),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_29),
.B1(n_23),
.B2(n_30),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_145),
.A2(n_49),
.B1(n_10),
.B2(n_11),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_64),
.B(n_30),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_150),
.B(n_151),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_2),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_153),
.B(n_155),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_94),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_4),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_4),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_4),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_168),
.B(n_180),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_61),
.A2(n_29),
.B1(n_23),
.B2(n_19),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_209),
.B1(n_49),
.B2(n_10),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_5),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_181),
.B(n_190),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_95),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_185),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_58),
.B(n_56),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_73),
.B(n_5),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_57),
.B(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_123),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_80),
.B(n_8),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_205),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_100),
.B(n_56),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_119),
.A2(n_29),
.B1(n_23),
.B2(n_51),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_69),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_214),
.A2(n_218),
.B1(n_226),
.B2(n_242),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_168),
.A2(n_84),
.B1(n_92),
.B2(n_89),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_215),
.A2(n_217),
.B1(n_219),
.B2(n_259),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_145),
.A2(n_87),
.B1(n_77),
.B2(n_72),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_109),
.B1(n_41),
.B2(n_51),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_170),
.A2(n_66),
.B1(n_71),
.B2(n_41),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_187),
.B1(n_125),
.B2(n_192),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_220),
.A2(n_221),
.B1(n_227),
.B2(n_240),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_268),
.B1(n_269),
.B2(n_276),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_9),
.B1(n_159),
.B2(n_194),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_186),
.A2(n_9),
.B1(n_209),
.B2(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_229),
.Y(n_330)
);

AO22x1_ASAP7_75t_SL g230 ( 
.A1(n_181),
.A2(n_193),
.B1(n_147),
.B2(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_231),
.B(n_255),
.Y(n_298)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_233),
.A2(n_248),
.B(n_282),
.Y(n_308)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_234),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_184),
.A2(n_162),
.B1(n_177),
.B2(n_210),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_147),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_254),
.Y(n_299)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_201),
.B1(n_176),
.B2(n_142),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_178),
.B1(n_180),
.B2(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_161),
.Y(n_243)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_130),
.A2(n_140),
.B(n_144),
.C(n_127),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_281),
.B(n_237),
.C(n_282),
.Y(n_296)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_173),
.A2(n_175),
.B1(n_200),
.B2(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_247),
.A2(n_260),
.B1(n_262),
.B2(n_267),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_156),
.B(n_160),
.C(n_162),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_206),
.Y(n_253)
);

BUFx4f_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_128),
.B(n_146),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_172),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_135),
.A2(n_176),
.B1(n_136),
.B2(n_142),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_177),
.A2(n_182),
.B1(n_169),
.B2(n_165),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_136),
.A2(n_199),
.B1(n_133),
.B2(n_182),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_175),
.A2(n_200),
.B1(n_195),
.B2(n_167),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_265),
.B1(n_283),
.B2(n_217),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_167),
.A2(n_179),
.B1(n_156),
.B2(n_199),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_266),
.B(n_273),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_148),
.A2(n_191),
.B1(n_154),
.B2(n_169),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_165),
.A2(n_163),
.B1(n_179),
.B2(n_183),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_165),
.A2(n_183),
.B1(n_132),
.B2(n_154),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_148),
.Y(n_271)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_154),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_139),
.A2(n_191),
.B1(n_132),
.B2(n_137),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_241),
.B1(n_233),
.B2(n_224),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_137),
.A2(n_145),
.B1(n_126),
.B2(n_112),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_171),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_278),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_168),
.A2(n_192),
.B1(n_190),
.B2(n_186),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_152),
.Y(n_284)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_261),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_290),
.B(n_310),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_222),
.B(n_235),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_293),
.B(n_296),
.Y(n_347)
);

AO21x2_ASAP7_75t_L g344 ( 
.A1(n_294),
.A2(n_274),
.B(n_278),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_307),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_230),
.B(n_238),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_295),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_231),
.B(n_256),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_315),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_261),
.Y(n_310)
);

NAND2x1p5_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_225),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_298),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_238),
.A2(n_256),
.B1(n_215),
.B2(n_244),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_332),
.B1(n_263),
.B2(n_265),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_254),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_213),
.C(n_279),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_229),
.C(n_234),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_272),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_317),
.B(n_334),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_264),
.B(n_255),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_318),
.B(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_212),
.B(n_216),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_324),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_212),
.B(n_216),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_249),
.B(n_284),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_335),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_248),
.B(n_219),
.CI(n_223),
.CON(n_331),
.SN(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_223),
.A2(n_246),
.B1(n_250),
.B2(n_262),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_246),
.B(n_250),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_333),
.B(n_315),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_251),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_249),
.B(n_228),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_362),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_291),
.A2(n_258),
.B1(n_245),
.B2(n_252),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_338),
.A2(n_346),
.B1(n_329),
.B2(n_301),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_308),
.A2(n_270),
.B(n_275),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_339),
.A2(n_350),
.B(n_361),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_291),
.A2(n_253),
.B1(n_239),
.B2(n_243),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_340),
.A2(n_344),
.B1(n_319),
.B2(n_323),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_352),
.C(n_363),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_307),
.A2(n_232),
.B1(n_257),
.B2(n_266),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_295),
.A2(n_273),
.B(n_277),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_296),
.B(n_271),
.C(n_278),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_321),
.B(n_271),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_353),
.B(n_356),
.Y(n_404)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_299),
.B(n_278),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_359),
.B(n_370),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_358),
.B(n_365),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_307),
.A2(n_324),
.B(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_309),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_312),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_294),
.B(n_303),
.C(n_325),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_368),
.C(n_285),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_285),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_288),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_373),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_292),
.A2(n_312),
.B(n_313),
.Y(n_370)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_287),
.Y(n_371)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_330),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_313),
.B(n_320),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_374),
.B(n_300),
.Y(n_397)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_371),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_322),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_380),
.B(n_382),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_351),
.Y(n_382)
);

A2O1A1O1Ixp25_ASAP7_75t_L g385 ( 
.A1(n_347),
.A2(n_331),
.B(n_302),
.C(n_286),
.D(n_285),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_385),
.A2(n_359),
.B(n_357),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_322),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_351),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_397),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_285),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_400),
.C(n_403),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_368),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_348),
.A2(n_286),
.B1(n_331),
.B2(n_304),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_392),
.A2(n_395),
.B1(n_401),
.B2(n_337),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_348),
.A2(n_304),
.B1(n_323),
.B2(n_328),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_320),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_396),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_398),
.A2(n_346),
.B1(n_338),
.B2(n_337),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_345),
.B(n_330),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_348),
.A2(n_328),
.B1(n_306),
.B2(n_297),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_342),
.B(n_297),
.C(n_306),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_379),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_407),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_410),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_414),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_345),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_384),
.A2(n_344),
.B1(n_365),
.B2(n_362),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_412),
.A2(n_416),
.B1(n_420),
.B2(n_424),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_413),
.A2(n_426),
.B1(n_429),
.B2(n_430),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_377),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_389),
.A2(n_357),
.B(n_370),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_415),
.A2(n_375),
.B(n_404),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_384),
.A2(n_344),
.B1(n_336),
.B2(n_361),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_381),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_417),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_383),
.B(n_361),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_419),
.B(n_400),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_382),
.A2(n_344),
.B1(n_339),
.B2(n_356),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_387),
.A2(n_344),
.B1(n_367),
.B2(n_340),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_381),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_427),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_404),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_428),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_378),
.A2(n_385),
.B1(n_389),
.B2(n_392),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_388),
.A2(n_352),
.B1(n_364),
.B2(n_374),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_398),
.A2(n_358),
.B1(n_350),
.B2(n_349),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_432),
.A2(n_399),
.B1(n_402),
.B2(n_394),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_433),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_403),
.C(n_391),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_441),
.C(n_408),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_446),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_440),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_415),
.A2(n_375),
.B(n_376),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_393),
.C(n_405),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_402),
.B1(n_399),
.B2(n_394),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_442),
.A2(n_432),
.B1(n_426),
.B2(n_409),
.Y(n_465)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_444),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_419),
.B(n_393),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_448),
.A2(n_452),
.B1(n_420),
.B2(n_424),
.Y(n_459)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_449),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_369),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_450),
.B(n_455),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_423),
.A2(n_390),
.B1(n_395),
.B2(n_366),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_410),
.B(n_401),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_412),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_418),
.B(n_372),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_431),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_465),
.B1(n_473),
.B2(n_476),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_468),
.C(n_469),
.Y(n_492)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_431),
.Y(n_464)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_407),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_444),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_430),
.C(n_411),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_429),
.C(n_427),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_474),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_447),
.A2(n_417),
.B1(n_406),
.B2(n_422),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_406),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_416),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_475),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_453),
.A2(n_456),
.B1(n_439),
.B2(n_436),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_414),
.C(n_354),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_477),
.B(n_478),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_390),
.C(n_373),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_453),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_483),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_464),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_445),
.Y(n_484)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_484),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_456),
.Y(n_485)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_485),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_461),
.A2(n_451),
.B1(n_448),
.B2(n_445),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_440),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_488),
.B(n_452),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_490),
.A2(n_491),
.B1(n_438),
.B2(n_472),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_439),
.B1(n_469),
.B2(n_438),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_486),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_496),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_460),
.C(n_475),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_502),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_492),
.B(n_468),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_503),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_478),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_489),
.A2(n_451),
.B(n_437),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_477),
.C(n_446),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_470),
.Y(n_515)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_505),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_499),
.A2(n_488),
.B1(n_482),
.B2(n_484),
.Y(n_507)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_507),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g509 ( 
.A(n_498),
.B(n_483),
.CI(n_484),
.CON(n_509),
.SN(n_509)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_511),
.Y(n_516)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_515),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_492),
.C(n_496),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_520),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_481),
.Y(n_519)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_519),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_502),
.C(n_504),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_508),
.A2(n_487),
.B(n_490),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_522),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_471),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_513),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_527),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_519),
.A2(n_513),
.B1(n_463),
.B2(n_442),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_516),
.B(n_523),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_525),
.B(n_524),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_526),
.A2(n_509),
.B(n_515),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_524),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_533),
.B1(n_531),
.B2(n_509),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_470),
.B(n_458),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_449),
.Y(n_536)
);


endmodule