module fake_jpeg_12534_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_23),
.C(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_10),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_14),
.B(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_17),
.B1(n_12),
.B2(n_14),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_23),
.B1(n_17),
.B2(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_17),
.B1(n_12),
.B2(n_15),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_26),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_1),
.B(n_4),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_13),
.B1(n_11),
.B2(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_35),
.B1(n_34),
.B2(n_9),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_9),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_40),
.C(n_43),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_41),
.B1(n_4),
.B2(n_6),
.Y(n_54)
);

AO22x1_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_44),
.B(n_46),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_41),
.C(n_4),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_54),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_48),
.C(n_49),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_5),
.Y(n_59)
);

AOI31xp67_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_55),
.A3(n_53),
.B(n_7),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.CI(n_6),
.CON(n_60),
.SN(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_7),
.C(n_37),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_60),
.B(n_37),
.Y(n_62)
);


endmodule