module fake_netlist_6_1084_n_598 (n_52, n_16, n_1, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_42, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_598);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_42;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_598;

wire n_591;
wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_125;
wire n_384;
wire n_297;
wire n_595;
wire n_524;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_92;
wire n_513;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_548;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_596;
wire n_123;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_99;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_5),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_7),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_25),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_27),
.Y(n_100)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_12),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_6),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_23),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_26),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g111 ( 
.A(n_37),
.B(n_67),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_18),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_46),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_0),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_0),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_34),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_32),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_12),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_18),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_50),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_3),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_82),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_29),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_70),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_13),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_39),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_60),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_33),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_48),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_42),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_86),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_35),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_24),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_15),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_31),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_16),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_80),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_49),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx2_ASAP7_75t_SL g154 ( 
.A(n_65),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_7),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_45),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_28),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_71),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_73),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_47),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_14),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_40),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_38),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_43),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_109),
.B(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_112),
.B(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_112),
.B(n_4),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_95),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_119),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_4),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_117),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_95),
.B(n_11),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

OAI22x1_ASAP7_75t_SL g201 ( 
.A1(n_119),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

AOI22x1_ASAP7_75t_SL g204 ( 
.A1(n_126),
.A2(n_30),
.B1(n_44),
.B2(n_51),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_94),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_156),
.A2(n_53),
.B(n_55),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_83),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_150),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_139),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_98),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_103),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_105),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_149),
.B(n_59),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_96),
.B(n_63),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

OR2x6_ASAP7_75t_L g240 ( 
.A(n_154),
.B(n_64),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

AOI22x1_ASAP7_75t_SL g244 ( 
.A1(n_126),
.A2(n_77),
.B1(n_110),
.B2(n_121),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_163),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_102),
.B(n_115),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_129),
.B(n_172),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_177),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

AND3x2_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_132),
.C(n_101),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_93),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_161),
.C(n_100),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_196),
.B(n_152),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_188),
.A2(n_101),
.B1(n_152),
.B2(n_122),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_122),
.B1(n_121),
.B2(n_110),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_133),
.B1(n_100),
.B2(n_108),
.Y(n_272)
);

OR2x6_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_111),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_99),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_181),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_184),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_187),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_182),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_142),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_217),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_180),
.A2(n_108),
.B1(n_162),
.B2(n_155),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_174),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_114),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_174),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_221),
.B(n_162),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_184),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_196),
.B(n_155),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_221),
.B(n_137),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_192),
.B(n_118),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_L g295 ( 
.A(n_188),
.B(n_130),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_221),
.B(n_130),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_221),
.B(n_193),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_183),
.B(n_134),
.C(n_137),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_193),
.B(n_134),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_178),
.B(n_140),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_178),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_182),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_191),
.A2(n_144),
.B1(n_146),
.B2(n_151),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_185),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_222),
.B(n_228),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_191),
.B(n_217),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_223),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_178),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_197),
.B(n_223),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_185),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_228),
.B(n_190),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_179),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_220),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_228),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_306),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_222),
.Y(n_319)
);

NAND2xp33_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_200),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_240),
.B1(n_227),
.B2(n_197),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_285),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_278),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_266),
.A2(n_240),
.B1(n_222),
.B2(n_227),
.Y(n_326)
);

NOR2x2_ASAP7_75t_L g327 ( 
.A(n_273),
.B(n_240),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_239),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_282),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g330 ( 
.A(n_267),
.B(n_219),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_222),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_229),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_289),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_272),
.B(n_189),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_190),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

NOR2x2_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_240),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_263),
.B(n_242),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_309),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_229),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_273),
.A2(n_245),
.B1(n_251),
.B2(n_250),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_231),
.B(n_233),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_238),
.Y(n_344)
);

NAND2x1_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_219),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_239),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_286),
.B(n_238),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_288),
.A2(n_242),
.B1(n_251),
.B2(n_250),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_267),
.B(n_195),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_239),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_299),
.B(n_249),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_L g354 ( 
.A(n_292),
.B(n_214),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_241),
.B1(n_249),
.B2(n_243),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_239),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_257),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_274),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_229),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_258),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_245),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_283),
.B(n_300),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_299),
.B(n_243),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_284),
.B(n_241),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_295),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_305),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_295),
.Y(n_369)
);

O2A1O1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_351),
.A2(n_232),
.B(n_236),
.C(n_237),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_275),
.Y(n_372)
);

AOI21xp33_ASAP7_75t_L g373 ( 
.A1(n_322),
.A2(n_269),
.B(n_307),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_353),
.A2(n_305),
.B1(n_279),
.B2(n_300),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_328),
.A2(n_219),
.B(n_268),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_262),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_330),
.A2(n_219),
.B1(n_252),
.B2(n_246),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g378 ( 
.A1(n_354),
.A2(n_226),
.B(n_224),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_293),
.Y(n_379)
);

CKINVDCx10_ASAP7_75t_R g380 ( 
.A(n_329),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_300),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_246),
.B1(n_252),
.B2(n_237),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_207),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_320),
.A2(n_268),
.B(n_271),
.Y(n_386)
);

O2A1O1Ixp5_ASAP7_75t_L g387 ( 
.A1(n_345),
.A2(n_265),
.B(n_252),
.C(n_246),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_320),
.A2(n_332),
.B(n_341),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_215),
.B1(n_310),
.B2(n_277),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_300),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_316),
.A2(n_318),
.B(n_364),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_192),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_265),
.B(n_294),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_280),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_204),
.B1(n_304),
.B2(n_302),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_352),
.A2(n_294),
.B(n_308),
.Y(n_398)
);

NOR2x1_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_201),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_312),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_319),
.B(n_340),
.Y(n_401)
);

A2O1A1Ixp33_ASAP7_75t_L g402 ( 
.A1(n_343),
.A2(n_194),
.B(n_213),
.C(n_225),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_342),
.B(n_194),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_213),
.B(n_224),
.C(n_225),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_313),
.A2(n_294),
.B(n_308),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_SL g407 ( 
.A(n_326),
.B(n_244),
.C(n_202),
.Y(n_407)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_201),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_340),
.A2(n_215),
.B1(n_220),
.B2(n_214),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_350),
.A2(n_215),
.B1(n_220),
.B2(n_214),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_333),
.A2(n_204),
.B1(n_244),
.B2(n_226),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_360),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_337),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_360),
.A2(n_294),
.B(n_308),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_355),
.A2(n_220),
.B1(n_214),
.B2(n_200),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_349),
.A2(n_214),
.B1(n_220),
.B2(n_208),
.Y(n_417)
);

AOI21xp33_ASAP7_75t_L g418 ( 
.A1(n_362),
.A2(n_210),
.B(n_212),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_360),
.A2(n_261),
.B(n_290),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_337),
.A2(n_308),
.B(n_301),
.Y(n_421)
);

A2O1A1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_347),
.A2(n_209),
.B(n_205),
.C(n_199),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_SL g423 ( 
.A1(n_347),
.A2(n_209),
.B(n_205),
.C(n_199),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_362),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_357),
.A2(n_301),
.B(n_276),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_358),
.A2(n_220),
.B1(n_208),
.B2(n_209),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_358),
.Y(n_429)
);

AOI22x1_ASAP7_75t_L g430 ( 
.A1(n_327),
.A2(n_208),
.B1(n_206),
.B2(n_203),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_338),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_367),
.B(n_338),
.Y(n_432)
);

AOI221x1_ASAP7_75t_L g433 ( 
.A1(n_377),
.A2(n_392),
.B1(n_391),
.B2(n_381),
.C(n_389),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_419),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_420),
.A2(n_301),
.B(n_276),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_374),
.A2(n_208),
.B1(n_205),
.B2(n_203),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_400),
.A2(n_301),
.B(n_276),
.Y(n_437)
);

NAND3x1_ASAP7_75t_L g438 ( 
.A(n_393),
.B(n_408),
.C(n_399),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_210),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_387),
.A2(n_206),
.B(n_207),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_388),
.A2(n_290),
.B(n_198),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

AO31x2_ASAP7_75t_L g443 ( 
.A1(n_378),
.A2(n_211),
.A3(n_212),
.B(n_179),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

AO31x2_ASAP7_75t_L g447 ( 
.A1(n_409),
.A2(n_179),
.A3(n_198),
.B(n_422),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_179),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_386),
.A2(n_179),
.B(n_198),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_403),
.A2(n_198),
.B(n_412),
.Y(n_450)
);

AOI221x1_ASAP7_75t_L g451 ( 
.A1(n_396),
.A2(n_198),
.B1(n_390),
.B2(n_417),
.C(n_407),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_368),
.B(n_424),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_372),
.B(n_383),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_385),
.A2(n_413),
.B(n_398),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_394),
.A2(n_425),
.B(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_430),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_431),
.Y(n_457)
);

AOI221x1_ASAP7_75t_L g458 ( 
.A1(n_405),
.A2(n_416),
.B1(n_427),
.B2(n_410),
.C(n_418),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g459 ( 
.A1(n_376),
.A2(n_401),
.B1(n_411),
.B2(n_397),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_395),
.A2(n_414),
.B(n_406),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

INVx3_ASAP7_75t_SL g462 ( 
.A(n_376),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_401),
.A2(n_423),
.B(n_380),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_380),
.B(n_367),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_380),
.Y(n_469)
);

AOI31xp67_ASAP7_75t_L g470 ( 
.A1(n_381),
.A2(n_391),
.A3(n_385),
.B(n_371),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_426),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_372),
.B(n_329),
.Y(n_473)
);

AOI221xp5_ASAP7_75t_L g474 ( 
.A1(n_373),
.A2(n_351),
.B1(n_267),
.B2(n_322),
.C(n_393),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_389),
.A2(n_320),
.B(n_314),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_384),
.B(n_368),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_424),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

A2O1A1Ixp33_ASAP7_75t_L g480 ( 
.A1(n_369),
.A2(n_323),
.B(n_367),
.C(n_373),
.Y(n_480)
);

NAND3x1_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_408),
.C(n_399),
.Y(n_481)
);

AO32x2_ASAP7_75t_L g482 ( 
.A1(n_377),
.A2(n_382),
.A3(n_322),
.B1(n_409),
.B2(n_390),
.Y(n_482)
);

AOI221xp5_ASAP7_75t_SL g483 ( 
.A1(n_402),
.A2(n_351),
.B1(n_322),
.B2(n_323),
.C(n_367),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_375),
.A2(n_387),
.B(n_420),
.Y(n_484)
);

AOI221xp5_ASAP7_75t_L g485 ( 
.A1(n_474),
.A2(n_459),
.B1(n_483),
.B2(n_432),
.C(n_465),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_453),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_459),
.A2(n_434),
.B1(n_468),
.B2(n_472),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_445),
.Y(n_490)
);

AO31x2_ASAP7_75t_L g491 ( 
.A1(n_433),
.A2(n_451),
.A3(n_458),
.B(n_436),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_449),
.A2(n_454),
.B(n_461),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_482),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_439),
.B(n_452),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_475),
.A2(n_456),
.B(n_457),
.C(n_476),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_463),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_440),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_437),
.B(n_441),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

OAI21x1_ASAP7_75t_SL g502 ( 
.A1(n_464),
.A2(n_450),
.B(n_460),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_471),
.B(n_477),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_477),
.A2(n_438),
.B(n_481),
.Y(n_505)
);

NAND2x1p5_ASAP7_75t_L g506 ( 
.A(n_446),
.B(n_477),
.Y(n_506)
);

BUFx4f_ASAP7_75t_SL g507 ( 
.A(n_462),
.Y(n_507)
);

AO31x2_ASAP7_75t_L g508 ( 
.A1(n_470),
.A2(n_482),
.A3(n_443),
.B(n_484),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_467),
.B(n_455),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_469),
.B(n_447),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_447),
.B(n_393),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_471),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_323),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_487),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_514),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_499),
.Y(n_517)
);

NOR2x1_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_490),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_513),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_495),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_511),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_494),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_511),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_488),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_497),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_509),
.Y(n_528)
);

CKINVDCx11_ASAP7_75t_R g529 ( 
.A(n_503),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_509),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_517),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_510),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_508),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_504),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_492),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_491),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_521),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_SL g539 ( 
.A(n_526),
.B(n_505),
.C(n_506),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_506),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

AO21x2_ASAP7_75t_L g543 ( 
.A1(n_531),
.A2(n_509),
.B(n_500),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_501),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_519),
.B(n_501),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_533),
.B(n_530),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_515),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_520),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_543),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_521),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_538),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_543),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_541),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_532),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_543),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_532),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_524),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_528),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_553),
.B(n_536),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_528),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_542),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_554),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_534),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_556),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_542),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_547),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_555),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_555),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_552),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_564),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_552),
.Y(n_571)
);

O2A1O1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_565),
.A2(n_539),
.B(n_526),
.C(n_540),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_562),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_529),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_549),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_570),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_570),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_575),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_573),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_575),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_576),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_579),
.A2(n_572),
.B(n_574),
.C(n_577),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_578),
.B(n_571),
.Y(n_583)
);

OAI221xp5_ASAP7_75t_L g584 ( 
.A1(n_582),
.A2(n_546),
.B1(n_580),
.B2(n_571),
.C(n_568),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_581),
.A2(n_546),
.B(n_567),
.Y(n_585)
);

OAI211xp5_ASAP7_75t_SL g586 ( 
.A1(n_584),
.A2(n_585),
.B(n_583),
.C(n_580),
.Y(n_586)
);

OAI211xp5_ASAP7_75t_SL g587 ( 
.A1(n_584),
.A2(n_544),
.B(n_518),
.C(n_537),
.Y(n_587)
);

AOI211xp5_ASAP7_75t_L g588 ( 
.A1(n_586),
.A2(n_567),
.B(n_537),
.C(n_527),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_587),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_569),
.Y(n_590)
);

NAND4xp75_ASAP7_75t_L g591 ( 
.A(n_588),
.B(n_518),
.C(n_569),
.D(n_568),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_591),
.A2(n_567),
.B1(n_558),
.B2(n_560),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_590),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_593),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_594),
.A2(n_507),
.B1(n_558),
.B2(n_560),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_595),
.A2(n_524),
.B(n_515),
.C(n_527),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_596),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_597),
.A2(n_501),
.B(n_512),
.Y(n_598)
);


endmodule