module fake_jpeg_835_n_42 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_42);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_6),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_15),
.B(n_17),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B(n_14),
.C(n_16),
.D(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_15),
.B1(n_14),
.B2(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_16),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_32),
.B1(n_26),
.B2(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_3),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_12),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_4),
.C(n_5),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_34),
.C(n_33),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_36),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_4),
.C2(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);


endmodule