module fake_ariane_239_n_2865 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2865);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2865;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2663;
wire n_559;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_762;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_1491;
wire n_931;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_2147;
wire n_867;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_727;
wire n_590;
wire n_699;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2418;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_742;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_2448;
wire n_812;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_1700;
wire n_862;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_1659;
wire n_885;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_2647;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_1968;
wire n_918;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_1653;
wire n_872;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_1663;
wire n_919;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_1809;
wire n_765;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2324;
wire n_2153;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_671;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_2297;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_2673;
wire n_1591;
wire n_664;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_537;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_803;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_548;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_444),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_524),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_522),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_130),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_376),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_373),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_290),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_251),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_309),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_426),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_333),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_471),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_414),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_124),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_68),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_176),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_383),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_490),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_434),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_412),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_219),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_84),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_103),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_112),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_157),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_485),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_406),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_116),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_188),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_378),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_117),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_48),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_266),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_329),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_94),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_520),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_204),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_364),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_224),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_517),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_238),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_495),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_462),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_134),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_102),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_60),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_120),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_111),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_10),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_28),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_504),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_415),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_62),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_329),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_348),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_9),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_18),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_246),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_243),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_222),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_80),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_422),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_33),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_394),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_493),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_2),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_116),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_230),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_438),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_389),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_67),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_62),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_432),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_122),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_435),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_194),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_366),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_147),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_162),
.Y(n_606)
);

CKINVDCx14_ASAP7_75t_R g607 ( 
.A(n_442),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_173),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_245),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_31),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_404),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_478),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_441),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_269),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_134),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_310),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_100),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_374),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_510),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_526),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_501),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_421),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_74),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_258),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_206),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_319),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_402),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_392),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_335),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_275),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_183),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_400),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_443),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_165),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_377),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_391),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_169),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_499),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_511),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_312),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_228),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_473),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_202),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_301),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_262),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_440),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_25),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_28),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_188),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_416),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_371),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_494),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_121),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_57),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_191),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_428),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_375),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_297),
.Y(n_658)
);

CKINVDCx14_ASAP7_75t_R g659 ( 
.A(n_156),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_496),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_457),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_45),
.Y(n_662)
);

BUFx2_ASAP7_75t_SL g663 ( 
.A(n_129),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_298),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_156),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_449),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_447),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_0),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_58),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_361),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_95),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_107),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_350),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_60),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_497),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_135),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_290),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_78),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_353),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_321),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_85),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_204),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_328),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_36),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_27),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_179),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_353),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_152),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_158),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_463),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_106),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_26),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_386),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_112),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_44),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_293),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_70),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_149),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_72),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_507),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_487),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_513),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_166),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_291),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_271),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_179),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_121),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_260),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_262),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_500),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_425),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_399),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_445),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_503),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_88),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_488),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_396),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_120),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_211),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_318),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_361),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_180),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_45),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_299),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_344),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_519),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_18),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_486),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_76),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_481),
.Y(n_730)
);

CKINVDCx11_ASAP7_75t_R g731 ( 
.A(n_450),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_436),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_472),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_475),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_234),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_0),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_304),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_76),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_506),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_508),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_489),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_417),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_349),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_193),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_113),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_505),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_315),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_81),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_515),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_10),
.Y(n_750)
);

CKINVDCx16_ASAP7_75t_R g751 ( 
.A(n_315),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_408),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_88),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_304),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_195),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_351),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_32),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_461),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_476),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_350),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_470),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_319),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_80),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_218),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_407),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_24),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_333),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_190),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_327),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_292),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_107),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_73),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_12),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_388),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_355),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_71),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_431),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_191),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_458),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_232),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_123),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_227),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_96),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_479),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_498),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_429),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_122),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_284),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_29),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_446),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_433),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_424),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_516),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_284),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_142),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_195),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_301),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_380),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_322),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_71),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_477),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_288),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_410),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_459),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_206),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_448),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_401),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_217),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_390),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_181),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_521),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_381),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_287),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_85),
.Y(n_814)
);

BUFx5_ASAP7_75t_L g815 ( 
.A(n_90),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_232),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_430),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_452),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_56),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_20),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_512),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_79),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_403),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_126),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_379),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_337),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_165),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_14),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_234),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_317),
.Y(n_830)
);

BUFx10_ASAP7_75t_L g831 ( 
.A(n_456),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_306),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_169),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_397),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_395),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_61),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_269),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_162),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_133),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_365),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_326),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_320),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_214),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_525),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_292),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_209),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_323),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_468),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_55),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_148),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_69),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_464),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_372),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_393),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_111),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_311),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_320),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_514),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_418),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_349),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_277),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_302),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_243),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_411),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_483),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_370),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_423),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_170),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_199),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_67),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_96),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_61),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_491),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_265),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_149),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_356),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_368),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_398),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_124),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_310),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_100),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_482),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_427),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_155),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_265),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_5),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_460),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_300),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_252),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_352),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_127),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_465),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_193),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_260),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_145),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_439),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_146),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_324),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_405),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_95),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_213),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_159),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_247),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_502),
.Y(n_904)
);

BUFx10_ASAP7_75t_L g905 ( 
.A(n_47),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_226),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_224),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_330),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_474),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_259),
.Y(n_910)
);

BUFx5_ASAP7_75t_L g911 ( 
.A(n_313),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_189),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_196),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_79),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_342),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_518),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_413),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_454),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_210),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_87),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_198),
.Y(n_921)
);

CKINVDCx16_ASAP7_75t_R g922 ( 
.A(n_141),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_145),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_466),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_210),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_66),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_480),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_264),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_336),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_367),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_409),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_233),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_9),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_259),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_492),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_360),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_36),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_523),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_419),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_286),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_420),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_382),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_323),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_127),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_385),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_185),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_437),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_453),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_117),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_387),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_509),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_469),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_190),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_484),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_384),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_229),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_467),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_455),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_82),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_15),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_317),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_659),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_623),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_623),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_623),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_561),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_557),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_561),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_574),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_574),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_585),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_644),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_585),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_637),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_637),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_685),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_685),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_815),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_815),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_691),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_691),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_736),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_634),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_736),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_764),
.Y(n_985)
);

INVxp33_ASAP7_75t_SL g986 ( 
.A(n_540),
.Y(n_986)
);

INVxp33_ASAP7_75t_L g987 ( 
.A(n_894),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_764),
.Y(n_988)
);

INVxp33_ASAP7_75t_L g989 ( 
.A(n_933),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_750),
.Y(n_990)
);

CKINVDCx16_ASAP7_75t_R g991 ( 
.A(n_737),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_778),
.Y(n_992)
);

INVxp33_ASAP7_75t_SL g993 ( 
.A(n_530),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_778),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_937),
.Y(n_995)
);

CKINVDCx16_ASAP7_75t_R g996 ( 
.A(n_751),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_937),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_961),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_641),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_961),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_815),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_815),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_815),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_815),
.Y(n_1004)
);

INVxp67_ASAP7_75t_SL g1005 ( 
.A(n_624),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_815),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_815),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_911),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_731),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_911),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_911),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_911),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_726),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_911),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_662),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_624),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_911),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_911),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_911),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_549),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_564),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_718),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_624),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_624),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_795),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_565),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_624),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_533),
.Y(n_1028)
);

CKINVDCx14_ASAP7_75t_R g1029 ( 
.A(n_607),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_570),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_571),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_584),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_586),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_588),
.Y(n_1034)
);

CKINVDCx16_ASAP7_75t_R g1035 ( 
.A(n_840),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_922),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_1013),
.Y(n_1037)
);

OA21x2_ASAP7_75t_L g1038 ( 
.A1(n_1001),
.A2(n_544),
.B(n_538),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_1023),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1028),
.B(n_635),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_978),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1023),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1024),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_1024),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1013),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1013),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_986),
.A2(n_727),
.B1(n_738),
.B2(n_725),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1029),
.B(n_730),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_978),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_1036),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_977),
.B(n_784),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_1013),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_979),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_1002),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_979),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1003),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_994),
.B(n_963),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_1004),
.A2(n_568),
.B(n_552),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_1006),
.A2(n_602),
.B(n_577),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_1007),
.A2(n_613),
.B(n_611),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1008),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_964),
.B(n_548),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_SL g1063 ( 
.A1(n_983),
.A2(n_771),
.B1(n_799),
.B2(n_770),
.Y(n_1063)
);

BUFx8_ASAP7_75t_L g1064 ( 
.A(n_1036),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1029),
.B(n_620),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_1010),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1011),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_966),
.B(n_968),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_1009),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1012),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_SL g1071 ( 
.A1(n_983),
.A2(n_820),
.B1(n_822),
.B2(n_814),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_1014),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1017),
.A2(n_632),
.B(n_622),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1018),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_969),
.B(n_590),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_991),
.Y(n_1076)
);

CKINVDCx8_ASAP7_75t_R g1077 ( 
.A(n_1009),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_965),
.B(n_1005),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1019),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_967),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_970),
.B(n_590),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_999),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1016),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1027),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_986),
.A2(n_989),
.B1(n_987),
.B2(n_972),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_971),
.B(n_536),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_973),
.B(n_636),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1020),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1021),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_990),
.A2(n_888),
.B1(n_903),
.B2(n_875),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_L g1091 ( 
.A(n_974),
.B(n_536),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_975),
.B(n_548),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_976),
.B(n_590),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1026),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_1030),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_996),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1031),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1069),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1069),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1040),
.B(n_987),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1080),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1082),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1056),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1054),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1056),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_1050),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1088),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1067),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_1077),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1077),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1064),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_R g1112 ( 
.A(n_1050),
.B(n_993),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1064),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1088),
.Y(n_1114)
);

CKINVDCx16_ASAP7_75t_R g1115 ( 
.A(n_1076),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1083),
.B(n_962),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1067),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1083),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1064),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_1057),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1064),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1096),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1063),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1063),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1084),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1047),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1084),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1071),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1057),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1071),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1089),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1070),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_1047),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1040),
.B(n_989),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1090),
.Y(n_1135)
);

BUFx10_ASAP7_75t_L g1136 ( 
.A(n_1057),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1090),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1070),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1054),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1089),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1095),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1095),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1051),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1051),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1095),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1094),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1057),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1095),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_1075),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1054),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1053),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1085),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1053),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_1078),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1048),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1154),
.B(n_1120),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1103),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1154),
.B(n_1053),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1147),
.B(n_1075),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1100),
.B(n_1035),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1118),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1150),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1125),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1127),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1131),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1147),
.B(n_1081),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1152),
.A2(n_1058),
.B1(n_1059),
.B2(n_1038),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1143),
.B(n_1065),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1154),
.B(n_1053),
.Y(n_1169)
);

AND2x6_ASAP7_75t_SL g1170 ( 
.A(n_1134),
.B(n_608),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1140),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1120),
.B(n_1041),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1155),
.B(n_1081),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1146),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_1104),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1151),
.B(n_1041),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1151),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1102),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1155),
.B(n_1093),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1144),
.A2(n_1093),
.B1(n_993),
.B2(n_1078),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1152),
.A2(n_1058),
.B1(n_1059),
.B2(n_1038),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1150),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1104),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1153),
.B(n_1049),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1120),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1106),
.B(n_972),
.Y(n_1186)
);

AND2x2_ASAP7_75t_SL g1187 ( 
.A(n_1153),
.B(n_532),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_1129),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1129),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1103),
.B(n_1049),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1107),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1122),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1115),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1105),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1114),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1105),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1110),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1108),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1112),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1108),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1117),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1129),
.Y(n_1203)
);

AND2x2_ASAP7_75t_SL g1204 ( 
.A(n_1104),
.B(n_532),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1136),
.A2(n_1078),
.B1(n_545),
.B2(n_758),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1136),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1098),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1117),
.B(n_1055),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1132),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1132),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1136),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1149),
.B(n_1025),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1139),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1126),
.A2(n_1092),
.B1(n_1062),
.B2(n_663),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1138),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1138),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1141),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1139),
.Y(n_1218)
);

OAI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1116),
.A2(n_868),
.B(n_615),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1139),
.A2(n_1055),
.B(n_1061),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1142),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1145),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1113),
.B(n_1068),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1149),
.B(n_962),
.C(n_1061),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1148),
.B(n_1078),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1121),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1111),
.B(n_1068),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1135),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1137),
.B(n_1074),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1099),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1111),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_L g1232 ( 
.A(n_1123),
.B(n_1079),
.C(n_1074),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1128),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1176),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1204),
.A2(n_925),
.B1(n_926),
.B2(n_915),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1177),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1176),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1192),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1177),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1184),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1160),
.B(n_1124),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1198),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1192),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1178),
.B(n_1094),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1159),
.B(n_1119),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1157),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_1228),
.A2(n_1133),
.B1(n_1126),
.B2(n_1130),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1159),
.B(n_1119),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1168),
.A2(n_1073),
.B(n_1079),
.C(n_876),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1173),
.B(n_999),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1194),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1207),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1161),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1199),
.Y(n_1254)
);

NAND2x1p5_ASAP7_75t_L g1255 ( 
.A(n_1230),
.B(n_1095),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1193),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1173),
.A2(n_759),
.B1(n_811),
.B2(n_529),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1179),
.B(n_1015),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1168),
.B(n_1097),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1163),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1184),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1201),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1189),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1196),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1182),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1229),
.B(n_1097),
.Y(n_1266)
);

AO22x2_ASAP7_75t_L g1267 ( 
.A1(n_1214),
.A2(n_1133),
.B1(n_1130),
.B2(n_1128),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1209),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1197),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1202),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1210),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1215),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1189),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1200),
.B(n_1179),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1200),
.B(n_1015),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1190),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1204),
.A2(n_1164),
.B1(n_1225),
.B2(n_1171),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1166),
.B(n_1062),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1225),
.A2(n_947),
.B1(n_944),
.B2(n_928),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1166),
.B(n_1062),
.Y(n_1281)
);

OAI221xp5_ASAP7_75t_L g1282 ( 
.A1(n_1180),
.A2(n_855),
.B1(n_754),
.B2(n_530),
.C(n_537),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1229),
.B(n_1097),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1212),
.B(n_1097),
.C(n_1022),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1216),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1190),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1185),
.B(n_1188),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1189),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1165),
.B(n_1097),
.Y(n_1289)
);

NOR2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1226),
.B(n_1062),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1217),
.B(n_1086),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1186),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1185),
.B(n_1092),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1208),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1208),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1174),
.B(n_1092),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1217),
.B(n_1086),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1191),
.Y(n_1298)
);

AO22x2_ASAP7_75t_L g1299 ( 
.A1(n_1214),
.A2(n_1022),
.B1(n_1092),
.B2(n_868),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1223),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1188),
.B(n_1032),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1195),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1222),
.B(n_1221),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1211),
.B(n_1223),
.Y(n_1304)
);

AO22x2_ASAP7_75t_L g1305 ( 
.A1(n_1214),
.A2(n_907),
.B1(n_932),
.B2(n_615),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1182),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1162),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1189),
.B(n_527),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1203),
.B(n_1206),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1218),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1206),
.B(n_527),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1227),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1213),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1203),
.B(n_1087),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1227),
.B(n_980),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1206),
.B(n_1211),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1231),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1213),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1213),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1232),
.Y(n_1321)
);

AO22x2_ASAP7_75t_L g1322 ( 
.A1(n_1233),
.A2(n_932),
.B1(n_907),
.B2(n_614),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1206),
.B(n_1033),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1205),
.B(n_1226),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1224),
.B(n_981),
.Y(n_1325)
);

BUFx4_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1162),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1158),
.A2(n_1073),
.B(n_1058),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1187),
.B(n_1091),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1156),
.B(n_1034),
.Y(n_1330)
);

AO22x2_ASAP7_75t_L g1331 ( 
.A1(n_1172),
.A2(n_614),
.B1(n_715),
.B2(n_575),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1172),
.A2(n_657),
.B(n_661),
.C(n_638),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1162),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1187),
.B(n_1091),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1220),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1175),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1274),
.A2(n_1158),
.B(n_1169),
.C(n_1219),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1234),
.A2(n_1240),
.B(n_1237),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1234),
.A2(n_1169),
.B(n_1156),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1277),
.A2(n_848),
.B(n_712),
.C(n_713),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1264),
.B(n_1175),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1237),
.A2(n_1181),
.B(n_1167),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1240),
.A2(n_1183),
.B(n_1175),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1261),
.A2(n_1183),
.B(n_1175),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1257),
.B(n_1183),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1261),
.A2(n_1183),
.B(n_1181),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1276),
.A2(n_1167),
.B(n_1058),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1298),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1276),
.A2(n_1059),
.B(n_1038),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1286),
.A2(n_1059),
.B(n_1038),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1243),
.B(n_528),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1252),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_L g1353 ( 
.A(n_1250),
.B(n_594),
.C(n_593),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1282),
.A2(n_603),
.B(n_606),
.C(n_599),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1241),
.B(n_982),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1302),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1286),
.A2(n_848),
.B(n_617),
.C(n_625),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1294),
.A2(n_1060),
.B(n_1054),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1298),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1304),
.B(n_1044),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1238),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1294),
.A2(n_1060),
.B(n_1054),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1269),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1295),
.B(n_984),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1328),
.A2(n_1335),
.B(n_1259),
.Y(n_1365)
);

NAND2x1_ASAP7_75t_L g1366 ( 
.A(n_1273),
.B(n_1066),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1295),
.A2(n_1060),
.B(n_717),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1304),
.B(n_1287),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1321),
.A2(n_734),
.B(n_739),
.C(n_693),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1279),
.B(n_985),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1287),
.B(n_988),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1315),
.A2(n_1060),
.B(n_1066),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1279),
.B(n_992),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1318),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1258),
.A2(n_604),
.B1(n_605),
.B2(n_601),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1273),
.B(n_1039),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1310),
.A2(n_1072),
.B(n_1066),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1242),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1281),
.B(n_995),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1265),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1235),
.A2(n_705),
.B1(n_720),
.B2(n_669),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1267),
.A2(n_705),
.B1(n_720),
.B2(n_669),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1253),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1289),
.A2(n_1072),
.B(n_1066),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1281),
.B(n_997),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1292),
.B(n_998),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1266),
.A2(n_1072),
.B(n_1066),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1249),
.A2(n_777),
.B(n_746),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1283),
.A2(n_818),
.B(n_823),
.C(n_807),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1296),
.A2(n_1072),
.B(n_592),
.Y(n_1390)
);

AO32x1_ASAP7_75t_L g1391 ( 
.A1(n_1269),
.A2(n_1043),
.A3(n_1042),
.B1(n_679),
.B2(n_715),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1311),
.A2(n_854),
.B(n_835),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1317),
.A2(n_1072),
.B(n_592),
.Y(n_1393)
);

INVx6_ASAP7_75t_SL g1394 ( 
.A(n_1245),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1280),
.B(n_534),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1260),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1323),
.B(n_1000),
.Y(n_1397)
);

AND2x6_ASAP7_75t_SL g1398 ( 
.A(n_1275),
.B(n_609),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1323),
.B(n_534),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1265),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1256),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1270),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1301),
.B(n_535),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1270),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1271),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1301),
.B(n_535),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1265),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1244),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1267),
.A2(n_705),
.B1(n_720),
.B2(n_669),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1324),
.A2(n_640),
.B(n_643),
.C(n_630),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1300),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1303),
.A2(n_658),
.B(n_673),
.C(n_654),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1314),
.A2(n_600),
.B(n_580),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1271),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1319),
.A2(n_600),
.B(n_580),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1309),
.A2(n_677),
.B(n_680),
.C(n_676),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1236),
.A2(n_878),
.B(n_859),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1239),
.A2(n_941),
.B(n_899),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1246),
.Y(n_1419)
);

AO22x1_ASAP7_75t_L g1420 ( 
.A1(n_1245),
.A2(n_541),
.B1(n_542),
.B2(n_537),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1320),
.A2(n_652),
.B(n_627),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1330),
.B(n_541),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1330),
.B(n_542),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1293),
.B(n_547),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1293),
.B(n_547),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1278),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1312),
.A2(n_652),
.B(n_627),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1251),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1263),
.A2(n_701),
.B(n_666),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1306),
.A2(n_701),
.B(n_666),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1288),
.B(n_1039),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1254),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1248),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1288),
.A2(n_732),
.B(n_711),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1354),
.A2(n_1332),
.B(n_1334),
.C(n_1329),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1338),
.A2(n_1307),
.B(n_1278),
.Y(n_1436)
);

INVx3_ASAP7_75t_SL g1437 ( 
.A(n_1352),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1352),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1355),
.B(n_1316),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1361),
.B(n_1248),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1353),
.B(n_1313),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1374),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1401),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1395),
.A2(n_1326),
.B1(n_1284),
.B2(n_551),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1356),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1368),
.B(n_1327),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1433),
.B(n_1325),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1378),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1387),
.A2(n_1307),
.B(n_1278),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1368),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1343),
.A2(n_1344),
.B(n_1358),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1411),
.Y(n_1452)
);

BUFx8_ASAP7_75t_SL g1453 ( 
.A(n_1371),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1420),
.B(n_1291),
.Y(n_1454)
);

INVx5_ASAP7_75t_L g1455 ( 
.A(n_1380),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1394),
.Y(n_1456)
);

INVxp67_ASAP7_75t_SL g1457 ( 
.A(n_1346),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1371),
.B(n_1345),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1392),
.A2(n_1290),
.B(n_1333),
.C(n_1308),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1348),
.B(n_1299),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1383),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1380),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1408),
.B(n_1307),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1359),
.B(n_1299),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1375),
.B(n_1305),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1398),
.B(n_1297),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1396),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1386),
.B(n_1262),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1340),
.A2(n_1336),
.B(n_1272),
.C(n_1285),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1394),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1363),
.B(n_1305),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1414),
.B(n_1268),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1402),
.B(n_1247),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1380),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1404),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1412),
.A2(n_569),
.B(n_650),
.C(n_646),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1369),
.A2(n_684),
.B(n_687),
.C(n_681),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1405),
.B(n_1247),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1362),
.A2(n_1255),
.B(n_1331),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1357),
.A2(n_689),
.B(n_694),
.C(n_688),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1364),
.B(n_1322),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1370),
.B(n_1322),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1419),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1360),
.B(n_1331),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1373),
.B(n_550),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1400),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1428),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1403),
.A2(n_567),
.B1(n_581),
.B2(n_555),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1384),
.A2(n_732),
.B(n_711),
.Y(n_1490)
);

AOI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1365),
.A2(n_1046),
.B(n_1045),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1432),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1379),
.B(n_550),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1372),
.A2(n_858),
.B(n_733),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1400),
.Y(n_1495)
);

BUFx2_ASAP7_75t_SL g1496 ( 
.A(n_1407),
.Y(n_1496)
);

OA22x2_ASAP7_75t_L g1497 ( 
.A1(n_1422),
.A2(n_554),
.B1(n_555),
.B2(n_551),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1337),
.A2(n_569),
.B(n_650),
.C(n_646),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1406),
.A2(n_558),
.B1(n_560),
.B2(n_554),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1416),
.A2(n_699),
.B(n_703),
.C(n_696),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1397),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1385),
.Y(n_1502)
);

INVx8_ASAP7_75t_L g1503 ( 
.A(n_1407),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1341),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1410),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1339),
.A2(n_858),
.B(n_733),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1377),
.A2(n_909),
.B(n_896),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1347),
.A2(n_909),
.B(n_896),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1349),
.A2(n_955),
.B(n_948),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1351),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1423),
.B(n_558),
.Y(n_1511)
);

CKINVDCx8_ASAP7_75t_R g1512 ( 
.A(n_1382),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1417),
.B(n_562),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1381),
.A2(n_959),
.B1(n_595),
.B2(n_560),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1350),
.A2(n_955),
.B(n_945),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1399),
.A2(n_563),
.B1(n_929),
.B2(n_579),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1434),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1409),
.A2(n_708),
.B1(n_721),
.B2(n_707),
.C(n_704),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1426),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1418),
.B(n_559),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_SL g1521 ( 
.A(n_1342),
.B(n_710),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1388),
.B(n_1044),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1366),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1431),
.B(n_1044),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1389),
.A2(n_927),
.B(n_761),
.C(n_575),
.Y(n_1525)
);

INVx3_ASAP7_75t_SL g1526 ( 
.A(n_1427),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1429),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1413),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1367),
.A2(n_679),
.B(n_533),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1431),
.B(n_559),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1391),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1415),
.B(n_563),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1421),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1393),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1376),
.B(n_567),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1376),
.B(n_1039),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1452),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1461),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1450),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1455),
.B(n_1450),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1468),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1445),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1455),
.B(n_1390),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1442),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1463),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1442),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1520),
.B(n_572),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1466),
.A2(n_729),
.B1(n_905),
.B2(n_874),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1450),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1492),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1484),
.Y(n_1551)
);

BUFx12f_ASAP7_75t_L g1552 ( 
.A(n_1510),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1457),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1476),
.B(n_1430),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1475),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1501),
.B(n_722),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1531),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1480),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1463),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1437),
.Y(n_1560)
);

BUFx8_ASAP7_75t_L g1561 ( 
.A(n_1448),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1460),
.B(n_724),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1455),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1488),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1473),
.Y(n_1565)
);

BUFx2_ASAP7_75t_R g1566 ( 
.A(n_1453),
.Y(n_1566)
);

INVx5_ASAP7_75t_L g1567 ( 
.A(n_1485),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1473),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1465),
.B(n_747),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1469),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1439),
.B(n_729),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1472),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1443),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1463),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1438),
.Y(n_1575)
);

BUFx2_ASAP7_75t_R g1576 ( 
.A(n_1512),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1438),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1504),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1487),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1496),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1521),
.A2(n_573),
.B1(n_576),
.B2(n_572),
.Y(n_1581)
);

BUFx12f_ASAP7_75t_L g1582 ( 
.A(n_1438),
.Y(n_1582)
);

BUFx12f_ASAP7_75t_L g1583 ( 
.A(n_1487),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1503),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1474),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1503),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1446),
.B(n_1458),
.Y(n_1587)
);

INVx8_ASAP7_75t_L g1588 ( 
.A(n_1446),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1479),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1462),
.B(n_573),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1440),
.B(n_729),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1536),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1456),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1495),
.Y(n_1594)
);

BUFx2_ASAP7_75t_SL g1595 ( 
.A(n_1471),
.Y(n_1595)
);

CKINVDCx6p67_ASAP7_75t_R g1596 ( 
.A(n_1441),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1447),
.B(n_874),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1536),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1519),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1502),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1464),
.B(n_1039),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1467),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1485),
.B(n_1042),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1454),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1482),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1483),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1435),
.B(n_753),
.Y(n_1607)
);

BUFx2_ASAP7_75t_SL g1608 ( 
.A(n_1497),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1436),
.B(n_1043),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1444),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1523),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1491),
.Y(n_1612)
);

INVx5_ASAP7_75t_L g1613 ( 
.A(n_1526),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1459),
.Y(n_1614)
);

INVx5_ASAP7_75t_L g1615 ( 
.A(n_1470),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1528),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1486),
.B(n_874),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1522),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1533),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1538),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1616),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1547),
.A2(n_1481),
.B(n_1498),
.C(n_1477),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1543),
.A2(n_1451),
.B(n_1494),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1553),
.A2(n_1508),
.B(n_1449),
.Y(n_1624)
);

CKINVDCx20_ASAP7_75t_R g1625 ( 
.A(n_1561),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1613),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1607),
.A2(n_1513),
.B(n_1532),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1558),
.A2(n_1515),
.B(n_1509),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1541),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1598),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1564),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1619),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1547),
.A2(n_1506),
.B(n_1500),
.Y(n_1633)
);

BUFx10_ASAP7_75t_L g1634 ( 
.A(n_1560),
.Y(n_1634)
);

BUFx2_ASAP7_75t_R g1635 ( 
.A(n_1610),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1607),
.A2(n_1505),
.B(n_1478),
.C(n_1525),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_SL g1637 ( 
.A1(n_1580),
.A2(n_1575),
.B(n_1553),
.C(n_1581),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1543),
.A2(n_1534),
.B(n_1527),
.Y(n_1638)
);

NAND2x1_ASAP7_75t_L g1639 ( 
.A(n_1577),
.B(n_1517),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1554),
.A2(n_1507),
.B(n_1490),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1554),
.A2(n_1529),
.B(n_1524),
.Y(n_1641)
);

CKINVDCx6p67_ASAP7_75t_R g1642 ( 
.A(n_1552),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1551),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1590),
.A2(n_1499),
.B(n_1489),
.C(n_1516),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1613),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1606),
.B(n_1605),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1615),
.B(n_1535),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1548),
.A2(n_1518),
.B1(n_905),
.B2(n_769),
.Y(n_1649)
);

BUFx4f_ASAP7_75t_L g1650 ( 
.A(n_1540),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1583),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1582),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1572),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1598),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1548),
.A2(n_905),
.B1(n_769),
.B2(n_780),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1557),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1585),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1589),
.B(n_1511),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1590),
.A2(n_1514),
.B(n_1493),
.C(n_1530),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1555),
.B(n_756),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1550),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1596),
.A2(n_579),
.B1(n_581),
.B2(n_576),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1537),
.B(n_757),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1587),
.B(n_762),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1618),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1570),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1544),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1614),
.A2(n_766),
.B(n_763),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1557),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1587),
.B(n_775),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1578),
.Y(n_1672)
);

AOI22x1_ASAP7_75t_L g1673 ( 
.A1(n_1577),
.A2(n_583),
.B1(n_587),
.B2(n_582),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1613),
.B(n_761),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1612),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1618),
.Y(n_1676)
);

AO31x2_ASAP7_75t_L g1677 ( 
.A1(n_1542),
.A2(n_1391),
.A3(n_723),
.B(n_843),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1625),
.A2(n_1608),
.B1(n_1615),
.B2(n_1567),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1621),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1621),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1657),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1632),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1632),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1620),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1670),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1639),
.Y(n_1687)
);

BUFx10_ASAP7_75t_L g1688 ( 
.A(n_1668),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1657),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1670),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1638),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1631),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1643),
.B(n_1618),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1627),
.A2(n_1615),
.B(n_1597),
.Y(n_1694)
);

AOI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1648),
.A2(n_1569),
.B(n_1562),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1654),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1672),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1675),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1658),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1676),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1630),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1644),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1675),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1618),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1667),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1626),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1677),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1626),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1669),
.A2(n_1567),
.B1(n_1633),
.B2(n_1604),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1666),
.B(n_1559),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1647),
.Y(n_1714)
);

AO21x1_ASAP7_75t_SL g1715 ( 
.A1(n_1637),
.A2(n_1569),
.B(n_1562),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1666),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1622),
.A2(n_1576),
.B1(n_1580),
.B2(n_1567),
.Y(n_1717)
);

AO21x1_ASAP7_75t_L g1718 ( 
.A1(n_1645),
.A2(n_1556),
.B(n_796),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1646),
.Y(n_1719)
);

CKINVDCx11_ASAP7_75t_R g1720 ( 
.A(n_1625),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1623),
.A2(n_1592),
.B(n_1545),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1646),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1641),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1622),
.A2(n_1617),
.B(n_1591),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1653),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1677),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1664),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_R g1728 ( 
.A(n_1693),
.B(n_1651),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1717),
.A2(n_1656),
.B1(n_1649),
.B2(n_1567),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1653),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1700),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1681),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1689),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1682),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1720),
.B(n_1651),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1703),
.B(n_1637),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1682),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1679),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1714),
.B(n_1661),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1715),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1679),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1679),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_1688),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1684),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_R g1745 ( 
.A(n_1694),
.B(n_1573),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1714),
.B(n_1659),
.Y(n_1746)
);

OAI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1717),
.A2(n_1656),
.B1(n_1600),
.B2(n_1649),
.C1(n_1565),
.C2(n_1665),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1718),
.A2(n_1671),
.B1(n_1571),
.B2(n_1600),
.Y(n_1748)
);

CKINVDCx16_ASAP7_75t_R g1749 ( 
.A(n_1688),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_SL g1750 ( 
.A(n_1724),
.B(n_1663),
.C(n_1660),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1704),
.B(n_1713),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1680),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1642),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1719),
.B(n_1652),
.Y(n_1754)
);

AO32x2_ASAP7_75t_L g1755 ( 
.A1(n_1706),
.A2(n_1678),
.A3(n_1705),
.B1(n_1716),
.B2(n_1683),
.Y(n_1755)
);

NAND2xp33_ASAP7_75t_R g1756 ( 
.A(n_1694),
.B(n_1579),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1688),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1719),
.B(n_1634),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1680),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1719),
.B(n_1652),
.Y(n_1760)
);

CKINVDCx16_ASAP7_75t_R g1761 ( 
.A(n_1688),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1718),
.A2(n_1724),
.B1(n_1712),
.B2(n_1715),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1710),
.B(n_1630),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1703),
.B(n_1624),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1711),
.A2(n_1628),
.B(n_1636),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1698),
.B(n_1628),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1716),
.B(n_1634),
.Y(n_1767)
);

NAND2xp33_ASAP7_75t_R g1768 ( 
.A(n_1696),
.B(n_1566),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1680),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1701),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1710),
.B(n_1630),
.Y(n_1771)
);

AO31x2_ASAP7_75t_L g1772 ( 
.A1(n_1691),
.A2(n_1636),
.A3(n_1568),
.B(n_1556),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1683),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1684),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_R g1775 ( 
.A(n_1696),
.B(n_1566),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1686),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_R g1777 ( 
.A(n_1710),
.B(n_1561),
.Y(n_1777)
);

NOR2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1687),
.B(n_1602),
.Y(n_1778)
);

BUFx4f_ASAP7_75t_SL g1779 ( 
.A(n_1701),
.Y(n_1779)
);

BUFx4f_ASAP7_75t_SL g1780 ( 
.A(n_1701),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1738),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1764),
.B(n_1698),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1698),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1734),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1778),
.B(n_1706),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1742),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1750),
.A2(n_1678),
.B1(n_1611),
.B2(n_1707),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1758),
.B(n_1635),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1752),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1764),
.B(n_1705),
.Y(n_1792)
);

AO21x2_ASAP7_75t_L g1793 ( 
.A1(n_1765),
.A2(n_1709),
.B(n_1708),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1759),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1737),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1744),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1732),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1733),
.B(n_1699),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1730),
.B(n_1722),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1730),
.B(n_1722),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1767),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1755),
.B(n_1722),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1755),
.B(n_1722),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1755),
.B(n_1727),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1739),
.B(n_1686),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1736),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1774),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1754),
.B(n_1706),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1773),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1776),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1746),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1786),
.B(n_1749),
.Y(n_1813)
);

AO31x2_ASAP7_75t_L g1814 ( 
.A1(n_1784),
.A2(n_1736),
.A3(n_1795),
.B(n_1787),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1807),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1796),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1805),
.A2(n_1750),
.B1(n_1762),
.B2(n_1748),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1789),
.A2(n_1762),
.B1(n_1748),
.B2(n_1740),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1803),
.A2(n_1766),
.B(n_1765),
.Y(n_1819)
);

O2A1O1Ixp5_ASAP7_75t_L g1820 ( 
.A1(n_1803),
.A2(n_1747),
.B(n_1766),
.C(n_1760),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1809),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1796),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1809),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1808),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1804),
.A2(n_1747),
.B(n_1740),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1808),
.Y(n_1826)
);

AOI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1804),
.A2(n_1745),
.B(n_800),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1812),
.B(n_1692),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1811),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1811),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1782),
.A2(n_1711),
.B(n_1723),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1784),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1795),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1797),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1805),
.A2(n_1756),
.B1(n_1775),
.B2(n_1768),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1798),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1806),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1806),
.Y(n_1838)
);

INVx4_ASAP7_75t_R g1839 ( 
.A(n_1785),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1812),
.A2(n_1729),
.B1(n_1707),
.B2(n_1702),
.Y(n_1840)
);

OR2x6_ASAP7_75t_L g1841 ( 
.A(n_1786),
.B(n_1711),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1792),
.Y(n_1842)
);

CKINVDCx14_ASAP7_75t_R g1843 ( 
.A(n_1790),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1837),
.B(n_1838),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1821),
.B(n_1799),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1826),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1815),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1829),
.Y(n_1848)
);

NOR3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1818),
.B(n_1728),
.C(n_1761),
.Y(n_1849)
);

AO21x2_ASAP7_75t_L g1850 ( 
.A1(n_1825),
.A2(n_1792),
.B(n_1782),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1821),
.B(n_1799),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1823),
.B(n_1800),
.Y(n_1852)
);

INVxp67_ASAP7_75t_SL g1853 ( 
.A(n_1835),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1836),
.B(n_1783),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1830),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1841),
.B(n_1786),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1842),
.B(n_1783),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1817),
.A2(n_1793),
.B1(n_1787),
.B2(n_1788),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1832),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1833),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1828),
.B(n_1785),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1827),
.A2(n_1793),
.B1(n_1787),
.B2(n_1788),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1839),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1819),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1834),
.B(n_1802),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1814),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1816),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1843),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1841),
.Y(n_1869)
);

AND3x1_ASAP7_75t_L g1870 ( 
.A(n_1825),
.B(n_1753),
.C(n_1800),
.Y(n_1870)
);

AO21x2_ASAP7_75t_L g1871 ( 
.A1(n_1831),
.A2(n_1793),
.B(n_1695),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1814),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1814),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1822),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1818),
.B(n_1699),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1827),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1868),
.Y(n_1877)
);

AND2x4_ASAP7_75t_SL g1878 ( 
.A(n_1863),
.B(n_1743),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_R g1879 ( 
.A(n_1863),
.B(n_1847),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1865),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1870),
.B(n_1823),
.Y(n_1881)
);

NAND4xp25_ASAP7_75t_L g1882 ( 
.A(n_1865),
.B(n_1820),
.C(n_1813),
.D(n_1831),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1875),
.B(n_1824),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1850),
.B(n_1840),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1841),
.Y(n_1885)
);

INVxp67_ASAP7_75t_SL g1886 ( 
.A(n_1864),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1845),
.B(n_1809),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1853),
.A2(n_1793),
.B1(n_1820),
.B2(n_1788),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1844),
.B(n_1692),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1844),
.B(n_1781),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1850),
.B(n_1809),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1873),
.Y(n_1892)
);

OR2x6_ASAP7_75t_L g1893 ( 
.A(n_1876),
.B(n_1674),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1851),
.B(n_1786),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1846),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1848),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1851),
.B(n_1754),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_SL g1898 ( 
.A(n_1869),
.B(n_1576),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1855),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1859),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1850),
.B(n_1760),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1854),
.B(n_1702),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1852),
.B(n_1757),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1864),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1873),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1849),
.B(n_1763),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1871),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1877),
.B(n_1852),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1893),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1880),
.B(n_1860),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1893),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1878),
.B(n_1856),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1896),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1899),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1899),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1895),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1893),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1878),
.B(n_1856),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1902),
.B(n_1857),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1900),
.Y(n_1920)
);

OAI22xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1884),
.A2(n_1872),
.B1(n_1866),
.B2(n_1869),
.Y(n_1921)
);

AOI211x1_ASAP7_75t_SL g1922 ( 
.A1(n_1882),
.A2(n_1864),
.B(n_1872),
.C(n_1866),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1886),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1883),
.B(n_1857),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1892),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1879),
.B(n_1864),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1889),
.B(n_1861),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1892),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1889),
.B(n_1861),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1890),
.B(n_1867),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1905),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1905),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1890),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1897),
.B(n_1856),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1897),
.B(n_1869),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1901),
.B(n_1874),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1904),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1885),
.B(n_1871),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1907),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1906),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1907),
.B(n_1858),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1881),
.B(n_1735),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1888),
.B(n_1871),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1881),
.B(n_1862),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1885),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1893),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1891),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1887),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1887),
.B(n_723),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1903),
.B(n_1777),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1903),
.B(n_1763),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1912),
.B(n_1894),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1939),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1908),
.B(n_1937),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1942),
.B(n_1894),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1949),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1912),
.B(n_1906),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1949),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1918),
.B(n_1934),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1918),
.B(n_1906),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1914),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1915),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1945),
.B(n_1898),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1940),
.B(n_1595),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1922),
.A2(n_1674),
.B1(n_845),
.B2(n_881),
.C(n_843),
.Y(n_1965)
);

NOR2xp67_ASAP7_75t_L g1966 ( 
.A(n_1923),
.B(n_1),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1943),
.A2(n_1944),
.B1(n_1938),
.B2(n_1941),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1910),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1926),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1951),
.B(n_1687),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1923),
.B(n_776),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1948),
.B(n_1950),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1935),
.B(n_1546),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1938),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1935),
.B(n_1687),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1910),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1924),
.B(n_802),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1925),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1919),
.B(n_1770),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1927),
.B(n_805),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_SL g1981 ( 
.A(n_1913),
.B(n_1586),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1928),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1931),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1926),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1947),
.B(n_1929),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1916),
.B(n_1771),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1943),
.A2(n_845),
.B1(n_881),
.B2(n_780),
.Y(n_1987)
);

INVxp33_ASAP7_75t_SL g1988 ( 
.A(n_1932),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1930),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1936),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1920),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1933),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1941),
.B(n_816),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1921),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1909),
.B(n_1911),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1917),
.B(n_1687),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1946),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1922),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1921),
.B(n_824),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1942),
.B(n_1771),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1938),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1939),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1908),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1908),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1908),
.B(n_828),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1942),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1939),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_1942),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1908),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1908),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1937),
.B(n_1586),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1939),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1938),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1942),
.B(n_1725),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1942),
.B(n_1725),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_2006),
.B(n_1593),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_2003),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2009),
.B(n_2004),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_2010),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1989),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2009),
.B(n_833),
.Y(n_2021)
);

INVxp33_ASAP7_75t_SL g2022 ( 
.A(n_2008),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1989),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1989),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1990),
.B(n_836),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2005),
.B(n_837),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_1983),
.B(n_839),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1980),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1977),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1966),
.B(n_856),
.Y(n_2030)
);

HB1xp67_ASAP7_75t_L g2031 ( 
.A(n_1972),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_1972),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1963),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1971),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1988),
.B(n_860),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1988),
.B(n_877),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1994),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1955),
.B(n_1593),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1983),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_L g2040 ( 
.A(n_1974),
.B(n_879),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1959),
.B(n_1593),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1953),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1974),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_1969),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2002),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1985),
.B(n_890),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2007),
.Y(n_2047)
);

OAI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_1967),
.A2(n_1673),
.B1(n_900),
.B2(n_906),
.C(n_895),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1968),
.B(n_893),
.Y(n_2049)
);

NOR2x1_ASAP7_75t_L g2050 ( 
.A(n_2001),
.B(n_912),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1963),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2012),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1954),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_1984),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1961),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1962),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1976),
.B(n_934),
.Y(n_2057)
);

INVxp67_ASAP7_75t_SL g2058 ( 
.A(n_1998),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1955),
.B(n_946),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1992),
.B(n_956),
.Y(n_2060)
);

AND2x4_ASAP7_75t_SL g2061 ( 
.A(n_1959),
.B(n_1952),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1952),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1952),
.B(n_960),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2001),
.B(n_582),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1978),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1982),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_2013),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2013),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1957),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_1991),
.B(n_1),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1957),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1999),
.Y(n_2072)
);

NAND3xp33_ASAP7_75t_SL g2073 ( 
.A(n_1967),
.B(n_587),
.C(n_583),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1960),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_L g2075 ( 
.A(n_1987),
.B(n_1965),
.C(n_1993),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1960),
.B(n_1706),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1964),
.B(n_595),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1956),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1964),
.Y(n_2079)
);

INVxp67_ASAP7_75t_L g2080 ( 
.A(n_1981),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1986),
.B(n_598),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2000),
.B(n_1979),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2014),
.B(n_1725),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2014),
.B(n_1725),
.Y(n_2084)
);

AOI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1987),
.A2(n_898),
.B1(n_901),
.B2(n_598),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_1996),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_SL g2087 ( 
.A(n_1973),
.B(n_898),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1958),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1995),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2015),
.B(n_1584),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2015),
.B(n_1584),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1973),
.B(n_2011),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1975),
.B(n_901),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_1973),
.B(n_2),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_1995),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1997),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1975),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1970),
.B(n_902),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1997),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1996),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1970),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2009),
.B(n_902),
.Y(n_2102)
);

OAI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_2022),
.A2(n_2054),
.B(n_2044),
.Y(n_2103)
);

NAND4xp25_ASAP7_75t_L g2104 ( 
.A(n_2032),
.B(n_1563),
.C(n_910),
.D(n_913),
.Y(n_2104)
);

OAI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_2058),
.A2(n_913),
.B1(n_914),
.B2(n_910),
.C(n_908),
.Y(n_2105)
);

OAI21xp5_ASAP7_75t_SL g2106 ( 
.A1(n_2044),
.A2(n_2054),
.B(n_2031),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2037),
.A2(n_919),
.B1(n_920),
.B2(n_908),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2019),
.Y(n_2108)
);

OAI21xp33_ASAP7_75t_L g2109 ( 
.A1(n_2061),
.A2(n_919),
.B(n_914),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2043),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2033),
.A2(n_1780),
.B1(n_1779),
.B2(n_921),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2062),
.B(n_920),
.Y(n_2112)
);

OAI221xp5_ASAP7_75t_L g2113 ( 
.A1(n_2095),
.A2(n_929),
.B1(n_930),
.B2(n_923),
.C(n_921),
.Y(n_2113)
);

O2A1O1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_2073),
.A2(n_2048),
.B(n_2067),
.C(n_2051),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_2087),
.A2(n_930),
.B1(n_940),
.B2(n_923),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2018),
.Y(n_2116)
);

AOI332xp33_ASAP7_75t_L g2117 ( 
.A1(n_2020),
.A2(n_949),
.A3(n_940),
.B1(n_959),
.B2(n_953),
.B3(n_943),
.C1(n_936),
.C2(n_11),
.Y(n_2117)
);

OAI32xp33_ASAP7_75t_L g2118 ( 
.A1(n_2039),
.A2(n_949),
.A3(n_953),
.B1(n_943),
.B2(n_936),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2089),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2082),
.B(n_610),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2087),
.A2(n_1791),
.B1(n_1794),
.B2(n_1781),
.Y(n_2121)
);

OAI21xp5_ASAP7_75t_SL g2122 ( 
.A1(n_2017),
.A2(n_1695),
.B(n_1701),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2027),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2069),
.B(n_616),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2059),
.B(n_3),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2072),
.A2(n_1791),
.B1(n_1794),
.B2(n_1781),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2023),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2098),
.B(n_626),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2071),
.B(n_629),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2094),
.Y(n_2130)
);

OAI21xp33_ASAP7_75t_L g2131 ( 
.A1(n_2074),
.A2(n_645),
.B(n_631),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2024),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2086),
.B(n_647),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_SL g2134 ( 
.A1(n_2053),
.A2(n_649),
.B1(n_651),
.B2(n_648),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2080),
.A2(n_1780),
.B1(n_1779),
.B2(n_1791),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2093),
.B(n_653),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_2070),
.B(n_655),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2100),
.B(n_664),
.Y(n_2138)
);

A2O1A1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_2046),
.A2(n_668),
.B(n_670),
.C(n_665),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2025),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2041),
.B(n_671),
.Y(n_2141)
);

OAI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_2016),
.A2(n_674),
.B(n_672),
.Y(n_2142)
);

AOI21xp33_ASAP7_75t_SL g2143 ( 
.A1(n_2102),
.A2(n_3),
.B(n_4),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2097),
.B(n_678),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2038),
.A2(n_683),
.B(n_682),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2079),
.A2(n_1801),
.B1(n_1810),
.B2(n_1794),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2101),
.B(n_686),
.Y(n_2147)
);

OAI21xp5_ASAP7_75t_SL g2148 ( 
.A1(n_2092),
.A2(n_2101),
.B(n_2076),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2090),
.B(n_692),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2063),
.Y(n_2150)
);

XNOR2x1_ASAP7_75t_L g2151 ( 
.A(n_2072),
.B(n_695),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2081),
.A2(n_1810),
.B1(n_1801),
.B2(n_698),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2092),
.A2(n_1810),
.B1(n_1801),
.B2(n_706),
.Y(n_2153)
);

INVxp67_ASAP7_75t_L g2154 ( 
.A(n_2040),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_2068),
.Y(n_2155)
);

O2A1O1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_2035),
.A2(n_927),
.B(n_709),
.C(n_719),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2091),
.B(n_697),
.Y(n_2157)
);

AOI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_2034),
.A2(n_2029),
.B1(n_2028),
.B2(n_2096),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2099),
.A2(n_735),
.B1(n_744),
.B2(n_743),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2026),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2036),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2077),
.A2(n_748),
.B1(n_755),
.B2(n_745),
.Y(n_2162)
);

AOI21xp33_ASAP7_75t_SL g2163 ( 
.A1(n_2078),
.A2(n_4),
.B(n_5),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_2021),
.B(n_760),
.Y(n_2164)
);

O2A1O1Ixp33_ASAP7_75t_L g2165 ( 
.A1(n_2042),
.A2(n_768),
.B(n_772),
.C(n_767),
.Y(n_2165)
);

OAI22x1_ASAP7_75t_L g2166 ( 
.A1(n_2085),
.A2(n_1563),
.B1(n_781),
.B2(n_782),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2030),
.Y(n_2167)
);

OAI21xp33_ASAP7_75t_L g2168 ( 
.A1(n_2088),
.A2(n_783),
.B(n_773),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_2064),
.B(n_6),
.Y(n_2169)
);

OAI221xp5_ASAP7_75t_L g2170 ( 
.A1(n_2085),
.A2(n_789),
.B1(n_794),
.B2(n_788),
.C(n_787),
.Y(n_2170)
);

NAND3xp33_ASAP7_75t_L g2171 ( 
.A(n_2045),
.B(n_808),
.C(n_797),
.Y(n_2171)
);

INVx1_ASAP7_75t_SL g2172 ( 
.A(n_2060),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2047),
.B(n_810),
.Y(n_2173)
);

AOI211x1_ASAP7_75t_L g2174 ( 
.A1(n_2052),
.A2(n_1723),
.B(n_8),
.C(n_6),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2049),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2065),
.B(n_813),
.Y(n_2176)
);

AOI211xp5_ASAP7_75t_SL g2177 ( 
.A1(n_2066),
.A2(n_2056),
.B(n_2055),
.C(n_2057),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2050),
.B(n_819),
.Y(n_2178)
);

AOI222xp33_ASAP7_75t_L g2179 ( 
.A1(n_2075),
.A2(n_827),
.B1(n_829),
.B2(n_832),
.C1(n_830),
.C2(n_826),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2075),
.Y(n_2180)
);

OAI21xp33_ASAP7_75t_SL g2181 ( 
.A1(n_2083),
.A2(n_2084),
.B(n_1721),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2061),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2061),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2031),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2022),
.B(n_838),
.Y(n_2185)
);

OAI221xp5_ASAP7_75t_SL g2186 ( 
.A1(n_2044),
.A2(n_1691),
.B1(n_1592),
.B2(n_1545),
.C(n_1697),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_2022),
.B(n_841),
.Y(n_2187)
);

OAI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_2044),
.A2(n_846),
.B1(n_847),
.B2(n_842),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2031),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2022),
.B(n_849),
.Y(n_2190)
);

NAND2xp33_ASAP7_75t_L g2191 ( 
.A(n_2044),
.B(n_850),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2031),
.Y(n_2192)
);

OAI32xp33_ASAP7_75t_L g2193 ( 
.A1(n_2044),
.A2(n_861),
.A3(n_862),
.B1(n_857),
.B2(n_851),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2037),
.A2(n_869),
.B1(n_870),
.B2(n_866),
.C(n_863),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_2022),
.B(n_871),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2044),
.A2(n_880),
.B(n_872),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2031),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2031),
.Y(n_2198)
);

AOI222xp33_ASAP7_75t_L g2199 ( 
.A1(n_2037),
.A2(n_884),
.B1(n_886),
.B2(n_891),
.C1(n_889),
.C2(n_885),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2061),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2031),
.B(n_897),
.Y(n_2201)
);

AOI21xp33_ASAP7_75t_SL g2202 ( 
.A1(n_2022),
.A2(n_7),
.B(n_8),
.Y(n_2202)
);

OAI21xp33_ASAP7_75t_SL g2203 ( 
.A1(n_2058),
.A2(n_1721),
.B(n_7),
.Y(n_2203)
);

NOR3xp33_ASAP7_75t_L g2204 ( 
.A(n_2073),
.B(n_539),
.C(n_528),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2031),
.Y(n_2205)
);

OAI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_2022),
.A2(n_1650),
.B(n_1574),
.Y(n_2206)
);

NAND3xp33_ASAP7_75t_L g2207 ( 
.A(n_2031),
.B(n_1594),
.C(n_543),
.Y(n_2207)
);

INVx1_ASAP7_75t_SL g2208 ( 
.A(n_2044),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2031),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2031),
.Y(n_2210)
);

AOI21xp33_ASAP7_75t_L g2211 ( 
.A1(n_2044),
.A2(n_543),
.B(n_539),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2022),
.B(n_11),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_SL g2213 ( 
.A1(n_2058),
.A2(n_1701),
.B1(n_1594),
.B2(n_749),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2031),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2031),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2031),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2031),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2031),
.Y(n_2218)
);

OAI21xp33_ASAP7_75t_L g2219 ( 
.A1(n_2022),
.A2(n_1594),
.B(n_1691),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2031),
.B(n_12),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2044),
.A2(n_1650),
.B1(n_1701),
.B2(n_1594),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2032),
.B(n_13),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_2022),
.B(n_1630),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2031),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2031),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2022),
.B(n_13),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2022),
.B(n_14),
.Y(n_2227)
);

OAI31xp33_ASAP7_75t_L g2228 ( 
.A1(n_2037),
.A2(n_1603),
.A3(n_1540),
.B(n_612),
.Y(n_2228)
);

NOR3xp33_ASAP7_75t_SL g2229 ( 
.A(n_2018),
.B(n_553),
.C(n_546),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2037),
.A2(n_749),
.B1(n_831),
.B2(n_710),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2031),
.Y(n_2231)
);

INVx2_ASAP7_75t_SL g2232 ( 
.A(n_2061),
.Y(n_2232)
);

AOI21xp33_ASAP7_75t_SL g2233 ( 
.A1(n_2022),
.A2(n_15),
.B(n_16),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2031),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2031),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2031),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2022),
.B(n_16),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2022),
.B(n_17),
.Y(n_2238)
);

NOR2x1_ASAP7_75t_L g2239 ( 
.A(n_2044),
.B(n_17),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_2044),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2031),
.Y(n_2241)
);

OAI21xp33_ASAP7_75t_SL g2242 ( 
.A1(n_2058),
.A2(n_19),
.B(n_20),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2031),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_2061),
.B(n_19),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_2032),
.B(n_21),
.Y(n_2245)
);

OAI21xp33_ASAP7_75t_L g2246 ( 
.A1(n_2022),
.A2(n_1690),
.B(n_1685),
.Y(n_2246)
);

AOI32xp33_ASAP7_75t_L g2247 ( 
.A1(n_2044),
.A2(n_1603),
.A3(n_1772),
.B1(n_1697),
.B2(n_1683),
.Y(n_2247)
);

AOI21xp33_ASAP7_75t_SL g2248 ( 
.A1(n_2022),
.A2(n_21),
.B(n_22),
.Y(n_2248)
);

OAI21xp33_ASAP7_75t_L g2249 ( 
.A1(n_2022),
.A2(n_1690),
.B(n_1685),
.Y(n_2249)
);

INVx3_ASAP7_75t_L g2250 ( 
.A(n_2061),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2022),
.B(n_22),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2031),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2208),
.B(n_23),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2242),
.B(n_23),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2240),
.B(n_24),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2244),
.B(n_25),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2244),
.B(n_26),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_2202),
.B(n_27),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2120),
.B(n_2239),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2239),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2155),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2155),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2220),
.B(n_29),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2174),
.B(n_2233),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2103),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2248),
.B(n_30),
.Y(n_2266)
);

NAND3xp33_ASAP7_75t_SL g2267 ( 
.A(n_2106),
.B(n_553),
.C(n_546),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2201),
.B(n_30),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2110),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2250),
.B(n_2232),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2222),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2115),
.B(n_31),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2245),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2163),
.B(n_32),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_2250),
.B(n_33),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2184),
.B(n_2189),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2182),
.B(n_34),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2125),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2151),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2237),
.B(n_34),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2112),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2212),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2226),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2238),
.B(n_2130),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2123),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2137),
.B(n_35),
.Y(n_2286)
);

INVxp67_ASAP7_75t_SL g2287 ( 
.A(n_2191),
.Y(n_2287)
);

NOR2x1_ASAP7_75t_L g2288 ( 
.A(n_2104),
.B(n_35),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2166),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2227),
.Y(n_2290)
);

OAI31xp33_ASAP7_75t_L g2291 ( 
.A1(n_2180),
.A2(n_642),
.A3(n_690),
.B(n_531),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_2183),
.Y(n_2292)
);

INVxp67_ASAP7_75t_L g2293 ( 
.A(n_2251),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2192),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2197),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2200),
.B(n_37),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2149),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2198),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_2157),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2124),
.B(n_37),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2205),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2129),
.B(n_38),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2209),
.B(n_38),
.Y(n_2303)
);

NAND2x1_ASAP7_75t_L g2304 ( 
.A(n_2210),
.B(n_1655),
.Y(n_2304)
);

NOR2x1_ASAP7_75t_L g2305 ( 
.A(n_2214),
.B(n_39),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2215),
.B(n_39),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2216),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_2141),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2217),
.Y(n_2309)
);

NOR3xp33_ASAP7_75t_L g2310 ( 
.A(n_2114),
.B(n_562),
.C(n_556),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2218),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2203),
.B(n_1655),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2169),
.Y(n_2313)
);

NOR3xp33_ASAP7_75t_L g2314 ( 
.A(n_2105),
.B(n_566),
.C(n_556),
.Y(n_2314)
);

NOR2xp67_ASAP7_75t_L g2315 ( 
.A(n_2224),
.B(n_40),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2199),
.B(n_40),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2196),
.B(n_41),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2179),
.B(n_41),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2225),
.Y(n_2319)
);

CKINVDCx16_ASAP7_75t_R g2320 ( 
.A(n_2158),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2148),
.B(n_42),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2173),
.B(n_42),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2176),
.B(n_43),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_SL g2324 ( 
.A1(n_2177),
.A2(n_43),
.B(n_44),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2139),
.B(n_46),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2143),
.B(n_46),
.Y(n_2326)
);

INVxp67_ASAP7_75t_L g2327 ( 
.A(n_2178),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2231),
.B(n_47),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2204),
.B(n_48),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2140),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2234),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2150),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2161),
.B(n_49),
.Y(n_2333)
);

OAI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2235),
.A2(n_578),
.B(n_566),
.Y(n_2334)
);

INVx1_ASAP7_75t_SL g2335 ( 
.A(n_2185),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2236),
.B(n_49),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2241),
.B(n_50),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2243),
.B(n_50),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2252),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_2187),
.B(n_51),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_2108),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2147),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2138),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2133),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2119),
.B(n_51),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2229),
.B(n_2109),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2116),
.B(n_2188),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2128),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2195),
.B(n_52),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2136),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2190),
.B(n_52),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2144),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2193),
.B(n_53),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2223),
.B(n_53),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2127),
.B(n_54),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2134),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2132),
.B(n_54),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2171),
.B(n_55),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2107),
.B(n_56),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2172),
.B(n_57),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2113),
.B(n_2164),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2175),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2159),
.B(n_58),
.Y(n_2363)
);

INVx1_ASAP7_75t_SL g2364 ( 
.A(n_2211),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2131),
.B(n_59),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_2162),
.B(n_59),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2194),
.B(n_63),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2167),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2156),
.B(n_1655),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2118),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2168),
.B(n_2142),
.Y(n_2371)
);

INVxp67_ASAP7_75t_SL g2372 ( 
.A(n_2292),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2324),
.A2(n_2165),
.B(n_2145),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_2324),
.B(n_2320),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2292),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2315),
.B(n_2154),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_L g2377 ( 
.A(n_2259),
.B(n_2308),
.Y(n_2377)
);

OR2x6_ASAP7_75t_L g2378 ( 
.A(n_2277),
.B(n_2296),
.Y(n_2378)
);

A2O1A1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_2254),
.A2(n_2117),
.B(n_2207),
.C(n_2181),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2270),
.B(n_2213),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2260),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2315),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2265),
.B(n_2206),
.Y(n_2383)
);

OAI211xp5_ASAP7_75t_L g2384 ( 
.A1(n_2261),
.A2(n_2170),
.B(n_2228),
.C(n_2122),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2299),
.A2(n_2152),
.B1(n_2219),
.B2(n_2153),
.Y(n_2385)
);

AOI21xp33_ASAP7_75t_L g2386 ( 
.A1(n_2279),
.A2(n_2160),
.B(n_2230),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2263),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2264),
.B(n_2246),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2305),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2355),
.Y(n_2390)
);

AOI221xp5_ASAP7_75t_SL g2391 ( 
.A1(n_2262),
.A2(n_2221),
.B1(n_2111),
.B2(n_2135),
.C(n_2249),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2345),
.Y(n_2392)
);

INVxp67_ASAP7_75t_SL g2393 ( 
.A(n_2288),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2357),
.Y(n_2394)
);

OR2x2_ASAP7_75t_L g2395 ( 
.A(n_2253),
.B(n_2186),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2306),
.B(n_2121),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_2255),
.B(n_2146),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2306),
.B(n_2247),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2271),
.B(n_2126),
.Y(n_2399)
);

NAND2x1_ASAP7_75t_L g2400 ( 
.A(n_2303),
.B(n_1655),
.Y(n_2400)
);

INVxp67_ASAP7_75t_SL g2401 ( 
.A(n_2284),
.Y(n_2401)
);

NOR2x1_ASAP7_75t_L g2402 ( 
.A(n_2267),
.B(n_63),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2328),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2287),
.B(n_64),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2326),
.Y(n_2405)
);

NOR2x1_ASAP7_75t_L g2406 ( 
.A(n_2338),
.B(n_64),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2256),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2273),
.B(n_65),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_2341),
.B(n_710),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2313),
.Y(n_2410)
);

NOR3xp33_ASAP7_75t_L g2411 ( 
.A(n_2293),
.B(n_589),
.C(n_578),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2257),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2275),
.B(n_2297),
.Y(n_2413)
);

INVxp67_ASAP7_75t_L g2414 ( 
.A(n_2258),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_L g2415 ( 
.A(n_2321),
.B(n_591),
.C(n_589),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2274),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2266),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2281),
.B(n_2278),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2289),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2268),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2335),
.B(n_65),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2351),
.B(n_2332),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2360),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2276),
.B(n_66),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2322),
.Y(n_2425)
);

INVxp67_ASAP7_75t_SL g2426 ( 
.A(n_2323),
.Y(n_2426)
);

NOR2x1_ASAP7_75t_L g2427 ( 
.A(n_2336),
.B(n_68),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2317),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2282),
.B(n_69),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2280),
.B(n_70),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2283),
.B(n_72),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2366),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2294),
.B(n_73),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2290),
.B(n_74),
.Y(n_2434)
);

OR2x2_ASAP7_75t_L g2435 ( 
.A(n_2337),
.B(n_75),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2353),
.B(n_75),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2358),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2364),
.B(n_77),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2295),
.B(n_77),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2298),
.B(n_78),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2301),
.B(n_81),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2307),
.B(n_82),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2316),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2300),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2354),
.B(n_83),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2302),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2286),
.Y(n_2447)
);

AOI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2348),
.A2(n_1598),
.B1(n_1697),
.B2(n_1588),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2309),
.B(n_83),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2330),
.B(n_749),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2371),
.Y(n_2451)
);

NAND2x1p5_ASAP7_75t_L g2452 ( 
.A(n_2368),
.B(n_2356),
.Y(n_2452)
);

NAND3xp33_ASAP7_75t_L g2453 ( 
.A(n_2310),
.B(n_2269),
.C(n_2311),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2350),
.B(n_84),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2304),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2370),
.B(n_86),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2318),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2319),
.B(n_86),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2285),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2340),
.B(n_87),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2331),
.B(n_831),
.Y(n_2461)
);

INVx2_ASAP7_75t_SL g2462 ( 
.A(n_2339),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2346),
.B(n_2333),
.Y(n_2463)
);

OAI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2347),
.A2(n_1685),
.B1(n_1690),
.B2(n_1598),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2272),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2359),
.Y(n_2466)
);

AND2x4_ASAP7_75t_L g2467 ( 
.A(n_2362),
.B(n_89),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2329),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2325),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2327),
.B(n_89),
.Y(n_2470)
);

AOI221xp5_ASAP7_75t_L g2471 ( 
.A1(n_2352),
.A2(n_597),
.B1(n_904),
.B2(n_596),
.C(n_591),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2365),
.B(n_90),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2334),
.B(n_831),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2361),
.B(n_91),
.Y(n_2474)
);

OR2x2_ASAP7_75t_L g2475 ( 
.A(n_2344),
.B(n_91),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2367),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2363),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2349),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2343),
.B(n_2342),
.Y(n_2479)
);

AND3x1_ASAP7_75t_L g2480 ( 
.A(n_2314),
.B(n_92),
.C(n_93),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2369),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2291),
.B(n_92),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2291),
.B(n_2312),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2320),
.B(n_93),
.Y(n_2484)
);

NOR2x1_ASAP7_75t_L g2485 ( 
.A(n_2324),
.B(n_94),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2260),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2324),
.B(n_97),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2260),
.Y(n_2488)
);

OR2x2_ASAP7_75t_L g2489 ( 
.A(n_2292),
.B(n_97),
.Y(n_2489)
);

NOR2x1_ASAP7_75t_L g2490 ( 
.A(n_2292),
.B(n_98),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2260),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2292),
.Y(n_2492)
);

AND2x4_ASAP7_75t_SL g2493 ( 
.A(n_2270),
.B(n_1539),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2324),
.A2(n_597),
.B(n_596),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2260),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2260),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2320),
.B(n_98),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2260),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2320),
.B(n_99),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2260),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2260),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_2292),
.Y(n_2502)
);

INVxp67_ASAP7_75t_SL g2503 ( 
.A(n_2292),
.Y(n_2503)
);

NAND3xp33_ASAP7_75t_L g2504 ( 
.A(n_2324),
.B(n_916),
.C(n_904),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2320),
.B(n_99),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2320),
.B(n_101),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2320),
.B(n_101),
.Y(n_2507)
);

XOR2xp5_ASAP7_75t_L g2508 ( 
.A(n_2320),
.B(n_102),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2320),
.B(n_103),
.Y(n_2509)
);

AOI211xp5_ASAP7_75t_L g2510 ( 
.A1(n_2324),
.A2(n_917),
.B(n_918),
.C(n_916),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2324),
.B(n_104),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2270),
.B(n_104),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2320),
.B(n_105),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2260),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2320),
.B(n_105),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2260),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2270),
.B(n_106),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2270),
.B(n_108),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2320),
.B(n_108),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2260),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2372),
.B(n_109),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2502),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2503),
.Y(n_2523)
);

NOR2x1_ASAP7_75t_L g2524 ( 
.A(n_2375),
.B(n_109),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2378),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2508),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2492),
.B(n_917),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2389),
.B(n_110),
.Y(n_2528)
);

NOR3x1_ASAP7_75t_L g2529 ( 
.A(n_2453),
.B(n_110),
.C(n_113),
.Y(n_2529)
);

NOR2x1p5_ASAP7_75t_L g2530 ( 
.A(n_2401),
.B(n_114),
.Y(n_2530)
);

OAI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2452),
.A2(n_1601),
.B1(n_1549),
.B2(n_1539),
.Y(n_2531)
);

NOR2xp67_ASAP7_75t_L g2532 ( 
.A(n_2512),
.B(n_114),
.Y(n_2532)
);

AOI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2388),
.A2(n_1549),
.B1(n_1539),
.B2(n_1588),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2517),
.B(n_115),
.Y(n_2534)
);

NOR2x1_ASAP7_75t_L g2535 ( 
.A(n_2504),
.B(n_115),
.Y(n_2535)
);

AOI222xp33_ASAP7_75t_L g2536 ( 
.A1(n_2393),
.A2(n_867),
.B1(n_801),
.B2(n_951),
.C1(n_817),
.C2(n_779),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2374),
.B(n_118),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_SL g2538 ( 
.A(n_2518),
.B(n_918),
.Y(n_2538)
);

OAI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2485),
.A2(n_1601),
.B(n_931),
.Y(n_2539)
);

AOI211xp5_ASAP7_75t_SL g2540 ( 
.A1(n_2377),
.A2(n_123),
.B(n_118),
.C(n_119),
.Y(n_2540)
);

NAND3xp33_ASAP7_75t_L g2541 ( 
.A(n_2484),
.B(n_931),
.C(n_924),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2485),
.B(n_119),
.Y(n_2542)
);

NAND2x1_ASAP7_75t_L g2543 ( 
.A(n_2467),
.B(n_125),
.Y(n_2543)
);

OR3x1_ASAP7_75t_L g2544 ( 
.A(n_2381),
.B(n_125),
.C(n_126),
.Y(n_2544)
);

AOI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2380),
.A2(n_935),
.B(n_924),
.Y(n_2545)
);

OAI21xp33_ASAP7_75t_SL g2546 ( 
.A1(n_2462),
.A2(n_128),
.B(n_129),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2490),
.B(n_2451),
.Y(n_2547)
);

NAND3xp33_ASAP7_75t_L g2548 ( 
.A(n_2510),
.B(n_2459),
.C(n_2413),
.Y(n_2548)
);

NOR2xp67_ASAP7_75t_SL g2549 ( 
.A(n_2497),
.B(n_726),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2499),
.Y(n_2550)
);

O2A1O1Ixp5_ASAP7_75t_SL g2551 ( 
.A1(n_2486),
.A2(n_2488),
.B(n_2495),
.C(n_2491),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2467),
.B(n_128),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2487),
.B(n_130),
.Y(n_2553)
);

NOR4xp25_ASAP7_75t_L g2554 ( 
.A(n_2496),
.B(n_133),
.C(n_131),
.D(n_132),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2505),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2511),
.B(n_131),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2424),
.B(n_132),
.Y(n_2557)
);

NOR3xp33_ASAP7_75t_L g2558 ( 
.A(n_2506),
.B(n_938),
.C(n_935),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2507),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2509),
.Y(n_2560)
);

OAI21xp5_ASAP7_75t_SL g2561 ( 
.A1(n_2373),
.A2(n_135),
.B(n_136),
.Y(n_2561)
);

NOR3xp33_ASAP7_75t_L g2562 ( 
.A(n_2513),
.B(n_939),
.C(n_938),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2403),
.B(n_136),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2515),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2383),
.B(n_137),
.Y(n_2565)
);

NOR3x1_ASAP7_75t_L g2566 ( 
.A(n_2418),
.B(n_137),
.C(n_138),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2519),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2433),
.B(n_138),
.Y(n_2568)
);

OAI21xp33_ASAP7_75t_L g2569 ( 
.A1(n_2479),
.A2(n_942),
.B(n_939),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2441),
.B(n_139),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2457),
.A2(n_1549),
.B1(n_1539),
.B2(n_1588),
.Y(n_2571)
);

INVx1_ASAP7_75t_SL g2572 ( 
.A(n_2422),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2410),
.B(n_2402),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2449),
.B(n_139),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_2489),
.B(n_140),
.Y(n_2575)
);

NAND2xp33_ASAP7_75t_L g2576 ( 
.A(n_2379),
.B(n_942),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2390),
.B(n_140),
.Y(n_2577)
);

NAND3xp33_ASAP7_75t_SL g2578 ( 
.A(n_2376),
.B(n_952),
.C(n_950),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2406),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2427),
.Y(n_2580)
);

NOR3xp33_ASAP7_75t_SL g2581 ( 
.A(n_2384),
.B(n_952),
.C(n_950),
.Y(n_2581)
);

NOR2xp67_ASAP7_75t_L g2582 ( 
.A(n_2498),
.B(n_141),
.Y(n_2582)
);

OAI211xp5_ASAP7_75t_L g2583 ( 
.A1(n_2500),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2583)
);

NAND4xp25_ASAP7_75t_L g2584 ( 
.A(n_2391),
.B(n_146),
.C(n_143),
.D(n_144),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2493),
.B(n_147),
.Y(n_2585)
);

OAI21xp33_ASAP7_75t_SL g2586 ( 
.A1(n_2501),
.A2(n_148),
.B(n_150),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2458),
.B(n_150),
.Y(n_2587)
);

AOI21xp33_ASAP7_75t_SL g2588 ( 
.A1(n_2439),
.A2(n_151),
.B(n_152),
.Y(n_2588)
);

NOR2x1_ASAP7_75t_L g2589 ( 
.A(n_2514),
.B(n_151),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2427),
.Y(n_2590)
);

AOI211x1_ASAP7_75t_L g2591 ( 
.A1(n_2516),
.A2(n_157),
.B(n_153),
.C(n_154),
.Y(n_2591)
);

OAI21xp5_ASAP7_75t_SL g2592 ( 
.A1(n_2481),
.A2(n_153),
.B(n_154),
.Y(n_2592)
);

AOI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2404),
.A2(n_957),
.B(n_954),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2394),
.B(n_158),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2382),
.Y(n_2595)
);

INVx2_ASAP7_75t_SL g2596 ( 
.A(n_2440),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2475),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2435),
.Y(n_2598)
);

AOI222xp33_ASAP7_75t_L g2599 ( 
.A1(n_2483),
.A2(n_957),
.B1(n_958),
.B2(n_954),
.C1(n_882),
.C2(n_741),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2494),
.A2(n_958),
.B(n_159),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2392),
.B(n_160),
.Y(n_2601)
);

O2A1O1Ixp33_ASAP7_75t_L g2602 ( 
.A1(n_2473),
.A2(n_163),
.B(n_160),
.C(n_161),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2430),
.B(n_161),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2426),
.Y(n_2604)
);

AOI221x1_ASAP7_75t_L g2605 ( 
.A1(n_2520),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.C(n_167),
.Y(n_2605)
);

AND4x1_ASAP7_75t_L g2606 ( 
.A(n_2402),
.B(n_168),
.C(n_164),
.D(n_167),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2442),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_2421),
.B(n_168),
.Y(n_2608)
);

AOI221xp5_ASAP7_75t_L g2609 ( 
.A1(n_2586),
.A2(n_2463),
.B1(n_2468),
.B2(n_2417),
.C(n_2416),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2582),
.Y(n_2610)
);

AOI221xp5_ASAP7_75t_L g2611 ( 
.A1(n_2573),
.A2(n_2405),
.B1(n_2443),
.B2(n_2428),
.C(n_2478),
.Y(n_2611)
);

A2O1A1Ixp33_ASAP7_75t_L g2612 ( 
.A1(n_2546),
.A2(n_2399),
.B(n_2415),
.C(n_2414),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_R g2613 ( 
.A(n_2522),
.B(n_2445),
.Y(n_2613)
);

OAI211xp5_ASAP7_75t_L g2614 ( 
.A1(n_2523),
.A2(n_2455),
.B(n_2431),
.C(n_2434),
.Y(n_2614)
);

NAND4xp25_ASAP7_75t_L g2615 ( 
.A(n_2584),
.B(n_2386),
.C(n_2385),
.D(n_2387),
.Y(n_2615)
);

OAI211xp5_ASAP7_75t_L g2616 ( 
.A1(n_2604),
.A2(n_2429),
.B(n_2407),
.C(n_2412),
.Y(n_2616)
);

OAI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2572),
.A2(n_2408),
.B1(n_2436),
.B2(n_2454),
.Y(n_2617)
);

OAI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2547),
.A2(n_2400),
.B1(n_2396),
.B2(n_2398),
.C(n_2395),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2544),
.A2(n_2419),
.B1(n_2555),
.B2(n_2550),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2543),
.B(n_2378),
.Y(n_2620)
);

AOI221xp5_ASAP7_75t_SL g2621 ( 
.A1(n_2595),
.A2(n_2423),
.B1(n_2420),
.B2(n_2465),
.C(n_2447),
.Y(n_2621)
);

NAND4xp25_ASAP7_75t_L g2622 ( 
.A(n_2548),
.B(n_2425),
.C(n_2466),
.D(n_2446),
.Y(n_2622)
);

AOI222xp33_ASAP7_75t_L g2623 ( 
.A1(n_2580),
.A2(n_2450),
.B1(n_2432),
.B2(n_2444),
.C1(n_2476),
.C2(n_2477),
.Y(n_2623)
);

AOI211xp5_ASAP7_75t_SL g2624 ( 
.A1(n_2576),
.A2(n_2456),
.B(n_2411),
.C(n_2437),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2540),
.B(n_2474),
.Y(n_2625)
);

INVxp67_ASAP7_75t_SL g2626 ( 
.A(n_2566),
.Y(n_2626)
);

OAI221xp5_ASAP7_75t_L g2627 ( 
.A1(n_2561),
.A2(n_2592),
.B1(n_2539),
.B2(n_2589),
.C(n_2554),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2565),
.B(n_2480),
.Y(n_2628)
);

AOI221xp5_ASAP7_75t_SL g2629 ( 
.A1(n_2545),
.A2(n_2409),
.B1(n_2469),
.B2(n_2397),
.C(n_2461),
.Y(n_2629)
);

AOI221xp5_ASAP7_75t_L g2630 ( 
.A1(n_2593),
.A2(n_2438),
.B1(n_2472),
.B2(n_2460),
.C(n_2482),
.Y(n_2630)
);

AOI222xp33_ASAP7_75t_L g2631 ( 
.A1(n_2590),
.A2(n_2464),
.B1(n_2470),
.B2(n_2471),
.C1(n_2448),
.C2(n_882),
.Y(n_2631)
);

AOI211xp5_ASAP7_75t_L g2632 ( 
.A1(n_2578),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2559),
.A2(n_1549),
.B1(n_1709),
.B2(n_1708),
.Y(n_2633)
);

AOI211x1_ASAP7_75t_SL g2634 ( 
.A1(n_2525),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2634)
);

AOI221xp5_ASAP7_75t_L g2635 ( 
.A1(n_2579),
.A2(n_798),
.B1(n_882),
.B2(n_741),
.C(n_726),
.Y(n_2635)
);

NOR3xp33_ASAP7_75t_L g2636 ( 
.A(n_2526),
.B(n_619),
.C(n_618),
.Y(n_2636)
);

NAND3xp33_ASAP7_75t_SL g2637 ( 
.A(n_2551),
.B(n_628),
.C(n_621),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2606),
.B(n_174),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2530),
.Y(n_2639)
);

OA22x2_ASAP7_75t_L g2640 ( 
.A1(n_2596),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2640)
);

AOI211xp5_ASAP7_75t_SL g2641 ( 
.A1(n_2537),
.A2(n_178),
.B(n_175),
.C(n_177),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2557),
.Y(n_2642)
);

AOI322xp5_ASAP7_75t_L g2643 ( 
.A1(n_2560),
.A2(n_2567),
.A3(n_2564),
.B1(n_2598),
.B2(n_2524),
.C1(n_2597),
.C2(n_2607),
.Y(n_2643)
);

AND2x2_ASAP7_75t_SL g2644 ( 
.A(n_2529),
.B(n_177),
.Y(n_2644)
);

AOI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2521),
.A2(n_178),
.B(n_180),
.Y(n_2645)
);

AND4x2_ASAP7_75t_L g2646 ( 
.A(n_2600),
.B(n_183),
.C(n_181),
.D(n_182),
.Y(n_2646)
);

OAI321xp33_ASAP7_75t_L g2647 ( 
.A1(n_2571),
.A2(n_1609),
.A3(n_882),
.B1(n_741),
.B2(n_798),
.C(n_726),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2534),
.Y(n_2648)
);

NAND4xp25_ASAP7_75t_SL g2649 ( 
.A(n_2599),
.B(n_185),
.C(n_182),
.D(n_184),
.Y(n_2649)
);

NOR4xp25_ASAP7_75t_L g2650 ( 
.A(n_2542),
.B(n_187),
.C(n_184),
.D(n_186),
.Y(n_2650)
);

NAND5xp2_ASAP7_75t_L g2651 ( 
.A(n_2581),
.B(n_189),
.C(n_186),
.D(n_187),
.E(n_192),
.Y(n_2651)
);

OAI31xp33_ASAP7_75t_L g2652 ( 
.A1(n_2541),
.A2(n_196),
.A3(n_192),
.B(n_194),
.Y(n_2652)
);

AOI221xp5_ASAP7_75t_L g2653 ( 
.A1(n_2541),
.A2(n_798),
.B1(n_882),
.B2(n_741),
.C(n_726),
.Y(n_2653)
);

AOI21xp5_ASAP7_75t_SL g2654 ( 
.A1(n_2605),
.A2(n_197),
.B(n_198),
.Y(n_2654)
);

O2A1O1Ixp33_ASAP7_75t_L g2655 ( 
.A1(n_2527),
.A2(n_200),
.B(n_197),
.C(n_199),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2608),
.A2(n_1708),
.B1(n_1726),
.B2(n_1709),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2591),
.B(n_200),
.Y(n_2657)
);

AOI321xp33_ASAP7_75t_L g2658 ( 
.A1(n_2535),
.A2(n_2533),
.A3(n_2577),
.B1(n_2594),
.B2(n_2528),
.C(n_2562),
.Y(n_2658)
);

O2A1O1Ixp33_ASAP7_75t_L g2659 ( 
.A1(n_2602),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_2659)
);

NAND4xp25_ASAP7_75t_SL g2660 ( 
.A(n_2536),
.B(n_205),
.C(n_201),
.D(n_203),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_R g2661 ( 
.A(n_2538),
.B(n_205),
.Y(n_2661)
);

AOI221xp5_ASAP7_75t_L g2662 ( 
.A1(n_2558),
.A2(n_798),
.B1(n_741),
.B2(n_656),
.C(n_660),
.Y(n_2662)
);

NAND2xp33_ASAP7_75t_SL g2663 ( 
.A(n_2552),
.B(n_207),
.Y(n_2663)
);

NAND4xp25_ASAP7_75t_SL g2664 ( 
.A(n_2583),
.B(n_209),
.C(n_207),
.D(n_208),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2588),
.B(n_208),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2568),
.B(n_211),
.Y(n_2666)
);

OAI211xp5_ASAP7_75t_SL g2667 ( 
.A1(n_2611),
.A2(n_2569),
.B(n_2563),
.C(n_2553),
.Y(n_2667)
);

AOI21xp33_ASAP7_75t_L g2668 ( 
.A1(n_2626),
.A2(n_2549),
.B(n_2575),
.Y(n_2668)
);

AOI221xp5_ASAP7_75t_L g2669 ( 
.A1(n_2617),
.A2(n_2601),
.B1(n_2556),
.B2(n_2570),
.C(n_2587),
.Y(n_2669)
);

O2A1O1Ixp5_ASAP7_75t_L g2670 ( 
.A1(n_2616),
.A2(n_2603),
.B(n_2585),
.C(n_2574),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2640),
.Y(n_2671)
);

OAI211xp5_ASAP7_75t_SL g2672 ( 
.A1(n_2643),
.A2(n_2531),
.B(n_2532),
.C(n_214),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2640),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2644),
.B(n_798),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2634),
.B(n_212),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2610),
.Y(n_2676)
);

AND4x1_ASAP7_75t_L g2677 ( 
.A(n_2609),
.B(n_215),
.C(n_212),
.D(n_213),
.Y(n_2677)
);

AOI221xp5_ASAP7_75t_L g2678 ( 
.A1(n_2654),
.A2(n_667),
.B1(n_675),
.B2(n_639),
.C(n_633),
.Y(n_2678)
);

NAND4xp25_ASAP7_75t_L g2679 ( 
.A(n_2619),
.B(n_217),
.C(n_215),
.D(n_216),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2628),
.A2(n_702),
.B1(n_714),
.B2(n_700),
.Y(n_2680)
);

AOI21xp33_ASAP7_75t_L g2681 ( 
.A1(n_2620),
.A2(n_728),
.B(n_716),
.Y(n_2681)
);

OAI311xp33_ASAP7_75t_L g2682 ( 
.A1(n_2615),
.A2(n_219),
.A3(n_216),
.B1(n_218),
.C1(n_220),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2641),
.B(n_220),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2621),
.B(n_740),
.Y(n_2684)
);

AOI22xp5_ASAP7_75t_L g2685 ( 
.A1(n_2639),
.A2(n_752),
.B1(n_765),
.B2(n_742),
.Y(n_2685)
);

OAI211xp5_ASAP7_75t_SL g2686 ( 
.A1(n_2623),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_2686)
);

OAI21xp5_ASAP7_75t_L g2687 ( 
.A1(n_2612),
.A2(n_785),
.B(n_774),
.Y(n_2687)
);

AOI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2618),
.A2(n_791),
.B1(n_792),
.B2(n_790),
.C(n_786),
.Y(n_2688)
);

AOI211xp5_ASAP7_75t_L g2689 ( 
.A1(n_2614),
.A2(n_225),
.B(n_221),
.C(n_223),
.Y(n_2689)
);

NOR3xp33_ASAP7_75t_L g2690 ( 
.A(n_2622),
.B(n_803),
.C(n_793),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2651),
.B(n_225),
.Y(n_2691)
);

AOI222xp33_ASAP7_75t_SL g2692 ( 
.A1(n_2648),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.C1(n_229),
.C2(n_230),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2650),
.B(n_2638),
.Y(n_2693)
);

NAND5xp2_ASAP7_75t_SL g2694 ( 
.A(n_2627),
.B(n_235),
.C(n_231),
.D(n_233),
.E(n_236),
.Y(n_2694)
);

NOR3xp33_ASAP7_75t_L g2695 ( 
.A(n_2637),
.B(n_806),
.C(n_804),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2646),
.Y(n_2696)
);

AND4x1_ASAP7_75t_L g2697 ( 
.A(n_2632),
.B(n_236),
.C(n_231),
.D(n_235),
.Y(n_2697)
);

AOI221xp5_ASAP7_75t_L g2698 ( 
.A1(n_2630),
.A2(n_821),
.B1(n_825),
.B2(n_812),
.C(n_809),
.Y(n_2698)
);

AOI21xp33_ASAP7_75t_SL g2699 ( 
.A1(n_2657),
.A2(n_237),
.B(n_238),
.Y(n_2699)
);

AOI211xp5_ASAP7_75t_L g2700 ( 
.A1(n_2613),
.A2(n_240),
.B(n_237),
.C(n_239),
.Y(n_2700)
);

NAND4xp75_ASAP7_75t_L g2701 ( 
.A(n_2629),
.B(n_241),
.C(n_239),
.D(n_240),
.Y(n_2701)
);

OAI221xp5_ASAP7_75t_L g2702 ( 
.A1(n_2658),
.A2(n_2652),
.B1(n_2636),
.B2(n_2625),
.C(n_2659),
.Y(n_2702)
);

OAI21xp33_ASAP7_75t_L g2703 ( 
.A1(n_2696),
.A2(n_2664),
.B(n_2649),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2671),
.B(n_2660),
.Y(n_2704)
);

AOI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2676),
.A2(n_2672),
.B1(n_2691),
.B2(n_2673),
.Y(n_2705)
);

A2O1A1Ixp33_ASAP7_75t_L g2706 ( 
.A1(n_2678),
.A2(n_2655),
.B(n_2645),
.C(n_2665),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2701),
.B(n_2666),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2667),
.A2(n_2669),
.B1(n_2693),
.B2(n_2642),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2675),
.B(n_2663),
.Y(n_2709)
);

INVxp67_ASAP7_75t_SL g2710 ( 
.A(n_2683),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2697),
.B(n_2624),
.Y(n_2711)
);

INVxp67_ASAP7_75t_L g2712 ( 
.A(n_2692),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2677),
.Y(n_2713)
);

NAND3xp33_ASAP7_75t_SL g2714 ( 
.A(n_2689),
.B(n_2670),
.C(n_2674),
.Y(n_2714)
);

AOI211xp5_ASAP7_75t_L g2715 ( 
.A1(n_2679),
.A2(n_2662),
.B(n_2653),
.C(n_2647),
.Y(n_2715)
);

OAI321xp33_ASAP7_75t_L g2716 ( 
.A1(n_2702),
.A2(n_2635),
.A3(n_2633),
.B1(n_2631),
.B2(n_2656),
.C(n_2661),
.Y(n_2716)
);

AND2x4_ASAP7_75t_L g2717 ( 
.A(n_2684),
.B(n_2690),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2686),
.B(n_241),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2700),
.B(n_2695),
.Y(n_2719)
);

A2O1A1Ixp33_ASAP7_75t_L g2720 ( 
.A1(n_2680),
.A2(n_245),
.B(n_242),
.C(n_244),
.Y(n_2720)
);

NOR3xp33_ASAP7_75t_L g2721 ( 
.A(n_2668),
.B(n_844),
.C(n_834),
.Y(n_2721)
);

OAI21xp33_ASAP7_75t_L g2722 ( 
.A1(n_2688),
.A2(n_853),
.B(n_852),
.Y(n_2722)
);

NOR4xp25_ASAP7_75t_L g2723 ( 
.A(n_2714),
.B(n_2682),
.C(n_2687),
.D(n_2681),
.Y(n_2723)
);

NAND3xp33_ASAP7_75t_L g2724 ( 
.A(n_2708),
.B(n_2698),
.C(n_2699),
.Y(n_2724)
);

NAND3xp33_ASAP7_75t_SL g2725 ( 
.A(n_2705),
.B(n_2685),
.C(n_2694),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2710),
.A2(n_865),
.B1(n_873),
.B2(n_864),
.Y(n_2726)
);

NAND2x1p5_ASAP7_75t_L g2727 ( 
.A(n_2709),
.B(n_242),
.Y(n_2727)
);

NOR3x1_ASAP7_75t_L g2728 ( 
.A(n_2711),
.B(n_2707),
.C(n_2713),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2718),
.Y(n_2729)
);

NOR4xp75_ASAP7_75t_L g2730 ( 
.A(n_2703),
.B(n_247),
.C(n_244),
.D(n_246),
.Y(n_2730)
);

INVx1_ASAP7_75t_SL g2731 ( 
.A(n_2719),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2712),
.B(n_248),
.Y(n_2732)
);

BUFx2_ASAP7_75t_L g2733 ( 
.A(n_2720),
.Y(n_2733)
);

INVx2_ASAP7_75t_SL g2734 ( 
.A(n_2717),
.Y(n_2734)
);

AOI221xp5_ASAP7_75t_L g2735 ( 
.A1(n_2704),
.A2(n_883),
.B1(n_887),
.B2(n_892),
.C(n_251),
.Y(n_2735)
);

A2O1A1Ixp33_ASAP7_75t_L g2736 ( 
.A1(n_2706),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2717),
.B(n_249),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2715),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2721),
.B(n_250),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2734),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2727),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2729),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_R g2743 ( 
.A(n_2725),
.B(n_252),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2731),
.Y(n_2744)
);

OAI21xp5_ASAP7_75t_SL g2745 ( 
.A1(n_2738),
.A2(n_2722),
.B(n_2716),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2723),
.B(n_2728),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2732),
.B(n_253),
.Y(n_2747)
);

BUFx4f_ASAP7_75t_SL g2748 ( 
.A(n_2733),
.Y(n_2748)
);

BUFx6f_ASAP7_75t_L g2749 ( 
.A(n_2737),
.Y(n_2749)
);

NOR3xp33_ASAP7_75t_L g2750 ( 
.A(n_2724),
.B(n_253),
.C(n_254),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2730),
.Y(n_2751)
);

AOI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2739),
.A2(n_254),
.B(n_255),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2736),
.Y(n_2753)
);

CKINVDCx20_ASAP7_75t_R g2754 ( 
.A(n_2726),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2735),
.Y(n_2755)
);

CKINVDCx20_ASAP7_75t_R g2756 ( 
.A(n_2734),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2734),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2729),
.B(n_255),
.Y(n_2758)
);

CKINVDCx20_ASAP7_75t_R g2759 ( 
.A(n_2756),
.Y(n_2759)
);

AOI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2744),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2746),
.A2(n_261),
.B1(n_256),
.B2(n_257),
.Y(n_2761)
);

XOR2xp5_ASAP7_75t_L g2762 ( 
.A(n_2740),
.B(n_261),
.Y(n_2762)
);

AO22x2_ASAP7_75t_L g2763 ( 
.A1(n_2741),
.A2(n_266),
.B1(n_263),
.B2(n_264),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2757),
.B(n_263),
.Y(n_2764)
);

OAI21xp5_ASAP7_75t_L g2765 ( 
.A1(n_2752),
.A2(n_267),
.B(n_268),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2742),
.Y(n_2766)
);

HB1xp67_ASAP7_75t_L g2767 ( 
.A(n_2751),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2748),
.Y(n_2768)
);

OAI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2753),
.A2(n_267),
.B(n_268),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2749),
.Y(n_2770)
);

OAI22x1_ASAP7_75t_L g2771 ( 
.A1(n_2747),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2749),
.Y(n_2772)
);

INVxp67_ASAP7_75t_L g2773 ( 
.A(n_2749),
.Y(n_2773)
);

OA22x2_ASAP7_75t_L g2774 ( 
.A1(n_2745),
.A2(n_2755),
.B1(n_2758),
.B2(n_2743),
.Y(n_2774)
);

OAI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2754),
.A2(n_2750),
.B1(n_1609),
.B2(n_273),
.Y(n_2775)
);

AOI22x1_ASAP7_75t_L g2776 ( 
.A1(n_2744),
.A2(n_273),
.B1(n_270),
.B2(n_272),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2756),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2744),
.A2(n_1609),
.B1(n_276),
.B2(n_274),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2777),
.B(n_2759),
.Y(n_2779)
);

INVx4_ASAP7_75t_L g2780 ( 
.A(n_2770),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2766),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2763),
.Y(n_2782)
);

OR5x1_ASAP7_75t_L g2783 ( 
.A(n_2767),
.B(n_274),
.C(n_275),
.D(n_276),
.E(n_277),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2773),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_2784)
);

AND2x4_ASAP7_75t_SL g2785 ( 
.A(n_2768),
.B(n_278),
.Y(n_2785)
);

NOR3xp33_ASAP7_75t_L g2786 ( 
.A(n_2772),
.B(n_279),
.C(n_280),
.Y(n_2786)
);

OAI22xp5_ASAP7_75t_L g2787 ( 
.A1(n_2761),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2771),
.B(n_281),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2774),
.A2(n_1726),
.B1(n_1640),
.B2(n_1052),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2760),
.A2(n_285),
.B1(n_282),
.B2(n_283),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2764),
.B(n_2762),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2763),
.B(n_285),
.Y(n_2792)
);

XOR2x1_ASAP7_75t_L g2793 ( 
.A(n_2776),
.B(n_286),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2779),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2780),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2792),
.Y(n_2796)
);

INVxp67_ASAP7_75t_SL g2797 ( 
.A(n_2782),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2785),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2793),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2791),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2781),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2783),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2788),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2786),
.Y(n_2804)
);

BUFx2_ASAP7_75t_L g2805 ( 
.A(n_2784),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2787),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2790),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2802),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2794),
.A2(n_2795),
.B1(n_2799),
.B2(n_2797),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2794),
.A2(n_2769),
.B1(n_2765),
.B2(n_2789),
.Y(n_2810)
);

BUFx2_ASAP7_75t_L g2811 ( 
.A(n_2801),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2800),
.A2(n_2775),
.B1(n_2778),
.B2(n_289),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2798),
.B(n_2796),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2803),
.B(n_287),
.Y(n_2814)
);

INVx2_ASAP7_75t_SL g2815 ( 
.A(n_2805),
.Y(n_2815)
);

OAI22xp5_ASAP7_75t_SL g2816 ( 
.A1(n_2804),
.A2(n_291),
.B1(n_288),
.B2(n_289),
.Y(n_2816)
);

XNOR2x1_ASAP7_75t_L g2817 ( 
.A(n_2806),
.B(n_293),
.Y(n_2817)
);

AOI21x1_ASAP7_75t_L g2818 ( 
.A1(n_2807),
.A2(n_294),
.B(n_295),
.Y(n_2818)
);

INVx1_ASAP7_75t_SL g2819 ( 
.A(n_2794),
.Y(n_2819)
);

OAI322xp33_ASAP7_75t_L g2820 ( 
.A1(n_2794),
.A2(n_294),
.A3(n_295),
.B1(n_296),
.B2(n_297),
.C1(n_298),
.C2(n_299),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2794),
.A2(n_296),
.B1(n_300),
.B2(n_302),
.Y(n_2821)
);

OAI22x1_ASAP7_75t_L g2822 ( 
.A1(n_2794),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_2822)
);

OAI22xp5_ASAP7_75t_SL g2823 ( 
.A1(n_2794),
.A2(n_303),
.B1(n_305),
.B2(n_307),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2819),
.A2(n_307),
.B(n_308),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2815),
.B(n_308),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2811),
.B(n_309),
.Y(n_2826)
);

AO21x2_ASAP7_75t_L g2827 ( 
.A1(n_2809),
.A2(n_311),
.B(n_312),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_SL g2828 ( 
.A1(n_2813),
.A2(n_313),
.B1(n_314),
.B2(n_316),
.Y(n_2828)
);

OAI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2817),
.A2(n_314),
.B(n_316),
.Y(n_2829)
);

OAI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2810),
.A2(n_318),
.B(n_321),
.Y(n_2830)
);

AOI21xp5_ASAP7_75t_L g2831 ( 
.A1(n_2808),
.A2(n_322),
.B(n_324),
.Y(n_2831)
);

OA21x2_ASAP7_75t_L g2832 ( 
.A1(n_2818),
.A2(n_325),
.B(n_326),
.Y(n_2832)
);

AO21x2_ASAP7_75t_L g2833 ( 
.A1(n_2812),
.A2(n_325),
.B(n_327),
.Y(n_2833)
);

AOI22xp33_ASAP7_75t_L g2834 ( 
.A1(n_2823),
.A2(n_2822),
.B1(n_2816),
.B2(n_2814),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_R g2835 ( 
.A(n_2820),
.B(n_328),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2834),
.B(n_2821),
.Y(n_2836)
);

OAI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2824),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_2837)
);

OAI322xp33_ASAP7_75t_L g2838 ( 
.A1(n_2825),
.A2(n_331),
.A3(n_332),
.B1(n_334),
.B2(n_335),
.C1(n_336),
.C2(n_337),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2826),
.A2(n_2830),
.B1(n_2831),
.B2(n_2829),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2832),
.Y(n_2840)
);

INVx3_ASAP7_75t_L g2841 ( 
.A(n_2827),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2833),
.B(n_334),
.Y(n_2842)
);

XNOR2xp5_ASAP7_75t_L g2843 ( 
.A(n_2828),
.B(n_338),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2835),
.Y(n_2844)
);

AOI22xp33_ASAP7_75t_L g2845 ( 
.A1(n_2833),
.A2(n_1037),
.B1(n_1052),
.B2(n_340),
.Y(n_2845)
);

INVx1_ASAP7_75t_SL g2846 ( 
.A(n_2835),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2846),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_2847)
);

NOR2x1p5_ASAP7_75t_L g2848 ( 
.A(n_2840),
.B(n_339),
.Y(n_2848)
);

AOI221xp5_ASAP7_75t_L g2849 ( 
.A1(n_2841),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.C(n_344),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2844),
.A2(n_2842),
.B1(n_2843),
.B2(n_2836),
.Y(n_2850)
);

OAI222xp33_ASAP7_75t_L g2851 ( 
.A1(n_2845),
.A2(n_341),
.B1(n_343),
.B2(n_345),
.C1(n_346),
.C2(n_347),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2839),
.A2(n_345),
.B(n_346),
.Y(n_2852)
);

OA21x2_ASAP7_75t_L g2853 ( 
.A1(n_2837),
.A2(n_347),
.B(n_348),
.Y(n_2853)
);

OAI33xp33_ASAP7_75t_R g2854 ( 
.A1(n_2838),
.A2(n_351),
.A3(n_352),
.B1(n_354),
.B2(n_355),
.B3(n_356),
.Y(n_2854)
);

INVxp67_ASAP7_75t_SL g2855 ( 
.A(n_2840),
.Y(n_2855)
);

OAI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2840),
.A2(n_354),
.B(n_357),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2855),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2848),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_2858)
);

OAI31xp33_ASAP7_75t_L g2859 ( 
.A1(n_2851),
.A2(n_2850),
.A3(n_2852),
.B(n_2854),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2853),
.A2(n_1037),
.B1(n_1052),
.B2(n_364),
.Y(n_2860)
);

A2O1A1Ixp33_ASAP7_75t_SL g2861 ( 
.A1(n_2859),
.A2(n_2856),
.B(n_2847),
.C(n_2849),
.Y(n_2861)
);

OAI21xp5_ASAP7_75t_L g2862 ( 
.A1(n_2860),
.A2(n_362),
.B(n_363),
.Y(n_2862)
);

AO221x2_ASAP7_75t_L g2863 ( 
.A1(n_2858),
.A2(n_362),
.B1(n_363),
.B2(n_365),
.C(n_366),
.Y(n_2863)
);

AOI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2863),
.A2(n_2857),
.B1(n_2862),
.B2(n_2861),
.Y(n_2864)
);

AOI211xp5_ASAP7_75t_L g2865 ( 
.A1(n_2864),
.A2(n_367),
.B(n_368),
.C(n_369),
.Y(n_2865)
);


endmodule