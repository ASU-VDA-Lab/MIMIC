module fake_jpeg_19374_n_260 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_8),
.B(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx2_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_59),
.A2(n_70),
.B1(n_77),
.B2(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_62),
.B(n_67),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_19),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_26),
.B1(n_36),
.B2(n_18),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_68),
.B1(n_81),
.B2(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_26),
.B1(n_18),
.B2(n_37),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_80),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_30),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_45),
.B1(n_53),
.B2(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

HAxp5_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_19),
.CON(n_87),
.SN(n_87)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_35),
.B1(n_21),
.B2(n_27),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_21),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_34),
.B1(n_27),
.B2(n_24),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_97),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_54),
.B1(n_49),
.B2(n_47),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_113),
.B1(n_121),
.B2(n_78),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_24),
.B1(n_27),
.B2(n_35),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_47),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_68),
.C(n_58),
.Y(n_124)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_15),
.Y(n_114)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_24),
.B1(n_3),
.B2(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_146),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_79),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_104),
.B(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_R g131 ( 
.A(n_117),
.B(n_82),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_141),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_82),
.CI(n_84),
.CON(n_135),
.SN(n_135)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_137),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_63),
.B1(n_58),
.B2(n_72),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_142),
.B1(n_150),
.B2(n_111),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_11),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_63),
.B1(n_72),
.B2(n_78),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_84),
.C(n_85),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_147),
.C(n_101),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_60),
.B(n_4),
.C(n_5),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_14),
.C(n_13),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_173),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_120),
.B(n_115),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_94),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_116),
.B1(n_108),
.B2(n_93),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_134),
.B1(n_105),
.B2(n_125),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_148),
.B1(n_123),
.B2(n_134),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_94),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_172),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_99),
.B(n_102),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_131),
.B1(n_135),
.B2(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_153),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_189),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_195),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_196),
.B1(n_176),
.B2(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_146),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_151),
.C(n_163),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_201),
.C(n_204),
.Y(n_216)
);

XNOR2x2_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_168),
.C(n_161),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_206),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_209),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_166),
.C(n_154),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_147),
.C(n_10),
.Y(n_205)
);

NAND4xp25_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_10),
.C(n_184),
.D(n_7),
.Y(n_220)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_160),
.C(n_156),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_173),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_181),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_158),
.B(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_212),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_180),
.B1(n_194),
.B2(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_172),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

OAI22x1_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_193),
.B1(n_179),
.B2(n_177),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_218),
.B1(n_226),
.B2(n_213),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_5),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_186),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_191),
.C(n_195),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_197),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_202),
.B1(n_192),
.B2(n_194),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_198),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_229),
.C(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_201),
.C(n_207),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_223),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_234),
.B1(n_236),
.B2(n_215),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_208),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_180),
.B1(n_210),
.B2(n_179),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_215),
.B1(n_196),
.B2(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_188),
.B(n_222),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_6),
.B(n_7),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_227),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_245),
.B1(n_227),
.B2(n_239),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_233),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_119),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_143),
.C(n_8),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_143),
.C(n_105),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_8),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_255),
.C(n_257),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_9),
.Y(n_260)
);


endmodule