module real_jpeg_15106_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_311, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_311;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_68),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_68),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_3),
.A2(n_48),
.B1(n_53),
.B2(n_68),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_4),
.A2(n_35),
.B1(n_37),
.B2(n_167),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_4),
.A2(n_48),
.B1(n_53),
.B2(n_167),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_6),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_142),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_142),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_6),
.A2(n_48),
.B1(n_53),
.B2(n_142),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_7),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_188),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_7),
.A2(n_48),
.B1(n_53),
.B2(n_188),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_37),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_29),
.B1(n_64),
.B2(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_10),
.A2(n_29),
.B1(n_48),
.B2(n_53),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_11),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_43),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_11),
.A2(n_43),
.B1(n_48),
.B2(n_53),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_13),
.A2(n_61),
.B(n_64),
.C(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_13),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_13),
.B(n_103),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_181),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_13),
.A2(n_86),
.B1(n_89),
.B2(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_13),
.B(n_83),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_48),
.B1(n_53),
.B2(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_58),
.B1(n_64),
.B2(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_58),
.Y(n_114)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_104),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_84),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_21),
.B(n_74),
.CI(n_84),
.CON(n_306),
.SN(n_306)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_73),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_24),
.B(n_45),
.C(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_40),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_27),
.A2(n_32),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_28),
.A2(n_30),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g230 ( 
.A(n_28),
.B(n_181),
.CON(n_230),
.SN(n_230)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_30),
.A2(n_62),
.B(n_181),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_30),
.B(n_35),
.C(n_38),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_31),
.A2(n_113),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_31),
.A2(n_33),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_32),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_32),
.A2(n_41),
.B(n_114),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_32),
.A2(n_83),
.B1(n_184),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_32),
.A2(n_83),
.B1(n_217),
.B2(n_230),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_33),
.A2(n_82),
.B(n_115),
.Y(n_138)
);

OA22x2_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_34),
.A2(n_37),
.B(n_229),
.C(n_231),
.Y(n_228)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_37),
.B1(n_51),
.B2(n_54),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_37),
.B(n_251),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_44),
.A2(n_45),
.B1(n_112),
.B2(n_117),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_55),
.B(n_57),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_46),
.A2(n_55),
.B1(n_95),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_46),
.A2(n_55),
.B1(n_236),
.B2(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_46),
.A2(n_55),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_46),
.A2(n_55),
.B1(n_244),
.B2(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_79),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_47),
.A2(n_77),
.B(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_47),
.B(n_181),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g54 ( 
.A(n_51),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_51),
.B(n_53),
.C(n_181),
.Y(n_251)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_53),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_55),
.A2(n_57),
.B(n_96),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_55),
.Y(n_234)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_73),
.B1(n_107),
.B2(n_118),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_69),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_60),
.A2(n_99),
.B1(n_186),
.B2(n_189),
.Y(n_185)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_103),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_70),
.A2(n_103),
.B1(n_141),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_70),
.A2(n_103),
.B1(n_187),
.B2(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_75),
.B(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_76),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_114),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_92),
.B(n_97),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_97),
.B1(n_98),
.B2(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_85),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_85),
.A2(n_93),
.B1(n_94),
.B2(n_148),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B(n_90),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_86),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_86),
.A2(n_89),
.B1(n_259),
.B2(n_267),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_86),
.A2(n_130),
.B(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_87),
.A2(n_88),
.B1(n_160),
.B2(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_87),
.A2(n_91),
.B(n_162),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_87),
.A2(n_88),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_89),
.B(n_133),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_89),
.A2(n_131),
.B(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_89),
.B(n_181),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_102),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_99),
.A2(n_140),
.B(n_143),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_103),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_303),
.B(n_307),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_168),
.B(n_302),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_150),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_123),
.B(n_150),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_144),
.B2(n_149),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_124),
.B(n_145),
.C(n_146),
.Y(n_305)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_138),
.C(n_139),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_127),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_128),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_156),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_155),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_156),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.C(n_165),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_163),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_163),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_296),
.B(n_301),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_205),
.B1(n_221),
.B2(n_295),
.C(n_311),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_194),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_171),
.B(n_194),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_190),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_172),
.B(n_191),
.C(n_192),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.C(n_185),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_174),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_182),
.B(n_185),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_204),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_204),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_206),
.B(n_219),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_207),
.B(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_209),
.B(n_211),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_294),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_289),
.B(n_293),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_245),
.B(n_288),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_240),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_240),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_237),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_227),
.B(n_233),
.C(n_237),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_232),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_243),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_283),
.B(n_287),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_273),
.B(n_282),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_262),
.B(n_272),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_257),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_257),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_255),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_268),
.B(n_271),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_278),
.C(n_281),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_306),
.Y(n_310)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);


endmodule