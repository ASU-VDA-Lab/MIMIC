module fake_jpeg_801_n_99 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_14),
.C(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_36),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_0),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_32),
.B1(n_28),
.B2(n_33),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_39),
.B(n_38),
.C(n_30),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_32),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_54),
.B1(n_43),
.B2(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_58),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_39),
.B1(n_27),
.B2(n_29),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_29),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_43),
.C(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_64),
.Y(n_74)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_30),
.B1(n_28),
.B2(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_R g70 ( 
.A(n_69),
.B(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_78),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_35),
.B1(n_3),
.B2(n_5),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_79),
.B1(n_13),
.B2(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_63),
.C(n_10),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_85),
.B(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_18),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_91),
.B1(n_86),
.B2(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_90),
.B1(n_83),
.B2(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_88),
.B1(n_70),
.B2(n_21),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_19),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_20),
.B(n_22),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_26),
.C(n_23),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_24),
.Y(n_99)
);


endmodule