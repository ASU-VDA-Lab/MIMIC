module real_jpeg_9864_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_328, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_328;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_1),
.A2(n_20),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_1),
.B(n_33),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_45),
.B1(n_48),
.B2(n_53),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_1),
.A2(n_7),
.B(n_45),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_1),
.B(n_61),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_8),
.B(n_26),
.C(n_200),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_10),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_21),
.B1(n_45),
.B2(n_48),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_3),
.A2(n_21),
.B1(n_41),
.B2(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_10),
.B1(n_20),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_45),
.B1(n_48),
.B2(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_4),
.A2(n_41),
.B1(n_52),
.B2(n_57),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_57),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_7),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_7),
.B(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_8),
.A2(n_41),
.B1(n_52),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_26),
.B(n_62),
.C(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_8),
.B(n_26),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_10),
.A2(n_11),
.B1(n_20),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_11),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_11),
.A2(n_45),
.B1(n_48),
.B2(n_103),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_41),
.B1(n_52),
.B2(n_103),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_16),
.C(n_284),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_79),
.B(n_324),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_34),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_16),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_29),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_17),
.A2(n_25),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_18),
.B(n_101),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_22),
.B(n_31),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_22),
.A2(n_25),
.B(n_31),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_24),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_26),
.B(n_28),
.Y(n_130)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_27),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_29),
.B(n_114),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_32),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_33),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_35),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_71),
.C(n_73),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_36),
.A2(n_37),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_54),
.C(n_58),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_38),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_38),
.A2(n_105),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_38),
.A2(n_58),
.B1(n_59),
.B2(n_105),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_49),
.B(n_50),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_39),
.A2(n_96),
.B(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_40),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_40),
.B(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_40),
.B(n_97),
.Y(n_205)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_41),
.A2(n_53),
.B(n_63),
.Y(n_200)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_44),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_44),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_44),
.B(n_51),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_90),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_47),
.A2(n_52),
.B(n_53),
.C(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_48),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_49),
.B(n_53),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_49),
.A2(n_205),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_53),
.B(n_90),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_54),
.A2(n_55),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_67),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_62),
.B(n_70),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_62),
.A2(n_65),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_64),
.B(n_66),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_66),
.A2(n_143),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_71),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_71),
.A2(n_73),
.B1(n_248),
.B2(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_73),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_74),
.B(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_77),
.B(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_317),
.B(n_323),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_293),
.A3(n_312),
.B1(n_315),
.B2(n_316),
.C(n_328),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_271),
.B(n_292),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_252),
.B(n_270),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_151),
.B(n_234),
.C(n_251),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_134),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_85),
.B(n_134),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_110),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_99),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_87),
.B(n_99),
.C(n_110),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_88),
.B(n_95),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_93),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_89),
.A2(n_90),
.B(n_149),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_92),
.B(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_91),
.B(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_93),
.B(n_174),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_96),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_98),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_106),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_105),
.B(n_297),
.C(n_302),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_121),
.B1(n_122),
.B2(n_133),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_120),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_112),
.B(n_120),
.C(n_121),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_125),
.B(n_191),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_135),
.A2(n_136),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_142),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_143),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_233),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_227),
.B(n_232),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_212),
.B(n_226),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_193),
.B(n_211),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_181),
.B(n_192),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_170),
.B(n_180),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_162),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_166),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_175),
.B(n_179),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_183),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_202),
.B1(n_203),
.B2(n_210),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_197),
.A2(n_198),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_197),
.A2(n_198),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_197),
.A2(n_285),
.B(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_198),
.B(n_267),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_205),
.B(n_222),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_208),
.B(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_221),
.C(n_225),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_236),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_249),
.B2(n_250),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_243),
.C(n_250),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_241),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_254),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_269),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_265),
.B2(n_266),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_266),
.C(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_260),
.C(n_264),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_262),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_273),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_290),
.B2(n_291),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_281),
.B1(n_288),
.B2(n_289),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_289),
.C(n_291),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B(n_280),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_295),
.C(n_304),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_280),
.B(n_295),
.CI(n_304),
.CON(n_314),
.SN(n_314)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_282),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_283),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_305),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_297),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_307),
.C(n_311),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_320),
.Y(n_322)
);


endmodule