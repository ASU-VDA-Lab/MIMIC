module fake_netlist_6_3317_n_2778 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2778);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2778;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_873;
wire n_461;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_1550;
wire n_2703;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_405;
wire n_2660;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_2674;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_2733;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_411;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_420;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_2265;
wire n_2615;
wire n_414;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_924;
wire n_475;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_629;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g404 ( 
.A(n_237),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_258),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_281),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_341),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_358),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_128),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_176),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_236),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_41),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_311),
.Y(n_414)
);

BUFx10_ASAP7_75t_L g415 ( 
.A(n_275),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_88),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_7),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_174),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_200),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_63),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_296),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_151),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_44),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_19),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_2),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_95),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_183),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_321),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_270),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_371),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_266),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_110),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_356),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_18),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_20),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_114),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_151),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_328),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_228),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_324),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_110),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_231),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_75),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_345),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_53),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_132),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_116),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_317),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_242),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_129),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_306),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_158),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_251),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_129),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_347),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_9),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_19),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_87),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_139),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_111),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_294),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_155),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_262),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_40),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_111),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_237),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_130),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_283),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_11),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_336),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_109),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_160),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_261),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_359),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_8),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_292),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_287),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_125),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_72),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_163),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_145),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_142),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_102),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_210),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_332),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_337),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_171),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_59),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_379),
.Y(n_492)
);

BUFx5_ASAP7_75t_L g493 ( 
.A(n_62),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_119),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_51),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_210),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_382),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_41),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_257),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_58),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_236),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_159),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_307),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_37),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_94),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_227),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_183),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_355),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_94),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_393),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_331),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_263),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_254),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_327),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_58),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_167),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_35),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_301),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_167),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_351),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_277),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_184),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_232),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_230),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_20),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_357),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_165),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_4),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_113),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_189),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_118),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_135),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_124),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_66),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_349),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_244),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_365),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_172),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_64),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_383),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_310),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_313),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_218),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_187),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_398),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_217),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_165),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_208),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_288),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_56),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_22),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_149),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_23),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_93),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_304),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_109),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_113),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_255),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_2),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_136),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_259),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_377),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_297),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_85),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_103),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_85),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_250),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_253),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_369),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_228),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_222),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_293),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_84),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_243),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_264),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_83),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_335),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_390),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_244),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_93),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_123),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_380),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_140),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_308),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_3),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_81),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_83),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_107),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_114),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_289),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_133),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_350),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_240),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_170),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_238),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_249),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_13),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_51),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_342),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_224),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_102),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_177),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_75),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_21),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_216),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_400),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_239),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_333),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_239),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_63),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_256),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_79),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_403),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_158),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_173),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_13),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_376),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_62),
.Y(n_619)
);

CKINVDCx11_ASAP7_75t_R g620 ( 
.A(n_375),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_184),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_92),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_56),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_218),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_299),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_330),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_71),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_278),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_156),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_6),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_385),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_230),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_322),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_127),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_214),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_117),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_234),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_89),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_97),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_162),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_11),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_73),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_295),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_108),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_15),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_284),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_367),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_26),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_59),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_267),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_42),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_260),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_280),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_163),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_34),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_78),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_344),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_305),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_126),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_30),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_314),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_176),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_189),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_30),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_226),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_84),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_10),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_124),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_132),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_144),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_205),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_200),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_136),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_65),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_149),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_186),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_73),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_245),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_170),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_39),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_340),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_315),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_4),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_374),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_133),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_95),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_353),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_33),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_140),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_334),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_248),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_268),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_166),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_162),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_199),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_134),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_384),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_362),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_394),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_8),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_179),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_97),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_401),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_178),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_372),
.Y(n_705)
);

CKINVDCx16_ASAP7_75t_R g706 ( 
.A(n_173),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_213),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_190),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_107),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_192),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_42),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_493),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_R g713 ( 
.A(n_412),
.B(n_0),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_474),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_412),
.B(n_0),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_474),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_600),
.B(n_1),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_493),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_493),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_620),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_432),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_407),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_493),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_493),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_493),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_589),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_488),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_600),
.B(n_1),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_492),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_605),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_455),
.Y(n_731)
);

INVxp33_ASAP7_75t_SL g732 ( 
.A(n_605),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_546),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_493),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_493),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_493),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_408),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_414),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_617),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_455),
.B(n_3),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_497),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_617),
.B(n_5),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_497),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_421),
.Y(n_744)
);

CKINVDCx16_ASAP7_75t_R g745 ( 
.A(n_589),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_649),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_430),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_431),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_497),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_682),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_423),
.B(n_5),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_434),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_497),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_497),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_497),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_439),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_649),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_441),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_404),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_450),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_523),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_632),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_516),
.B(n_6),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_404),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_457),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_465),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_523),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_523),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_523),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_471),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_632),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_523),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_423),
.B(n_445),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_473),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_477),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_523),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_577),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_577),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_577),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_577),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_577),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_692),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_479),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_577),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_480),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_406),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_672),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_455),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_498),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_504),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_516),
.B(n_7),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_672),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_706),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_445),
.B(n_9),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_672),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_672),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_672),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_509),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_446),
.B(n_10),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_406),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_672),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_511),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_512),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_446),
.B(n_12),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_683),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_495),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_683),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_683),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_683),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_683),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_683),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_453),
.B(n_12),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_451),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_453),
.B(n_14),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_618),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_514),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_451),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_451),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_427),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_706),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_515),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_427),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_409),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_618),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_489),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_519),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_462),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_448),
.B(n_14),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_572),
.B(n_15),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_495),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_521),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_462),
.Y(n_832)
);

CKINVDCx16_ASAP7_75t_R g833 ( 
.A(n_486),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_582),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_582),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_586),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_527),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_586),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_536),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_665),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_538),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_541),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_542),
.Y(n_843)
);

CKINVDCx16_ASAP7_75t_R g844 ( 
.A(n_486),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_550),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_665),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_409),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_556),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_696),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_559),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_563),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_696),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_743),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_722),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_743),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_731),
.B(n_448),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_788),
.B(n_448),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_806),
.B(n_456),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_749),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_741),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_741),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_749),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_753),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_721),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_737),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_738),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_744),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_747),
.B(n_495),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_753),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_761),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_844),
.B(n_415),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_754),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_748),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_754),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_755),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_830),
.B(n_456),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_761),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_727),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_712),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_755),
.A2(n_476),
.B(n_467),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_712),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_752),
.B(n_687),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_756),
.B(n_576),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_736),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_767),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_784),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_828),
.B(n_456),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_729),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_828),
.B(n_687),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_784),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_767),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_768),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_768),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_733),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_742),
.B(n_678),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_769),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_758),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_769),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_772),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_795),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_SL g901 ( 
.A(n_825),
.B(n_415),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_736),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_795),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_760),
.B(n_687),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_765),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_797),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_772),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_797),
.B(n_690),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_750),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_776),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_776),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_766),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_732),
.A2(n_713),
.B1(n_715),
.B2(n_786),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_770),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_774),
.B(n_690),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_777),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_777),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_778),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_778),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_779),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_775),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_779),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_780),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_780),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_800),
.Y(n_925)
);

OA21x2_ASAP7_75t_L g926 ( 
.A1(n_781),
.A2(n_476),
.B(n_467),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_781),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_787),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_787),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_792),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_783),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_792),
.Y(n_932)
);

OA21x2_ASAP7_75t_L g933 ( 
.A1(n_796),
.A2(n_522),
.B(n_513),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_796),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_785),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_801),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_742),
.B(n_464),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_801),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_805),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_805),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_807),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_807),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_808),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_808),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_809),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_809),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_789),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_810),
.B(n_690),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_790),
.B(n_705),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_798),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_802),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_R g954 ( 
.A(n_720),
.B(n_564),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_726),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_803),
.B(n_705),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_811),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_811),
.B(n_705),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_819),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_819),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_782),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_718),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_815),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_835),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_816),
.B(n_463),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_771),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_821),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_718),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_719),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_835),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_826),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_719),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_837),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_740),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_723),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_723),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_844),
.B(n_415),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_975),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_965),
.B(n_463),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_968),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_856),
.B(n_745),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_906),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_870),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_955),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_975),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_976),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_974),
.B(n_839),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_870),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_883),
.A2(n_831),
.B1(n_843),
.B2(n_842),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_889),
.B(n_841),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_968),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_877),
.Y(n_992)
);

AND2x6_ASAP7_75t_L g993 ( 
.A(n_889),
.B(n_405),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_906),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_854),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_976),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_954),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_887),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_865),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_868),
.B(n_848),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_889),
.B(n_500),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_864),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_889),
.B(n_887),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_969),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_877),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_882),
.B(n_850),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_904),
.B(n_851),
.Y(n_1007)
);

INVx5_ASAP7_75t_L g1008 ( 
.A(n_895),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_969),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_962),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_908),
.B(n_813),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_937),
.B(n_745),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_906),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_856),
.B(n_793),
.Y(n_1014)
);

NOR2x1p5_ASAP7_75t_L g1015 ( 
.A(n_866),
.B(n_464),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_915),
.B(n_500),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_871),
.B(n_728),
.C(n_717),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_879),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_962),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_962),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_938),
.B(n_464),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_857),
.B(n_793),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_968),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_951),
.B(n_730),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_895),
.A2(n_773),
.B1(n_794),
.B2(n_751),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_879),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_968),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_968),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_968),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_972),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_972),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_956),
.B(n_724),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_857),
.B(n_820),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_858),
.B(n_876),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_972),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_913),
.A2(n_845),
.B1(n_746),
.B2(n_820),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_895),
.A2(n_804),
.B1(n_812),
.B2(n_799),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_895),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_R g1040 ( 
.A(n_963),
.B(n_714),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_972),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_972),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_972),
.Y(n_1043)
);

INVx3_ASAP7_75t_R g1044 ( 
.A(n_963),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_858),
.B(n_876),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_879),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_879),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_908),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_908),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_908),
.B(n_813),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_853),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_938),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_860),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_966),
.B(n_714),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_950),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_895),
.Y(n_1056)
);

INVx5_ASAP7_75t_L g1057 ( 
.A(n_895),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_895),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_925),
.Y(n_1059)
);

CKINVDCx8_ASAP7_75t_R g1060 ( 
.A(n_867),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_873),
.Y(n_1061)
);

AND2x6_ASAP7_75t_L g1062 ( 
.A(n_950),
.B(n_405),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_853),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_860),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_895),
.B(n_724),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_950),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_977),
.A2(n_824),
.B1(n_833),
.B2(n_716),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_886),
.B(n_678),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_855),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_924),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_855),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_859),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_878),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_913),
.A2(n_814),
.B1(n_763),
.B2(n_791),
.Y(n_1074)
);

AND2x6_ASAP7_75t_L g1075 ( 
.A(n_950),
.B(n_405),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_859),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_958),
.B(n_725),
.Y(n_1077)
);

NOR2x1p5_ASAP7_75t_L g1078 ( 
.A(n_897),
.B(n_553),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_958),
.B(n_633),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_888),
.Y(n_1080)
);

INVx8_ASAP7_75t_L g1081 ( 
.A(n_905),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_958),
.B(n_633),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_958),
.B(n_678),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_862),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_959),
.A2(n_823),
.B1(n_847),
.B2(n_764),
.C(n_759),
.Y(n_1085)
);

BUFx10_ASAP7_75t_L g1086 ( 
.A(n_912),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_894),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_959),
.B(n_553),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_862),
.B(n_725),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_863),
.B(n_734),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_914),
.B(n_678),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_924),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_863),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_921),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_931),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_869),
.B(n_734),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_960),
.B(n_553),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_861),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_861),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_935),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_869),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_861),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_872),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_948),
.B(n_716),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_952),
.B(n_678),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_909),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_890),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_880),
.B(n_643),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_880),
.A2(n_598),
.B1(n_666),
.B2(n_572),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_872),
.Y(n_1110)
);

AND2x6_ASAP7_75t_L g1111 ( 
.A(n_874),
.B(n_513),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_880),
.B(n_652),
.Y(n_1112)
);

CKINVDCx16_ASAP7_75t_R g1113 ( 
.A(n_901),
.Y(n_1113)
);

NAND3x1_ASAP7_75t_L g1114 ( 
.A(n_960),
.B(n_413),
.C(n_410),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_874),
.Y(n_1115)
);

AND2x6_ASAP7_75t_L g1116 ( 
.A(n_875),
.B(n_522),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_964),
.B(n_817),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_875),
.B(n_735),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_953),
.B(n_739),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_885),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_885),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_891),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_961),
.B(n_757),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_967),
.B(n_735),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_891),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_971),
.B(n_822),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_892),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_892),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_893),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_973),
.B(n_822),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_964),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_886),
.B(n_678),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_880),
.A2(n_658),
.B1(n_661),
.B2(n_653),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_893),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_932),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_926),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_896),
.B(n_598),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_970),
.B(n_817),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1032),
.B(n_881),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1024),
.B(n_483),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1048),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_997),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1024),
.B(n_487),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1049),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1000),
.B(n_881),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1035),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1000),
.B(n_881),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_997),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1035),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1006),
.B(n_881),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1034),
.A2(n_666),
.B(n_575),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1060),
.Y(n_1152)
);

AO22x1_ASAP7_75t_L g1153 ( 
.A1(n_1017),
.A2(n_413),
.B1(n_424),
.B2(n_410),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1017),
.B(n_829),
.C(n_417),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1055),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_1081),
.B(n_560),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1059),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1006),
.B(n_902),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1007),
.B(n_902),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1052),
.A2(n_440),
.B(n_447),
.C(n_424),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1053),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1055),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1066),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1007),
.B(n_902),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1018),
.B(n_902),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_995),
.B(n_999),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1081),
.B(n_560),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1053),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1018),
.B(n_896),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1126),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1073),
.Y(n_1171)
);

OAI221xp5_ASAP7_75t_L g1172 ( 
.A1(n_1038),
.A2(n_458),
.B1(n_459),
.B2(n_447),
.C(n_440),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1045),
.B(n_491),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1026),
.B(n_898),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1066),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1008),
.B(n_697),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1008),
.B(n_568),
.Y(n_1177)
);

INVxp67_ASAP7_75t_SL g1178 ( 
.A(n_1026),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1012),
.B(n_502),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1008),
.B(n_569),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1008),
.B(n_570),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_981),
.B(n_486),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1045),
.B(n_594),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1047),
.B(n_898),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1002),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1003),
.A2(n_884),
.B(n_899),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1011),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1039),
.B(n_573),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1052),
.B(n_987),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1047),
.B(n_899),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1011),
.Y(n_1191)
);

AND2x6_ASAP7_75t_SL g1192 ( 
.A(n_1123),
.B(n_458),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1124),
.B(n_907),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_989),
.B(n_970),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_L g1195 ( 
.A(n_1038),
.B(n_419),
.C(n_416),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1124),
.B(n_907),
.Y(n_1196)
);

AND2x6_ASAP7_75t_L g1197 ( 
.A(n_1133),
.B(n_543),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1011),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1039),
.B(n_578),
.Y(n_1199)
);

OR2x6_ASAP7_75t_L g1200 ( 
.A(n_1081),
.B(n_560),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_978),
.B(n_910),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_985),
.B(n_910),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1039),
.B(n_579),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1021),
.B(n_575),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1050),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1119),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1087),
.B(n_575),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1050),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1039),
.B(n_583),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1064),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1021),
.B(n_655),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_986),
.B(n_911),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1014),
.B(n_641),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1050),
.Y(n_1214)
);

INVx8_ASAP7_75t_L g1215 ( 
.A(n_1054),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1056),
.B(n_585),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1136),
.A2(n_933),
.B1(n_926),
.B2(n_460),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1056),
.B(n_593),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1022),
.B(n_486),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1130),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1056),
.B(n_607),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_998),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1046),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_996),
.B(n_911),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1122),
.B(n_916),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1033),
.B(n_677),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_998),
.B(n_420),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_990),
.B(n_425),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1056),
.B(n_609),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1104),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1101),
.B(n_1074),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1015),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1136),
.A2(n_933),
.B1(n_926),
.B2(n_460),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1025),
.A2(n_470),
.B(n_472),
.C(n_459),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1101),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1057),
.B(n_612),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1122),
.B(n_916),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1064),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1119),
.B(n_496),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1057),
.B(n_614),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1025),
.A2(n_562),
.B1(n_591),
.B2(n_543),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1128),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1128),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_933),
.B1(n_926),
.B2(n_472),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1129),
.B(n_918),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1129),
.B(n_918),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1046),
.B(n_982),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_982),
.B(n_928),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_994),
.B(n_928),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1054),
.B(n_655),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1098),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_994),
.B(n_929),
.Y(n_1252)
);

NAND2x1_ASAP7_75t_L g1253 ( 
.A(n_1058),
.B(n_890),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1117),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1098),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1013),
.B(n_929),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1013),
.B(n_930),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1078),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1131),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1099),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1099),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1040),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1051),
.B(n_930),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1095),
.B(n_655),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_980),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_L g1266 ( 
.A(n_993),
.B(n_631),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1109),
.A2(n_485),
.B(n_490),
.C(n_470),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1117),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_993),
.A2(n_684),
.B1(n_698),
.B2(n_650),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1102),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_993),
.A2(n_933),
.B1(n_490),
.B2(n_494),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1117),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1063),
.B(n_936),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1069),
.B(n_936),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1102),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1057),
.B(n_699),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1040),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1071),
.B(n_939),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1091),
.B(n_426),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1057),
.B(n_562),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1072),
.B(n_939),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1076),
.B(n_944),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1084),
.B(n_944),
.Y(n_1283)
);

INVx8_ASAP7_75t_L g1284 ( 
.A(n_1054),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1093),
.B(n_945),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1103),
.B(n_945),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1131),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1138),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1110),
.B(n_949),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1107),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_993),
.A2(n_597),
.B1(n_625),
.B2(n_591),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1058),
.B(n_597),
.Y(n_1292)
);

AO22x1_ASAP7_75t_L g1293 ( 
.A1(n_1037),
.A2(n_993),
.B1(n_1116),
.B2(n_1111),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1077),
.B(n_625),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1115),
.B(n_949),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1120),
.B(n_957),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1123),
.B(n_428),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_995),
.B(n_411),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1088),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1121),
.B(n_957),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1138),
.Y(n_1301)
);

NOR2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1002),
.B(n_433),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1108),
.A2(n_628),
.B1(n_646),
.B2(n_626),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1091),
.B(n_435),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1134),
.B(n_932),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1138),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1016),
.B(n_932),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_999),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1016),
.B(n_932),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1001),
.A2(n_884),
.B(n_919),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1065),
.B(n_626),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1108),
.B(n_628),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1088),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_983),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1107),
.Y(n_1316)
);

NAND2xp33_ASAP7_75t_L g1317 ( 
.A(n_1062),
.B(n_646),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1085),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1097),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_979),
.B(n_934),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1112),
.B(n_647),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1097),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1100),
.B(n_246),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_983),
.Y(n_1324)
);

NOR2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1080),
.B(n_436),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1004),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_988),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_979),
.B(n_934),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_984),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1137),
.A2(n_494),
.B(n_501),
.C(n_485),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1009),
.B(n_934),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1001),
.A2(n_884),
.B(n_919),
.Y(n_1332)
);

NAND2x1_ASAP7_75t_L g1333 ( 
.A(n_1062),
.B(n_890),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1079),
.A2(n_884),
.B(n_920),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1254),
.B(n_1105),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1171),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1172),
.A2(n_1075),
.B1(n_1062),
.B2(n_1111),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1189),
.B(n_1113),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1189),
.B(n_1105),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1155),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1206),
.B(n_1067),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1140),
.B(n_1061),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1193),
.B(n_1112),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1152),
.B(n_1080),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1178),
.A2(n_1031),
.B(n_991),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1142),
.Y(n_1346)
);

BUFx4f_ASAP7_75t_L g1347 ( 
.A(n_1215),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1196),
.B(n_1062),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1141),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1268),
.B(n_1272),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1155),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1140),
.B(n_1062),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1215),
.B(n_1123),
.Y(n_1353)
);

BUFx8_ASAP7_75t_L g1354 ( 
.A(n_1259),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1157),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1144),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1288),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1301),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1143),
.B(n_1061),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1222),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1143),
.B(n_1075),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1145),
.B(n_1075),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1262),
.B(n_1086),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1315),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1277),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1307),
.Y(n_1366)
);

AND3x1_ASAP7_75t_SL g1367 ( 
.A(n_1302),
.B(n_518),
.C(n_501),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1147),
.B(n_1150),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1315),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1185),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1148),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1158),
.B(n_1075),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_L g1373 ( 
.A(n_1287),
.B(n_1083),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1324),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1231),
.A2(n_1082),
.B1(n_1079),
.B2(n_1083),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1230),
.A2(n_1044),
.B1(n_418),
.B2(n_438),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1313),
.A2(n_1028),
.B(n_1027),
.Y(n_1377)
);

AND2x6_ASAP7_75t_SL g1378 ( 
.A(n_1207),
.B(n_1156),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1231),
.B(n_1086),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1307),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1155),
.B(n_1094),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1213),
.B(n_1094),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1327),
.Y(n_1383)
);

CKINVDCx6p67_ASAP7_75t_R g1384 ( 
.A(n_1309),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1213),
.B(n_1106),
.Y(n_1385)
);

AO22x1_ASAP7_75t_L g1386 ( 
.A1(n_1197),
.A2(n_442),
.B1(n_443),
.B2(n_437),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1215),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1166),
.B(n_422),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1155),
.B(n_980),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1159),
.B(n_1075),
.Y(n_1390)
);

INVx3_ASAP7_75t_SL g1391 ( 
.A(n_1284),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1164),
.B(n_1010),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1162),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1234),
.A2(n_1082),
.B(n_1137),
.C(n_1090),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1207),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1204),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1187),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1329),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1146),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1173),
.B(n_1019),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_R g1401 ( 
.A(n_1298),
.B(n_526),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1162),
.B(n_980),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1271),
.B(n_980),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1173),
.B(n_1020),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1191),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1333),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1313),
.A2(n_1132),
.B(n_1030),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1198),
.B(n_647),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_R g1409 ( 
.A(n_1232),
.B(n_529),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1205),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1149),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1284),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1183),
.B(n_1029),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1208),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1214),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1228),
.A2(n_1116),
.B1(n_1111),
.B2(n_1041),
.Y(n_1416)
);

INVx5_ASAP7_75t_L g1417 ( 
.A(n_1265),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1223),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1161),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1284),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1163),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1175),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1170),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1183),
.B(n_1036),
.Y(n_1424)
);

NAND2xp33_ASAP7_75t_SL g1425 ( 
.A(n_1271),
.B(n_574),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1250),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1228),
.B(n_1043),
.Y(n_1427)
);

AND2x6_ASAP7_75t_SL g1428 ( 
.A(n_1207),
.B(n_518),
.Y(n_1428)
);

NOR3xp33_ASAP7_75t_SL g1429 ( 
.A(n_1226),
.B(n_449),
.C(n_444),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1223),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1303),
.B(n_1111),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1179),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1326),
.Y(n_1433)
);

AND3x2_ASAP7_75t_SL g1434 ( 
.A(n_1153),
.B(n_587),
.C(n_584),
.Y(n_1434)
);

AND2x6_ASAP7_75t_L g1435 ( 
.A(n_1182),
.B(n_657),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1242),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1168),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1226),
.B(n_496),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1220),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1265),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1210),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1243),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1279),
.B(n_1111),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1217),
.B(n_1023),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

NOR3xp33_ASAP7_75t_SL g1446 ( 
.A(n_1154),
.B(n_454),
.C(n_452),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1197),
.A2(n_1116),
.B1(n_1092),
.B2(n_1070),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_R g1448 ( 
.A(n_1258),
.B(n_601),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1235),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1279),
.B(n_1116),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1238),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_L g1452 ( 
.A(n_1156),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1299),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1197),
.A2(n_1116),
.B1(n_1092),
.B2(n_1070),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1239),
.A2(n_630),
.B1(n_676),
.B2(n_624),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1251),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1255),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1319),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1322),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1305),
.B(n_1089),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1305),
.B(n_1096),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1260),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1156),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1167),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1261),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1225),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_R g1467 ( 
.A(n_1317),
.B(n_710),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1270),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1318),
.B(n_1118),
.Y(n_1469)
);

OR2x2_ASAP7_75t_SL g1470 ( 
.A(n_1195),
.B(n_520),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_R g1471 ( 
.A(n_1297),
.B(n_461),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1237),
.B(n_1135),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1234),
.A2(n_524),
.B(n_530),
.C(n_520),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1204),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1245),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1219),
.B(n_496),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1246),
.Y(n_1477)
);

AND2x2_ASAP7_75t_SL g1478 ( 
.A(n_1217),
.B(n_657),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1201),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1227),
.B(n_466),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1275),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1211),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1233),
.B(n_1227),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1211),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1194),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1264),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1469),
.B(n_1479),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1377),
.A2(n_1306),
.B(n_1186),
.Y(n_1488)
);

AOI211x1_ASAP7_75t_L g1489 ( 
.A1(n_1483),
.A2(n_1241),
.B(n_1151),
.C(n_1293),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1417),
.A2(n_1403),
.B(n_1247),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1469),
.B(n_1233),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1417),
.A2(n_1321),
.B(n_1165),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1466),
.B(n_1197),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1375),
.A2(n_1304),
.A3(n_1160),
.B(n_1330),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1475),
.B(n_1197),
.Y(n_1495)
);

AOI21xp33_ASAP7_75t_L g1496 ( 
.A1(n_1339),
.A2(n_1321),
.B(n_1294),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1477),
.B(n_1139),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1349),
.Y(n_1498)
);

NOR2x1_ASAP7_75t_SL g1499 ( 
.A(n_1417),
.B(n_1292),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1368),
.A2(n_1394),
.B(n_1343),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1342),
.B(n_1264),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1478),
.A2(n_1244),
.B1(n_1267),
.B2(n_1160),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1399),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1440),
.B(n_1323),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1478),
.B(n_1202),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1432),
.B(n_1264),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1474),
.B(n_1325),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1417),
.A2(n_1174),
.B(n_1169),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1403),
.A2(n_1190),
.B(n_1184),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1342),
.B(n_1212),
.Y(n_1510)
);

AO22x2_ASAP7_75t_L g1511 ( 
.A1(n_1438),
.A2(n_1434),
.B1(n_1338),
.B2(n_1480),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1359),
.B(n_1167),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1356),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1362),
.A2(n_1266),
.B(n_1253),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1372),
.A2(n_1292),
.B(n_1031),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1359),
.B(n_1224),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1344),
.Y(n_1517)
);

BUFx5_ASAP7_75t_L g1518 ( 
.A(n_1366),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1473),
.A2(n_1330),
.A3(n_1267),
.B(n_1310),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1385),
.B(n_1167),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1337),
.A2(n_1244),
.B1(n_1291),
.B2(n_1273),
.Y(n_1521)
);

AOI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1413),
.A2(n_1180),
.B(n_1177),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1390),
.A2(n_1450),
.B(n_1443),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1370),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1460),
.B(n_1263),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1337),
.A2(n_1274),
.B1(n_1281),
.B2(n_1278),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1426),
.B(n_1200),
.Y(n_1527)
);

NAND2x1p5_ASAP7_75t_L g1528 ( 
.A(n_1440),
.B(n_1418),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1357),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1365),
.B(n_1200),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1461),
.B(n_1282),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1355),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1379),
.A2(n_1283),
.B1(n_1286),
.B2(n_1285),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1444),
.A2(n_1312),
.B(n_1294),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1444),
.A2(n_1312),
.B(n_1320),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1345),
.A2(n_1308),
.B(n_1328),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1382),
.B(n_1289),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1402),
.A2(n_1331),
.B(n_1249),
.Y(n_1538)
);

AOI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1424),
.A2(n_1389),
.B(n_1427),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1402),
.A2(n_1252),
.B(n_1248),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1420),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_SL g1542 ( 
.A(n_1401),
.B(n_469),
.C(n_468),
.Y(n_1542)
);

O2A1O1Ixp5_ASAP7_75t_L g1543 ( 
.A1(n_1352),
.A2(n_1180),
.B(n_1181),
.C(n_1177),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1336),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1400),
.B(n_1404),
.Y(n_1545)
);

AO31x2_ASAP7_75t_L g1546 ( 
.A1(n_1473),
.A2(n_1257),
.A3(n_1256),
.B(n_1295),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1449),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1348),
.A2(n_991),
.B(n_1176),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1340),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1341),
.A2(n_1425),
.B(n_1379),
.C(n_1335),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1425),
.B(n_1296),
.Y(n_1551)
);

AO31x2_ASAP7_75t_L g1552 ( 
.A1(n_1361),
.A2(n_1300),
.A3(n_1316),
.B(n_1290),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1389),
.A2(n_1332),
.B(n_1311),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1439),
.B(n_1363),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1431),
.A2(n_1176),
.B(n_1042),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1341),
.B(n_1200),
.C(n_1269),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1392),
.A2(n_1334),
.B(n_1188),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_1358),
.C(n_1397),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1472),
.A2(n_1188),
.B(n_1181),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1335),
.B(n_988),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1470),
.A2(n_530),
.B1(n_531),
.B2(n_524),
.Y(n_1561)
);

CKINVDCx6p67_ASAP7_75t_R g1562 ( 
.A(n_1391),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1336),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1364),
.A2(n_1203),
.B(n_1199),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1405),
.A2(n_532),
.B1(n_535),
.B2(n_531),
.Y(n_1565)
);

AO31x2_ASAP7_75t_L g1566 ( 
.A1(n_1364),
.A2(n_691),
.A3(n_703),
.B(n_681),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1369),
.A2(n_1203),
.B(n_1199),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1410),
.B(n_1209),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1370),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1369),
.A2(n_691),
.A3(n_703),
.B(n_681),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1414),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1340),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1415),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1560),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1500),
.A2(n_1416),
.B(n_1447),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1550),
.A2(n_1338),
.B(n_1476),
.Y(n_1576)
);

AO21x1_ASAP7_75t_L g1577 ( 
.A1(n_1500),
.A2(n_1408),
.B(n_1381),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1558),
.B(n_1350),
.Y(n_1578)
);

AO21x2_ASAP7_75t_L g1579 ( 
.A1(n_1523),
.A2(n_1454),
.B(n_1407),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1544),
.Y(n_1580)
);

BUFx4f_ASAP7_75t_L g1581 ( 
.A(n_1528),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1487),
.B(n_1393),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1491),
.A2(n_1487),
.B1(n_1531),
.B2(n_1525),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1496),
.A2(n_1534),
.B(n_1535),
.Y(n_1584)
);

BUFx10_ASAP7_75t_L g1585 ( 
.A(n_1517),
.Y(n_1585)
);

OAI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1510),
.A2(n_1452),
.B1(n_1433),
.B2(n_1360),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1488),
.A2(n_1536),
.B(n_1559),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1514),
.A2(n_1381),
.B(n_1399),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1496),
.A2(n_1419),
.B(n_1411),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1531),
.B(n_1393),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1534),
.A2(n_1407),
.B(n_1446),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1505),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1509),
.A2(n_1429),
.B(n_1435),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1516),
.B(n_1360),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1535),
.A2(n_1419),
.B(n_1411),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1501),
.B(n_1363),
.Y(n_1597)
);

AO31x2_ASAP7_75t_L g1598 ( 
.A1(n_1502),
.A2(n_1441),
.A3(n_1456),
.B(n_1437),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1502),
.A2(n_1455),
.B1(n_1452),
.B2(n_1422),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1543),
.A2(n_1435),
.B(n_1408),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1532),
.Y(n_1601)
);

BUFx12f_ASAP7_75t_L g1602 ( 
.A(n_1541),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1538),
.A2(n_1441),
.B(n_1437),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1551),
.A2(n_1557),
.B(n_1522),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1564),
.A2(n_1457),
.B(n_1456),
.Y(n_1605)
);

O2A1O1Ixp5_ASAP7_75t_L g1606 ( 
.A1(n_1539),
.A2(n_1209),
.B(n_1218),
.C(n_1216),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1567),
.A2(n_1462),
.B(n_1457),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1503),
.Y(n_1608)
);

OAI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1561),
.A2(n_1401),
.B(n_1388),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1537),
.B(n_1346),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1511),
.A2(n_1435),
.B1(n_1485),
.B2(n_1350),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1518),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1555),
.A2(n_1465),
.B(n_1462),
.Y(n_1613)
);

OAI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1561),
.A2(n_1497),
.B1(n_1521),
.B2(n_1513),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1547),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1563),
.Y(n_1616)
);

BUFx2_ASAP7_75t_SL g1617 ( 
.A(n_1572),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1518),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1515),
.A2(n_1430),
.B(n_1418),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1518),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1557),
.A2(n_1548),
.B(n_1490),
.Y(n_1621)
);

BUFx10_ASAP7_75t_L g1622 ( 
.A(n_1507),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1507),
.B(n_1351),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1572),
.B(n_1351),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1518),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1497),
.B(n_1408),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1578),
.B(n_1511),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1598),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1612),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1598),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1598),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_SL g1632 ( 
.A(n_1609),
.B(n_1388),
.C(n_1467),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1608),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1601),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1626),
.B(n_1511),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1626),
.B(n_1494),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1371),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1599),
.A2(n_1376),
.B1(n_1512),
.B2(n_1467),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1598),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1609),
.A2(n_1542),
.B1(n_1556),
.B2(n_1435),
.Y(n_1641)
);

NAND2x1_ASAP7_75t_L g1642 ( 
.A(n_1578),
.B(n_1340),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1576),
.A2(n_1533),
.B(n_1495),
.Y(n_1643)
);

NAND4xp25_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1520),
.C(n_1565),
.D(n_1506),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1599),
.A2(n_1533),
.B1(n_1435),
.B2(n_1554),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1593),
.B(n_1423),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1595),
.B(n_1344),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_SL g1648 ( 
.A1(n_1575),
.A2(n_1521),
.B(n_1493),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1601),
.Y(n_1649)
);

BUFx12f_ASAP7_75t_L g1650 ( 
.A(n_1602),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1593),
.B(n_1498),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1598),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1598),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1578),
.B(n_1623),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1602),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1494),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_R g1657 ( 
.A(n_1616),
.B(n_1409),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1576),
.A2(n_1578),
.B1(n_1583),
.B2(n_1586),
.Y(n_1658)
);

AOI222xp33_ASAP7_75t_L g1659 ( 
.A1(n_1614),
.A2(n_639),
.B1(n_596),
.B2(n_636),
.C1(n_496),
.C2(n_539),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1608),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1596),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1583),
.B(n_1529),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1600),
.A2(n_1508),
.B(n_1492),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1578),
.B(n_1340),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1619),
.A2(n_1621),
.B(n_1600),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1623),
.B(n_1549),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1596),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1602),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1608),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1670)
);

CKINVDCx14_ASAP7_75t_R g1671 ( 
.A(n_1585),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1596),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1582),
.B(n_1573),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_SL g1674 ( 
.A1(n_1614),
.A2(n_1586),
.B(n_1591),
.C(n_1582),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1594),
.A2(n_1471),
.B1(n_1434),
.B2(n_1448),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1574),
.B(n_1482),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1675),
.A2(n_1471),
.B1(n_429),
.B2(n_415),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1633),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1639),
.A2(n_1611),
.B1(n_1530),
.B2(n_1527),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1659),
.A2(n_1611),
.B(n_1448),
.C(n_1409),
.Y(n_1680)
);

OAI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1645),
.A2(n_1644),
.B(n_1658),
.C(n_1647),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1632),
.A2(n_429),
.B1(n_1577),
.B2(n_1594),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1627),
.A2(n_1575),
.B1(n_1584),
.B2(n_1592),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1644),
.A2(n_1353),
.B1(n_1464),
.B2(n_1463),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1627),
.A2(n_429),
.B1(n_1577),
.B2(n_1592),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1633),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1645),
.A2(n_535),
.B(n_539),
.C(n_532),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1627),
.B(n_1577),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1627),
.A2(n_1638),
.B1(n_1635),
.B2(n_1654),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1674),
.A2(n_1386),
.B1(n_1565),
.B2(n_478),
.C(n_482),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1641),
.A2(n_1524),
.B1(n_1615),
.B2(n_1486),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1666),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1636),
.B(n_1584),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1628),
.Y(n_1694)
);

OAI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1646),
.A2(n_545),
.B(n_549),
.C(n_544),
.Y(n_1695)
);

O2A1O1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1643),
.A2(n_1615),
.B(n_1580),
.C(n_544),
.Y(n_1696)
);

AOI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1665),
.A2(n_1619),
.B(n_1587),
.Y(n_1697)
);

OAI211xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1649),
.A2(n_1580),
.B(n_549),
.C(n_552),
.Y(n_1698)
);

AOI33xp33_ASAP7_75t_L g1699 ( 
.A1(n_1635),
.A2(n_566),
.A3(n_552),
.B1(n_567),
.B2(n_555),
.B3(n_545),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1660),
.Y(n_1700)
);

OAI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1651),
.A2(n_566),
.B(n_567),
.C(n_555),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1670),
.B(n_1634),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1627),
.A2(n_429),
.B1(n_1592),
.B2(n_1395),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1671),
.A2(n_1616),
.B1(n_1347),
.B2(n_1353),
.Y(n_1704)
);

INVx4_ASAP7_75t_L g1705 ( 
.A(n_1666),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1660),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1642),
.A2(n_1587),
.B(n_1589),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1662),
.A2(n_1499),
.B(n_1504),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1648),
.A2(n_590),
.B(n_595),
.C(n_581),
.Y(n_1709)
);

AOI222xp33_ASAP7_75t_L g1710 ( 
.A1(n_1648),
.A2(n_610),
.B1(n_590),
.B2(n_616),
.C1(n_595),
.C2(n_581),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1654),
.A2(n_1592),
.B1(n_1458),
.B2(n_1353),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1628),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1661),
.A2(n_1587),
.B(n_1603),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1636),
.B(n_1584),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1654),
.A2(n_1458),
.B1(n_1569),
.B2(n_1568),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1669),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1654),
.A2(n_1664),
.B1(n_1656),
.B2(n_1650),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1669),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1664),
.A2(n_1623),
.B1(n_1459),
.B2(n_1445),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1664),
.A2(n_1668),
.B1(n_1650),
.B2(n_1666),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1629),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1676),
.A2(n_484),
.B1(n_499),
.B2(n_481),
.C(n_475),
.Y(n_1723)
);

AOI222xp33_ASAP7_75t_L g1724 ( 
.A1(n_1668),
.A2(n_623),
.B1(n_610),
.B2(n_629),
.C1(n_627),
.C2(n_616),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1657),
.A2(n_1384),
.B1(n_1591),
.B2(n_1581),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1661),
.A2(n_1603),
.B(n_1606),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1673),
.A2(n_1347),
.B1(n_1581),
.B2(n_1562),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1630),
.A2(n_506),
.B1(n_507),
.B2(n_505),
.C(n_503),
.Y(n_1728)
);

A2O1A1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1642),
.A2(n_1581),
.B(n_1526),
.C(n_1606),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1629),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1629),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1664),
.A2(n_1584),
.B1(n_1581),
.B2(n_1622),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1630),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1655),
.A2(n_1373),
.B1(n_1623),
.B2(n_1421),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1655),
.A2(n_1484),
.B1(n_1396),
.B2(n_1474),
.C(n_629),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1666),
.A2(n_1367),
.B1(n_1623),
.B2(n_1622),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1637),
.B(n_1584),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1637),
.B(n_1590),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1663),
.A2(n_1526),
.B1(n_1588),
.B2(n_1574),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1663),
.B(n_1398),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1663),
.B(n_1585),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1640),
.Y(n_1742)
);

OAI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1640),
.A2(n_1589),
.B(n_1504),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1653),
.A2(n_1588),
.B1(n_636),
.B2(n_639),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1653),
.B(n_1436),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1631),
.A2(n_1453),
.B1(n_1391),
.B2(n_1442),
.Y(n_1746)
);

OA21x2_ASAP7_75t_L g1747 ( 
.A1(n_1667),
.A2(n_1603),
.B(n_1605),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1631),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1652),
.A2(n_1489),
.B1(n_1412),
.B2(n_1387),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1652),
.B(n_1590),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1652),
.A2(n_1622),
.B1(n_1621),
.B2(n_636),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1667),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1672),
.B(n_1590),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1672),
.A2(n_627),
.B1(n_635),
.B2(n_623),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1675),
.A2(n_636),
.B1(n_639),
.B2(n_596),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1675),
.A2(n_639),
.B1(n_596),
.B2(n_1380),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1675),
.A2(n_596),
.B1(n_1585),
.B2(n_1453),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1638),
.B(n_1585),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1665),
.A2(n_1621),
.B(n_1604),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1639),
.A2(n_1387),
.B1(n_1412),
.B2(n_1453),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1635),
.B(n_1590),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1753),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1688),
.B(n_1589),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1753),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1731),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1759),
.B(n_1428),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1693),
.B(n_1604),
.Y(n_1768)
);

OA21x2_ASAP7_75t_L g1769 ( 
.A1(n_1760),
.A2(n_1607),
.B(n_1605),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1702),
.B(n_1378),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1740),
.B(n_1604),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1694),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1724),
.A2(n_638),
.B1(n_640),
.B2(n_635),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1693),
.B(n_1604),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1747),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1714),
.B(n_1596),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1714),
.B(n_1596),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1719),
.B(n_1621),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1719),
.B(n_1579),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1762),
.B(n_1579),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1747),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1688),
.B(n_1579),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1747),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1677),
.A2(n_1756),
.B1(n_1757),
.B2(n_1680),
.C(n_1758),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1694),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1712),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1681),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1712),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1692),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1692),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1688),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1742),
.Y(n_1792)
);

OAI33xp33_ASAP7_75t_L g1793 ( 
.A1(n_1755),
.A2(n_664),
.A3(n_640),
.B1(n_667),
.B2(n_654),
.B3(n_638),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1742),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1733),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1749),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1692),
.B(n_1612),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1738),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1762),
.B(n_1579),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1688),
.B(n_1566),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1738),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1737),
.B(n_1552),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1683),
.B(n_1566),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1754),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1737),
.B(n_1754),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1705),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1691),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1713),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1725),
.B(n_1192),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1678),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1713),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1705),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1748),
.B(n_1566),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1684),
.B(n_1622),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1739),
.B(n_1612),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1748),
.B(n_1570),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1751),
.B(n_1552),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1705),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1715),
.A2(n_1689),
.B1(n_1736),
.B2(n_1735),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1751),
.B(n_1570),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1726),
.B(n_1552),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1732),
.B(n_1570),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1730),
.B(n_1685),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1722),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1730),
.B(n_1605),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1713),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1686),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1700),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1706),
.B(n_1618),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1717),
.B(n_1607),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1716),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1743),
.B(n_1607),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1718),
.B(n_1618),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1726),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1726),
.B(n_1546),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1707),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1745),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1699),
.B(n_1696),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1707),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1729),
.B(n_1618),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1729),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1750),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1697),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1699),
.B(n_1620),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1746),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1711),
.B(n_1546),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1697),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1703),
.B(n_1679),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1687),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1710),
.B(n_1620),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1752),
.B(n_1546),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1727),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1709),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1682),
.B(n_1620),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1721),
.B(n_1625),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1704),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1701),
.Y(n_1857)
);

AND2x4_ASAP7_75t_SL g1858 ( 
.A(n_1720),
.B(n_1625),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1708),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1734),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1695),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1708),
.B(n_1625),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1761),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1744),
.B(n_1613),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1698),
.B(n_1613),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1690),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1728),
.B(n_1613),
.Y(n_1867)
);

OAI222xp33_ASAP7_75t_L g1868 ( 
.A1(n_1723),
.A2(n_669),
.B1(n_664),
.B2(n_671),
.C1(n_667),
.C2(n_654),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1731),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1753),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1753),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1693),
.B(n_669),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1694),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1694),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1694),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1762),
.B(n_1494),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1731),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1693),
.B(n_671),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1753),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1702),
.B(n_508),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1753),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1719),
.B(n_1624),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1753),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1702),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1702),
.B(n_510),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1693),
.B(n_679),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1753),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1693),
.B(n_679),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1762),
.B(n_827),
.Y(n_1889)
);

BUFx2_ASAP7_75t_SL g1890 ( 
.A(n_1753),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1692),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1694),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1702),
.B(n_517),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1753),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1694),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1731),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1677),
.A2(n_1617),
.B1(n_1528),
.B2(n_1114),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1693),
.B(n_686),
.Y(n_1898)
);

OA21x2_ASAP7_75t_L g1899 ( 
.A1(n_1760),
.A2(n_1540),
.B(n_1553),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1693),
.B(n_686),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1724),
.A2(n_689),
.B1(n_700),
.B2(n_688),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1694),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1759),
.B(n_1354),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1693),
.B(n_688),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1694),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1762),
.B(n_827),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1753),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1693),
.B(n_689),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1762),
.B(n_832),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1753),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1772),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1805),
.B(n_832),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1785),
.Y(n_1913)
);

OAI31xp33_ASAP7_75t_L g1914 ( 
.A1(n_1868),
.A2(n_701),
.A3(n_700),
.B(n_834),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1790),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1884),
.B(n_1872),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_1790),
.Y(n_1917)
);

OAI33xp33_ASAP7_75t_L g1918 ( 
.A1(n_1866),
.A2(n_701),
.A3(n_534),
.B1(n_528),
.B2(n_537),
.B3(n_533),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1773),
.A2(n_1901),
.B1(n_1784),
.B2(n_1809),
.C(n_1838),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1891),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1808),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1891),
.Y(n_1922)
);

OAI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1787),
.A2(n_547),
.B1(n_548),
.B2(n_540),
.C(n_525),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1819),
.A2(n_1367),
.B1(n_1624),
.B2(n_834),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1786),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1805),
.B(n_836),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1882),
.B(n_836),
.Y(n_1927)
);

NOR2x1_ASAP7_75t_SL g1928 ( 
.A(n_1890),
.B(n_1617),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1808),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1882),
.B(n_838),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1848),
.A2(n_840),
.B(n_838),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1843),
.A2(n_846),
.B(n_840),
.Y(n_1932)
);

OAI321xp33_ASAP7_75t_L g1933 ( 
.A1(n_1848),
.A2(n_852),
.A3(n_846),
.B1(n_849),
.B2(n_818),
.C(n_1453),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1798),
.B(n_818),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1788),
.Y(n_1935)
);

OR2x6_ASAP7_75t_L g1936 ( 
.A(n_1764),
.B(n_1624),
.Y(n_1936)
);

NAND3xp33_ASAP7_75t_L g1937 ( 
.A(n_1841),
.B(n_852),
.C(n_849),
.Y(n_1937)
);

OAI321xp33_ASAP7_75t_L g1938 ( 
.A1(n_1863),
.A2(n_1221),
.A3(n_1216),
.B1(n_1236),
.B2(n_1229),
.C(n_1218),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1792),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1891),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1798),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1794),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1891),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1793),
.A2(n_554),
.B1(n_557),
.B2(n_551),
.Y(n_1944)
);

AOI21x1_ASAP7_75t_L g1945 ( 
.A1(n_1852),
.A2(n_1878),
.B(n_1872),
.Y(n_1945)
);

OAI33xp33_ASAP7_75t_L g1946 ( 
.A1(n_1861),
.A2(n_571),
.A3(n_561),
.B1(n_580),
.B2(n_565),
.B3(n_558),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1873),
.Y(n_1947)
);

BUFx3_ASAP7_75t_L g1948 ( 
.A(n_1891),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1882),
.B(n_1624),
.Y(n_1949)
);

OAI221xp5_ASAP7_75t_L g1950 ( 
.A1(n_1807),
.A2(n_599),
.B1(n_602),
.B2(n_592),
.C(n_588),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1874),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1878),
.B(n_1886),
.Y(n_1952)
);

OAI211xp5_ASAP7_75t_L g1953 ( 
.A1(n_1863),
.A2(n_1857),
.B(n_1849),
.C(n_1853),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1886),
.B(n_1624),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1811),
.Y(n_1955)
);

INVx4_ASAP7_75t_L g1956 ( 
.A(n_1889),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1814),
.A2(n_604),
.B1(n_606),
.B2(n_603),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1888),
.B(n_1519),
.Y(n_1958)
);

AOI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1767),
.A2(n_613),
.B1(n_615),
.B2(n_611),
.C(n_608),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1888),
.B(n_1898),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1875),
.Y(n_1961)
);

AOI211xp5_ASAP7_75t_L g1962 ( 
.A1(n_1897),
.A2(n_621),
.B(n_622),
.C(n_619),
.Y(n_1962)
);

AO21x2_ASAP7_75t_L g1963 ( 
.A1(n_1847),
.A2(n_1839),
.B(n_1836),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1898),
.B(n_1519),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1801),
.B(n_16),
.Y(n_1965)
);

OR2x6_ASAP7_75t_L g1966 ( 
.A(n_1764),
.B(n_1418),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1892),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1845),
.A2(n_637),
.B1(n_642),
.B2(n_634),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1853),
.A2(n_645),
.B1(n_648),
.B2(n_644),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1900),
.B(n_1519),
.Y(n_1970)
);

AO21x2_ASAP7_75t_L g1971 ( 
.A1(n_1847),
.A2(n_1229),
.B(n_1221),
.Y(n_1971)
);

OR2x6_ASAP7_75t_SL g1972 ( 
.A(n_1889),
.B(n_651),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1801),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1842),
.A2(n_659),
.B1(n_660),
.B2(n_656),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1811),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1895),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1804),
.B(n_16),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1859),
.A2(n_1867),
.B(n_1771),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1860),
.A2(n_663),
.B1(n_668),
.B2(n_662),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1770),
.A2(n_673),
.B1(n_674),
.B2(n_670),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1806),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1900),
.B(n_17),
.Y(n_1982)
);

AOI33xp33_ASAP7_75t_L g1983 ( 
.A1(n_1904),
.A2(n_17),
.A3(n_18),
.B1(n_21),
.B2(n_22),
.B3(n_23),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1860),
.A2(n_680),
.B(n_685),
.C(n_675),
.Y(n_1984)
);

OAI31xp33_ASAP7_75t_SL g1985 ( 
.A1(n_1903),
.A2(n_1782),
.A3(n_1851),
.B(n_1803),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1871),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1880),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1826),
.Y(n_1988)
);

OAI221xp5_ASAP7_75t_SL g1989 ( 
.A1(n_1885),
.A2(n_695),
.B1(n_702),
.B2(n_694),
.C(n_693),
.Y(n_1989)
);

OAI222xp33_ASAP7_75t_SL g1990 ( 
.A1(n_1893),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.C1(n_27),
.C2(n_28),
.Y(n_1990)
);

AOI221x1_ASAP7_75t_L g1991 ( 
.A1(n_1904),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.C(n_28),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1856),
.A2(n_707),
.B1(n_708),
.B2(n_704),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1804),
.B(n_29),
.Y(n_1993)
);

BUFx3_ASAP7_75t_L g1994 ( 
.A(n_1806),
.Y(n_1994)
);

OAI21xp33_ASAP7_75t_L g1995 ( 
.A1(n_1908),
.A2(n_711),
.B(n_709),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1902),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1908),
.B(n_29),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_1806),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1826),
.Y(n_1999)
);

AO21x2_ASAP7_75t_L g2000 ( 
.A1(n_1836),
.A2(n_1240),
.B(n_1236),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1834),
.A2(n_1276),
.B(n_1240),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1905),
.Y(n_2002)
);

AOI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1837),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.C(n_34),
.Y(n_2003)
);

AOI211xp5_ASAP7_75t_SL g2004 ( 
.A1(n_1803),
.A2(n_1068),
.B(n_1451),
.C(n_1383),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1812),
.B(n_31),
.Y(n_2005)
);

INVx5_ASAP7_75t_SL g2006 ( 
.A(n_1764),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1795),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1906),
.B(n_32),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1828),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1775),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1867),
.A2(n_1518),
.B1(n_1354),
.B2(n_1383),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1831),
.Y(n_2012)
);

OAI33xp33_ASAP7_75t_L g2013 ( 
.A1(n_1906),
.A2(n_35),
.A3(n_36),
.B1(n_37),
.B2(n_38),
.B3(n_39),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_1789),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1876),
.B(n_36),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1810),
.Y(n_2016)
);

OAI221xp5_ASAP7_75t_L g2017 ( 
.A1(n_1859),
.A2(n_1374),
.B1(n_1276),
.B2(n_1451),
.C(n_1465),
.Y(n_2017)
);

INVxp67_ASAP7_75t_SL g2018 ( 
.A(n_1775),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1909),
.B(n_1418),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1871),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1862),
.A2(n_1430),
.B(n_1068),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1781),
.Y(n_2022)
);

INVxp67_ASAP7_75t_SL g2023 ( 
.A(n_1781),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1876),
.B(n_38),
.Y(n_2024)
);

OAI33xp33_ASAP7_75t_L g2025 ( 
.A1(n_1909),
.A2(n_40),
.A3(n_43),
.B1(n_44),
.B2(n_45),
.B3(n_46),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1780),
.B(n_43),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1766),
.B(n_45),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1850),
.A2(n_1354),
.B1(n_1430),
.B2(n_1374),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1812),
.Y(n_2029)
);

INVx4_ASAP7_75t_L g2030 ( 
.A(n_1812),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1783),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1810),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1827),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1763),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1844),
.A2(n_1851),
.B1(n_1854),
.B2(n_1840),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1780),
.B(n_46),
.Y(n_2036)
);

AOI33xp33_ASAP7_75t_L g2037 ( 
.A1(n_1800),
.A2(n_1782),
.A3(n_1822),
.B1(n_1823),
.B2(n_1840),
.B3(n_1820),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1778),
.B(n_47),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1763),
.Y(n_2039)
);

INVxp67_ASAP7_75t_SL g2040 ( 
.A(n_1783),
.Y(n_2040)
);

CKINVDCx8_ASAP7_75t_R g2041 ( 
.A(n_1797),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1854),
.A2(n_1468),
.B1(n_1481),
.B2(n_1430),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1846),
.A2(n_1481),
.B1(n_1468),
.B2(n_49),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1765),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1778),
.B(n_47),
.Y(n_2045)
);

AO21x2_ASAP7_75t_L g2046 ( 
.A1(n_1834),
.A2(n_1280),
.B(n_922),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1799),
.B(n_1778),
.Y(n_2047)
);

AO21x2_ASAP7_75t_L g2048 ( 
.A1(n_1835),
.A2(n_1800),
.B(n_1821),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1799),
.B(n_48),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2048),
.B(n_1791),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2048),
.B(n_1791),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1941),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2037),
.B(n_1768),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1941),
.Y(n_2054)
);

INVxp67_ASAP7_75t_L g2055 ( 
.A(n_1912),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1973),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_1986),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1921),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_2047),
.B(n_1817),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2037),
.B(n_1768),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2035),
.B(n_1823),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1973),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1987),
.B(n_1818),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1916),
.B(n_1774),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2009),
.B(n_2012),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1936),
.B(n_1774),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_1915),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1978),
.B(n_1840),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1915),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1919),
.A2(n_1846),
.B1(n_1864),
.B2(n_1830),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1936),
.B(n_1776),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2034),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2026),
.B(n_1779),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2039),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2036),
.B(n_1779),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1936),
.B(n_1776),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2006),
.B(n_1777),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_1986),
.B(n_1817),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2016),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2032),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2006),
.B(n_1777),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2020),
.B(n_1802),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2049),
.B(n_1869),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1921),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1911),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_2014),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1966),
.B(n_1948),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1966),
.B(n_1818),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2020),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1929),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1929),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1913),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2006),
.B(n_1764),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1926),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1985),
.B(n_1877),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1966),
.B(n_2044),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1994),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2044),
.B(n_1890),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1945),
.B(n_1956),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1917),
.B(n_1813),
.Y(n_2100)
);

NAND2xp67_ASAP7_75t_L g2101 ( 
.A(n_1927),
.B(n_1862),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1956),
.B(n_1896),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1925),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1935),
.Y(n_2104)
);

HB1xp67_ASAP7_75t_L g2105 ( 
.A(n_2007),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_1955),
.B(n_1802),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2033),
.B(n_1815),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1920),
.B(n_1813),
.Y(n_2108)
);

NOR3xp33_ASAP7_75t_SL g2109 ( 
.A(n_1953),
.B(n_1881),
.C(n_1879),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1943),
.B(n_1816),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1955),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1981),
.B(n_1816),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1948),
.B(n_1907),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1981),
.B(n_1820),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_1975),
.B(n_1907),
.Y(n_2115)
);

AND2x2_ASAP7_75t_SL g2116 ( 
.A(n_1983),
.B(n_1858),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1994),
.B(n_1879),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1939),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1942),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_1975),
.B(n_1821),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1947),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_1988),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1998),
.B(n_1832),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1934),
.B(n_1822),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2029),
.B(n_1830),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2029),
.B(n_2038),
.Y(n_2126)
);

AND2x4_ASAP7_75t_L g2127 ( 
.A(n_1940),
.B(n_2030),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1988),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1934),
.B(n_1829),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1951),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1934),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_1940),
.B(n_1881),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_1972),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2045),
.B(n_1835),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2030),
.B(n_1883),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1999),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1999),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_2010),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_1962),
.B(n_1865),
.C(n_1855),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1961),
.B(n_1829),
.Y(n_2140)
);

NOR3xp33_ASAP7_75t_L g2141 ( 
.A(n_1923),
.B(n_1865),
.C(n_1855),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1967),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2010),
.B(n_1765),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1976),
.B(n_1829),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_2041),
.B(n_1797),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2022),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2022),
.B(n_1870),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2031),
.B(n_1870),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2031),
.B(n_1996),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2002),
.B(n_1894),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2018),
.B(n_1894),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1952),
.B(n_1833),
.Y(n_2152)
);

BUFx2_ASAP7_75t_L g2153 ( 
.A(n_1922),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2018),
.B(n_2023),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1960),
.B(n_1833),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2023),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2015),
.B(n_1833),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2040),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1963),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2024),
.B(n_1824),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1930),
.B(n_1883),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1963),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2040),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1965),
.B(n_1910),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1965),
.B(n_1910),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1965),
.B(n_1887),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1983),
.B(n_1797),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1949),
.B(n_1887),
.Y(n_2168)
);

NAND2x1p5_ASAP7_75t_L g2169 ( 
.A(n_2019),
.B(n_1864),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_1938),
.A2(n_1864),
.B(n_1858),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1977),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1958),
.B(n_1825),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1993),
.Y(n_2173)
);

INVx4_ASAP7_75t_L g2174 ( 
.A(n_2005),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1964),
.B(n_1796),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_1987),
.B(n_1796),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_2005),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2027),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1970),
.B(n_1825),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2005),
.B(n_1899),
.Y(n_2180)
);

NOR2xp67_ASAP7_75t_L g2181 ( 
.A(n_2028),
.B(n_1931),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_2011),
.B(n_1406),
.Y(n_2182)
);

AND2x4_ASAP7_75t_L g2183 ( 
.A(n_1928),
.B(n_48),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_1982),
.B(n_1769),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1932),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_1932),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2142),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2094),
.B(n_2011),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_2174),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_2089),
.Y(n_2190)
);

AOI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2141),
.A2(n_1990),
.B1(n_1980),
.B2(n_1918),
.C(n_1979),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_2174),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2105),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2159),
.Y(n_2194)
);

NAND2x1_ASAP7_75t_L g2195 ( 
.A(n_2089),
.B(n_2127),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2050),
.B(n_2051),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2050),
.B(n_1954),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_2055),
.B(n_1918),
.Y(n_2198)
);

NAND2x1p5_ASAP7_75t_L g2199 ( 
.A(n_2145),
.B(n_1769),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2053),
.B(n_2008),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2053),
.B(n_2008),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2072),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2159),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2060),
.B(n_2004),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2174),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2093),
.B(n_1997),
.Y(n_2206)
);

OAI21xp33_ASAP7_75t_L g2207 ( 
.A1(n_2070),
.A2(n_1980),
.B(n_1992),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_2067),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2156),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2051),
.B(n_2001),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2074),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2162),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2071),
.B(n_2001),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2162),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2071),
.B(n_2000),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2184),
.B(n_1899),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2079),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2080),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2085),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2184),
.B(n_1899),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2092),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2076),
.B(n_2000),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2076),
.B(n_1971),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2103),
.Y(n_2224)
);

INVx1_ASAP7_75t_SL g2225 ( 
.A(n_2086),
.Y(n_2225)
);

INVxp67_ASAP7_75t_SL g2226 ( 
.A(n_2158),
.Y(n_2226)
);

INVxp33_ASAP7_75t_SL g2227 ( 
.A(n_2133),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2104),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2118),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_2127),
.Y(n_2230)
);

INVx2_ASAP7_75t_SL g2231 ( 
.A(n_2127),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2119),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2121),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2130),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2060),
.B(n_2043),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2061),
.B(n_2043),
.Y(n_2236)
);

BUFx2_ASAP7_75t_L g2237 ( 
.A(n_2067),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2059),
.B(n_1971),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2059),
.B(n_1769),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2178),
.B(n_2042),
.Y(n_2240)
);

NOR2xp67_ASAP7_75t_SL g2241 ( 
.A(n_2133),
.B(n_2139),
.Y(n_2241)
);

OAI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2116),
.A2(n_1924),
.B1(n_2003),
.B2(n_1957),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2068),
.B(n_2042),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2052),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2166),
.B(n_1968),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2054),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2056),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2062),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2095),
.B(n_2021),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2166),
.B(n_2140),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2144),
.B(n_2164),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2149),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2073),
.B(n_1937),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2075),
.B(n_2046),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2082),
.Y(n_2255)
);

NAND2x1p5_ASAP7_75t_L g2256 ( 
.A(n_2145),
.B(n_1990),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2082),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2164),
.B(n_1995),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2123),
.B(n_1974),
.Y(n_2259)
);

INVxp67_ASAP7_75t_L g2260 ( 
.A(n_2099),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2154),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2165),
.B(n_1974),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2093),
.B(n_1984),
.Y(n_2263)
);

AOI21xp33_ASAP7_75t_L g2264 ( 
.A1(n_2099),
.A2(n_1950),
.B(n_1992),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2150),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2165),
.B(n_1991),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2150),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2154),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_2135),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2066),
.B(n_1959),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2087),
.B(n_49),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2078),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2078),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_2083),
.B(n_2017),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2065),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2122),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2115),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2115),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2148),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2148),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2151),
.Y(n_2281)
);

INVxp67_ASAP7_75t_SL g2282 ( 
.A(n_2163),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2151),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2066),
.B(n_1914),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2106),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2112),
.B(n_2114),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2122),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_2116),
.A2(n_1946),
.B1(n_2025),
.B2(n_2013),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2152),
.B(n_1969),
.Y(n_2289)
);

INVxp67_ASAP7_75t_SL g2290 ( 
.A(n_2122),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2176),
.B(n_1946),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2124),
.B(n_2160),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2143),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2143),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_2069),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2138),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2147),
.Y(n_2297)
);

A2O1A1Ixp33_ASAP7_75t_L g2298 ( 
.A1(n_2181),
.A2(n_1989),
.B(n_1944),
.C(n_1933),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2147),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2284),
.B(n_2200),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_2253),
.B(n_2292),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2201),
.B(n_2134),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2243),
.B(n_2157),
.Y(n_2303)
);

INVx2_ASAP7_75t_SL g2304 ( 
.A(n_2195),
.Y(n_2304)
);

BUFx2_ASAP7_75t_L g2305 ( 
.A(n_2208),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2198),
.B(n_2134),
.Y(n_2306)
);

NOR2x1_ASAP7_75t_L g2307 ( 
.A(n_2237),
.B(n_2183),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2202),
.Y(n_2308)
);

AND4x1_ASAP7_75t_L g2309 ( 
.A(n_2241),
.B(n_2109),
.C(n_2013),
.D(n_2025),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2194),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2249),
.B(n_2155),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2211),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2197),
.B(n_2108),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2194),
.Y(n_2314)
);

NAND2xp33_ASAP7_75t_L g2315 ( 
.A(n_2256),
.B(n_2167),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2209),
.Y(n_2316)
);

INVx1_ASAP7_75t_SL g2317 ( 
.A(n_2225),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2217),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2198),
.B(n_2171),
.Y(n_2319)
);

OAI221xp5_ASAP7_75t_L g2320 ( 
.A1(n_2264),
.A2(n_2167),
.B1(n_2170),
.B2(n_2173),
.C(n_2107),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_2227),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2203),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2197),
.B(n_2108),
.Y(n_2323)
);

INVx3_ASAP7_75t_SL g2324 ( 
.A(n_2271),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2227),
.B(n_2063),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2206),
.B(n_2110),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2206),
.B(n_2110),
.Y(n_2327)
);

OR2x2_ASAP7_75t_L g2328 ( 
.A(n_2204),
.B(n_2274),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2218),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2286),
.B(n_2112),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2259),
.B(n_2131),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_2209),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2219),
.Y(n_2333)
);

NOR2x1_ASAP7_75t_L g2334 ( 
.A(n_2263),
.B(n_2183),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2189),
.B(n_2114),
.Y(n_2335)
);

NAND5xp2_ASAP7_75t_SL g2336 ( 
.A(n_2288),
.B(n_2177),
.C(n_2126),
.D(n_2180),
.E(n_2125),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2266),
.B(n_2064),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2192),
.B(n_2205),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2271),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2203),
.Y(n_2340)
);

AOI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2207),
.A2(n_2182),
.B1(n_1944),
.B2(n_2183),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2212),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2212),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2230),
.B(n_2100),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2214),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2242),
.A2(n_2182),
.B1(n_2177),
.B2(n_2161),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2221),
.Y(n_2347)
);

INVx1_ASAP7_75t_SL g2348 ( 
.A(n_2295),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_2190),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2262),
.B(n_2101),
.Y(n_2350)
);

OAI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2256),
.A2(n_2169),
.B1(n_2129),
.B2(n_2087),
.Y(n_2351)
);

OAI221xp5_ASAP7_75t_L g2352 ( 
.A1(n_2191),
.A2(n_2102),
.B1(n_2169),
.B2(n_2069),
.C(n_2175),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2224),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2228),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2190),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2229),
.Y(n_2356)
);

NOR2x1_ASAP7_75t_L g2357 ( 
.A(n_2271),
.B(n_2153),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2214),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2232),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_R g2360 ( 
.A(n_2288),
.B(n_50),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2276),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2233),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2231),
.B(n_2087),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_R g2364 ( 
.A(n_2291),
.B(n_50),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2291),
.B(n_2168),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2230),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2234),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2235),
.B(n_2168),
.Y(n_2368)
);

INVxp67_ASAP7_75t_L g2369 ( 
.A(n_2188),
.Y(n_2369)
);

AO22x1_ASAP7_75t_L g2370 ( 
.A1(n_2260),
.A2(n_2057),
.B1(n_2126),
.B2(n_2097),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2270),
.B(n_2275),
.Y(n_2371)
);

AND2x2_ASAP7_75t_SL g2372 ( 
.A(n_2236),
.B(n_2088),
.Y(n_2372)
);

O2A1O1Ixp33_ASAP7_75t_SL g2373 ( 
.A1(n_2298),
.A2(n_2097),
.B(n_2120),
.C(n_2179),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2240),
.B(n_2172),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_R g2375 ( 
.A(n_2260),
.B(n_52),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2230),
.B(n_2172),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_2231),
.B(n_2180),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2245),
.B(n_2135),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2187),
.B(n_2096),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2250),
.B(n_2125),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2193),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2244),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2246),
.Y(n_2383)
);

INVx1_ASAP7_75t_SL g2384 ( 
.A(n_2258),
.Y(n_2384)
);

INVx1_ASAP7_75t_SL g2385 ( 
.A(n_2289),
.Y(n_2385)
);

NAND3xp33_ASAP7_75t_L g2386 ( 
.A(n_2298),
.B(n_2185),
.C(n_2096),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2276),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2251),
.B(n_2132),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2277),
.B(n_2132),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2247),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2278),
.B(n_2132),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2269),
.B(n_2077),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2281),
.B(n_2120),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2283),
.B(n_2077),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2248),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2255),
.Y(n_2396)
);

OA21x2_ASAP7_75t_L g2397 ( 
.A1(n_2290),
.A2(n_2084),
.B(n_2058),
.Y(n_2397)
);

INVxp67_ASAP7_75t_L g2398 ( 
.A(n_2226),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2199),
.Y(n_2399)
);

AOI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2223),
.A2(n_2081),
.B1(n_2088),
.B2(n_2135),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2287),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2226),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2279),
.B(n_2098),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_2254),
.B(n_2285),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2280),
.B(n_2098),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2265),
.B(n_2117),
.Y(n_2406)
);

A2O1A1Ixp33_ASAP7_75t_SL g2407 ( 
.A1(n_2369),
.A2(n_2210),
.B(n_2268),
.C(n_2261),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2316),
.Y(n_2408)
);

INVx1_ASAP7_75t_SL g2409 ( 
.A(n_2321),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2386),
.A2(n_2199),
.B1(n_2196),
.B2(n_2257),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2316),
.Y(n_2411)
);

AOI211x1_ASAP7_75t_L g2412 ( 
.A1(n_2309),
.A2(n_2196),
.B(n_2273),
.C(n_2272),
.Y(n_2412)
);

OAI221xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2341),
.A2(n_2210),
.B1(n_2282),
.B2(n_2220),
.C(n_2216),
.Y(n_2413)
);

INVxp67_ASAP7_75t_SL g2414 ( 
.A(n_2315),
.Y(n_2414)
);

INVxp67_ASAP7_75t_SL g2415 ( 
.A(n_2315),
.Y(n_2415)
);

OAI321xp33_ASAP7_75t_L g2416 ( 
.A1(n_2352),
.A2(n_2215),
.A3(n_2213),
.B1(n_2222),
.B2(n_2238),
.C(n_2239),
.Y(n_2416)
);

OAI21xp33_ASAP7_75t_L g2417 ( 
.A1(n_2360),
.A2(n_2215),
.B(n_2213),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2321),
.B(n_2325),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2349),
.Y(n_2419)
);

OAI22xp33_ASAP7_75t_L g2420 ( 
.A1(n_2320),
.A2(n_2290),
.B1(n_2186),
.B2(n_2252),
.Y(n_2420)
);

HB1xp67_ASAP7_75t_L g2421 ( 
.A(n_2349),
.Y(n_2421)
);

OAI221xp5_ASAP7_75t_SL g2422 ( 
.A1(n_2341),
.A2(n_2267),
.B1(n_2294),
.B2(n_2297),
.C(n_2293),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2325),
.B(n_2299),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2332),
.Y(n_2424)
);

OAI321xp33_ASAP7_75t_L g2425 ( 
.A1(n_2351),
.A2(n_2296),
.A3(n_2287),
.B1(n_2146),
.B2(n_2137),
.C(n_2136),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2326),
.B(n_2117),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2332),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2372),
.A2(n_2088),
.B1(n_2117),
.B2(n_2296),
.Y(n_2428)
);

AOI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2372),
.A2(n_2186),
.B1(n_2113),
.B2(n_2084),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2346),
.A2(n_2186),
.B1(n_2113),
.B2(n_2138),
.Y(n_2430)
);

INVx1_ASAP7_75t_SL g2431 ( 
.A(n_2364),
.Y(n_2431)
);

NAND4xp25_ASAP7_75t_L g2432 ( 
.A(n_2328),
.B(n_2113),
.C(n_2090),
.D(n_2091),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2308),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2336),
.A2(n_2138),
.B1(n_2090),
.B2(n_2091),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2312),
.Y(n_2435)
);

OR2x2_ASAP7_75t_L g2436 ( 
.A(n_2301),
.B(n_2058),
.Y(n_2436)
);

AOI21xp33_ASAP7_75t_L g2437 ( 
.A1(n_2319),
.A2(n_2128),
.B(n_2111),
.Y(n_2437)
);

OR2x2_ASAP7_75t_L g2438 ( 
.A(n_2371),
.B(n_2111),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2318),
.Y(n_2439)
);

INVxp33_ASAP7_75t_L g2440 ( 
.A(n_2364),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2385),
.B(n_2128),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2329),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2333),
.Y(n_2443)
);

AOI321xp33_ASAP7_75t_L g2444 ( 
.A1(n_2334),
.A2(n_2146),
.A3(n_2137),
.B1(n_2136),
.B2(n_55),
.C(n_57),
.Y(n_2444)
);

AOI21xp33_ASAP7_75t_L g2445 ( 
.A1(n_2350),
.A2(n_52),
.B(n_53),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2365),
.B(n_54),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2384),
.B(n_54),
.Y(n_2447)
);

AOI21xp33_ASAP7_75t_L g2448 ( 
.A1(n_2307),
.A2(n_55),
.B(n_57),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2317),
.B(n_920),
.Y(n_2449)
);

CKINVDCx20_ASAP7_75t_R g2450 ( 
.A(n_2339),
.Y(n_2450)
);

HB1xp67_ASAP7_75t_L g2451 ( 
.A(n_2355),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2347),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2353),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2300),
.B(n_60),
.Y(n_2454)
);

O2A1O1Ixp33_ASAP7_75t_L g2455 ( 
.A1(n_2360),
.A2(n_64),
.B(n_60),
.C(n_61),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2348),
.B(n_61),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2327),
.B(n_65),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2354),
.Y(n_2458)
);

INVxp67_ASAP7_75t_SL g2459 ( 
.A(n_2355),
.Y(n_2459)
);

NAND2x1_ASAP7_75t_SL g2460 ( 
.A(n_2357),
.B(n_66),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2366),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2303),
.B(n_67),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2306),
.B(n_2305),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2398),
.Y(n_2464)
);

NAND4xp25_ASAP7_75t_L g2465 ( 
.A(n_2373),
.B(n_69),
.C(n_67),
.D(n_68),
.Y(n_2465)
);

AOI31xp33_ASAP7_75t_L g2466 ( 
.A1(n_2373),
.A2(n_70),
.A3(n_68),
.B(n_69),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2324),
.B(n_70),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2324),
.B(n_71),
.Y(n_2468)
);

NOR2xp67_ASAP7_75t_L g2469 ( 
.A(n_2304),
.B(n_74),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2338),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2335),
.B(n_76),
.Y(n_2471)
);

AOI21xp33_ASAP7_75t_SL g2472 ( 
.A1(n_2370),
.A2(n_77),
.B(n_78),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2380),
.B(n_77),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_2331),
.A2(n_79),
.B(n_80),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2375),
.B(n_922),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2375),
.B(n_80),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2356),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2378),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_2478)
);

NAND3xp33_ASAP7_75t_L g2479 ( 
.A(n_2398),
.B(n_82),
.C(n_86),
.Y(n_2479)
);

NAND3x1_ASAP7_75t_L g2480 ( 
.A(n_2366),
.B(n_87),
.C(n_88),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2368),
.B(n_89),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2313),
.B(n_90),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2378),
.B(n_90),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2381),
.B(n_91),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2359),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2362),
.Y(n_2486)
);

OAI322xp33_ASAP7_75t_L g2487 ( 
.A1(n_2402),
.A2(n_91),
.A3(n_92),
.B1(n_96),
.B2(n_98),
.C1(n_99),
.C2(n_100),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2374),
.B(n_96),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2363),
.Y(n_2489)
);

NOR2xp67_ASAP7_75t_L g2490 ( 
.A(n_2400),
.B(n_98),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2419),
.Y(n_2491)
);

NAND2x1p5_ASAP7_75t_L g2492 ( 
.A(n_2469),
.B(n_2363),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2419),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2412),
.B(n_2367),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2474),
.B(n_2311),
.Y(n_2495)
);

OAI21xp33_ASAP7_75t_L g2496 ( 
.A1(n_2417),
.A2(n_2337),
.B(n_2379),
.Y(n_2496)
);

AOI211xp5_ASAP7_75t_SL g2497 ( 
.A1(n_2466),
.A2(n_2396),
.B(n_2363),
.C(n_2392),
.Y(n_2497)
);

AOI321xp33_ASAP7_75t_L g2498 ( 
.A1(n_2414),
.A2(n_2302),
.A3(n_2382),
.B1(n_2390),
.B2(n_2395),
.C(n_2383),
.Y(n_2498)
);

OR2x2_ASAP7_75t_L g2499 ( 
.A(n_2463),
.B(n_2404),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2431),
.B(n_2323),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2421),
.Y(n_2501)
);

AOI21xp33_ASAP7_75t_SL g2502 ( 
.A1(n_2440),
.A2(n_2396),
.B(n_2399),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2468),
.B(n_2330),
.Y(n_2503)
);

AOI22xp33_ASAP7_75t_L g2504 ( 
.A1(n_2465),
.A2(n_2377),
.B1(n_2391),
.B2(n_2389),
.Y(n_2504)
);

BUFx2_ASAP7_75t_L g2505 ( 
.A(n_2460),
.Y(n_2505)
);

NOR2x1_ASAP7_75t_L g2506 ( 
.A(n_2450),
.B(n_2397),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2421),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2415),
.A2(n_2405),
.B(n_2403),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_L g2509 ( 
.A(n_2451),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2415),
.A2(n_2344),
.B1(n_2377),
.B2(n_2376),
.Y(n_2510)
);

AOI322xp5_ASAP7_75t_L g2511 ( 
.A1(n_2476),
.A2(n_2377),
.A3(n_2388),
.B1(n_2406),
.B2(n_2310),
.C1(n_2345),
.C2(n_2314),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_2409),
.B(n_2394),
.Y(n_2512)
);

AOI21xp33_ASAP7_75t_L g2513 ( 
.A1(n_2455),
.A2(n_2314),
.B(n_2310),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2470),
.B(n_2489),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2418),
.B(n_2393),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_2467),
.B(n_2361),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2472),
.B(n_2361),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2426),
.B(n_2387),
.Y(n_2518)
);

INVxp67_ASAP7_75t_SL g2519 ( 
.A(n_2480),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2451),
.Y(n_2520)
);

AOI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_2448),
.A2(n_2401),
.B(n_2387),
.Y(n_2521)
);

NAND3xp33_ASAP7_75t_L g2522 ( 
.A(n_2444),
.B(n_2340),
.C(n_2322),
.Y(n_2522)
);

OAI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2490),
.A2(n_2397),
.B1(n_2401),
.B2(n_2340),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2459),
.Y(n_2524)
);

NAND3xp33_ASAP7_75t_SL g2525 ( 
.A(n_2455),
.B(n_2342),
.C(n_2322),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2462),
.B(n_2342),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2423),
.B(n_2343),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2459),
.Y(n_2528)
);

AOI22xp5_ASAP7_75t_L g2529 ( 
.A1(n_2410),
.A2(n_2345),
.B1(n_2358),
.B2(n_2343),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2464),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2464),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2408),
.B(n_2358),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2457),
.B(n_2397),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2471),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2473),
.B(n_99),
.Y(n_2535)
);

AOI21xp33_ASAP7_75t_L g2536 ( 
.A1(n_2479),
.A2(n_100),
.B(n_101),
.Y(n_2536)
);

OAI21xp33_ASAP7_75t_L g2537 ( 
.A1(n_2413),
.A2(n_101),
.B(n_103),
.Y(n_2537)
);

NOR3xp33_ASAP7_75t_L g2538 ( 
.A(n_2413),
.B(n_1280),
.C(n_104),
.Y(n_2538)
);

OAI21xp5_ASAP7_75t_SL g2539 ( 
.A1(n_2445),
.A2(n_104),
.B(n_105),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2428),
.B(n_105),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2420),
.A2(n_923),
.B1(n_927),
.B2(n_917),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2411),
.B(n_106),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2424),
.Y(n_2543)
);

XOR2x2_ASAP7_75t_L g2544 ( 
.A(n_2478),
.B(n_108),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2461),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2454),
.B(n_2484),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2427),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2407),
.A2(n_112),
.B(n_115),
.Y(n_2548)
);

AOI22xp33_ASAP7_75t_L g2549 ( 
.A1(n_2420),
.A2(n_923),
.B1(n_927),
.B2(n_917),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2433),
.Y(n_2550)
);

INVxp67_ASAP7_75t_L g2551 ( 
.A(n_2475),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2435),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2439),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2442),
.Y(n_2554)
);

OAI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2422),
.A2(n_116),
.B1(n_112),
.B2(n_115),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2416),
.B(n_1406),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2482),
.B(n_117),
.Y(n_2557)
);

AND2x2_ASAP7_75t_SL g2558 ( 
.A(n_2483),
.B(n_118),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2429),
.B(n_119),
.Y(n_2559)
);

OAI21xp33_ASAP7_75t_SL g2560 ( 
.A1(n_2432),
.A2(n_120),
.B(n_121),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2447),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2438),
.B(n_120),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2446),
.B(n_121),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2456),
.B(n_2441),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2488),
.B(n_122),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2481),
.B(n_2443),
.Y(n_2566)
);

AO22x1_ASAP7_75t_L g2567 ( 
.A1(n_2430),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2436),
.B(n_126),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2509),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2519),
.B(n_2497),
.Y(n_2570)
);

AOI21xp33_ASAP7_75t_L g2571 ( 
.A1(n_2537),
.A2(n_2453),
.B(n_2452),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2497),
.B(n_2458),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2505),
.B(n_2477),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2524),
.Y(n_2574)
);

CKINVDCx20_ASAP7_75t_R g2575 ( 
.A(n_2544),
.Y(n_2575)
);

INVx4_ASAP7_75t_L g2576 ( 
.A(n_2542),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2528),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2534),
.B(n_2485),
.Y(n_2578)
);

OR2x2_ASAP7_75t_L g2579 ( 
.A(n_2500),
.B(n_2486),
.Y(n_2579)
);

NOR3xp33_ASAP7_75t_SL g2580 ( 
.A(n_2525),
.B(n_2555),
.C(n_2560),
.Y(n_2580)
);

XOR2xp5_ASAP7_75t_L g2581 ( 
.A(n_2492),
.B(n_2449),
.Y(n_2581)
);

OAI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2548),
.A2(n_2555),
.B1(n_2495),
.B2(n_2492),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2491),
.Y(n_2583)
);

AND3x2_ASAP7_75t_L g2584 ( 
.A(n_2538),
.B(n_2487),
.C(n_2425),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2493),
.Y(n_2585)
);

NAND2xp33_ASAP7_75t_R g2586 ( 
.A(n_2540),
.B(n_127),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2501),
.Y(n_2587)
);

OR2x2_ASAP7_75t_L g2588 ( 
.A(n_2561),
.B(n_2437),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2561),
.B(n_2434),
.Y(n_2589)
);

NOR3xp33_ASAP7_75t_SL g2590 ( 
.A(n_2512),
.B(n_128),
.C(n_130),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2494),
.B(n_2522),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2558),
.B(n_131),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2542),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2551),
.B(n_2546),
.Y(n_2594)
);

AOI21xp33_ASAP7_75t_SL g2595 ( 
.A1(n_2536),
.A2(n_131),
.B(n_134),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2507),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2515),
.B(n_135),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2520),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2494),
.B(n_137),
.Y(n_2599)
);

NOR3xp33_ASAP7_75t_L g2600 ( 
.A(n_2502),
.B(n_137),
.C(n_138),
.Y(n_2600)
);

INVx1_ASAP7_75t_SL g2601 ( 
.A(n_2506),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2530),
.Y(n_2602)
);

INVxp67_ASAP7_75t_L g2603 ( 
.A(n_2517),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2564),
.B(n_138),
.Y(n_2604)
);

OAI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2539),
.A2(n_139),
.B(n_141),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2566),
.B(n_141),
.Y(n_2606)
);

BUFx2_ASAP7_75t_L g2607 ( 
.A(n_2531),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2568),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2526),
.Y(n_2609)
);

INVxp67_ASAP7_75t_L g2610 ( 
.A(n_2514),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2516),
.B(n_142),
.Y(n_2611)
);

NOR2x1_ASAP7_75t_L g2612 ( 
.A(n_2539),
.B(n_143),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2562),
.Y(n_2613)
);

AOI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2523),
.A2(n_143),
.B(n_144),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2532),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2532),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2567),
.B(n_146),
.Y(n_2617)
);

OAI222xp33_ASAP7_75t_L g2618 ( 
.A1(n_2523),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.C1(n_152),
.C2(n_153),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2503),
.B(n_148),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2559),
.B(n_150),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2543),
.Y(n_2621)
);

NAND2xp33_ASAP7_75t_L g2622 ( 
.A(n_2499),
.B(n_152),
.Y(n_2622)
);

OAI21xp33_ASAP7_75t_L g2623 ( 
.A1(n_2496),
.A2(n_2511),
.B(n_2510),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_2527),
.B(n_154),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2547),
.Y(n_2625)
);

AOI211xp5_ASAP7_75t_L g2626 ( 
.A1(n_2582),
.A2(n_2513),
.B(n_2556),
.C(n_2508),
.Y(n_2626)
);

INVxp67_ASAP7_75t_SL g2627 ( 
.A(n_2622),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2607),
.Y(n_2628)
);

NAND3xp33_ASAP7_75t_L g2629 ( 
.A(n_2580),
.B(n_2498),
.C(n_2513),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2593),
.B(n_2504),
.Y(n_2630)
);

NOR3xp33_ASAP7_75t_L g2631 ( 
.A(n_2570),
.B(n_2563),
.C(n_2565),
.Y(n_2631)
);

NAND5xp2_ASAP7_75t_L g2632 ( 
.A(n_2623),
.B(n_2529),
.C(n_2521),
.D(n_2553),
.E(n_2552),
.Y(n_2632)
);

AND2x4_ASAP7_75t_L g2633 ( 
.A(n_2576),
.B(n_2545),
.Y(n_2633)
);

NAND4xp25_ASAP7_75t_L g2634 ( 
.A(n_2591),
.B(n_2554),
.C(n_2550),
.D(n_2535),
.Y(n_2634)
);

AOI211xp5_ASAP7_75t_L g2635 ( 
.A1(n_2582),
.A2(n_2533),
.B(n_2557),
.C(n_2518),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2576),
.Y(n_2636)
);

NOR4xp25_ASAP7_75t_L g2637 ( 
.A(n_2601),
.B(n_2549),
.C(n_2541),
.D(n_156),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2612),
.B(n_154),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2569),
.Y(n_2639)
);

NAND3xp33_ASAP7_75t_L g2640 ( 
.A(n_2600),
.B(n_157),
.C(n_159),
.Y(n_2640)
);

AOI222xp33_ASAP7_75t_L g2641 ( 
.A1(n_2572),
.A2(n_161),
.B1(n_164),
.B2(n_166),
.C1(n_168),
.C2(n_169),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2613),
.Y(n_2642)
);

NOR3xp33_ASAP7_75t_L g2643 ( 
.A(n_2599),
.B(n_168),
.C(n_169),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2608),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2575),
.B(n_171),
.Y(n_2645)
);

INVxp67_ASAP7_75t_L g2646 ( 
.A(n_2586),
.Y(n_2646)
);

NOR3xp33_ASAP7_75t_L g2647 ( 
.A(n_2594),
.B(n_172),
.C(n_174),
.Y(n_2647)
);

NOR3xp33_ASAP7_75t_L g2648 ( 
.A(n_2603),
.B(n_175),
.C(n_177),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2574),
.Y(n_2649)
);

INVxp67_ASAP7_75t_L g2650 ( 
.A(n_2617),
.Y(n_2650)
);

NAND4xp25_ASAP7_75t_L g2651 ( 
.A(n_2589),
.B(n_175),
.C(n_178),
.D(n_179),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2610),
.B(n_180),
.Y(n_2652)
);

AOI221x1_ASAP7_75t_L g2653 ( 
.A1(n_2614),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.C(n_185),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_SL g2654 ( 
.A(n_2618),
.B(n_2592),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2577),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2602),
.Y(n_2656)
);

NAND3xp33_ASAP7_75t_L g2657 ( 
.A(n_2584),
.B(n_181),
.C(n_182),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2605),
.B(n_185),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2605),
.B(n_2619),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2601),
.B(n_917),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2590),
.B(n_941),
.Y(n_2661)
);

INVx2_ASAP7_75t_SL g2662 ( 
.A(n_2579),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2583),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2606),
.B(n_188),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2585),
.Y(n_2665)
);

NOR3xp33_ASAP7_75t_L g2666 ( 
.A(n_2611),
.B(n_188),
.C(n_190),
.Y(n_2666)
);

NOR3x1_ASAP7_75t_L g2667 ( 
.A(n_2573),
.B(n_191),
.C(n_192),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2628),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2629),
.A2(n_2581),
.B1(n_2609),
.B2(n_2598),
.Y(n_2669)
);

OAI211xp5_ASAP7_75t_SL g2670 ( 
.A1(n_2626),
.A2(n_2571),
.B(n_2588),
.C(n_2587),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2630),
.B(n_2597),
.Y(n_2671)
);

AOI21xp33_ASAP7_75t_L g2672 ( 
.A1(n_2646),
.A2(n_2578),
.B(n_2596),
.Y(n_2672)
);

AOI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2657),
.A2(n_2604),
.B1(n_2620),
.B2(n_2616),
.Y(n_2673)
);

AOI211xp5_ASAP7_75t_L g2674 ( 
.A1(n_2632),
.A2(n_2595),
.B(n_2615),
.C(n_2621),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2646),
.B(n_2624),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2627),
.B(n_2625),
.Y(n_2676)
);

INVx2_ASAP7_75t_SL g2677 ( 
.A(n_2633),
.Y(n_2677)
);

OAI221xp5_ASAP7_75t_SL g2678 ( 
.A1(n_2635),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.C(n_196),
.Y(n_2678)
);

O2A1O1Ixp33_ASAP7_75t_L g2679 ( 
.A1(n_2659),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_2679)
);

NAND3xp33_ASAP7_75t_L g2680 ( 
.A(n_2654),
.B(n_197),
.C(n_198),
.Y(n_2680)
);

OAI31xp33_ASAP7_75t_L g2681 ( 
.A1(n_2640),
.A2(n_2651),
.A3(n_2643),
.B(n_2666),
.Y(n_2681)
);

XOR2x2_ASAP7_75t_L g2682 ( 
.A(n_2645),
.B(n_201),
.Y(n_2682)
);

A2O1A1Ixp33_ASAP7_75t_L g2683 ( 
.A1(n_2643),
.A2(n_202),
.B(n_203),
.C(n_204),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2662),
.Y(n_2684)
);

NAND4xp25_ASAP7_75t_L g2685 ( 
.A(n_2631),
.B(n_203),
.C(n_204),
.D(n_205),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_SL g2686 ( 
.A(n_2641),
.B(n_206),
.C(n_207),
.D(n_208),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2633),
.B(n_206),
.Y(n_2687)
);

OAI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2637),
.A2(n_207),
.B(n_209),
.Y(n_2688)
);

OAI211xp5_ASAP7_75t_L g2689 ( 
.A1(n_2653),
.A2(n_209),
.B(n_211),
.C(n_212),
.Y(n_2689)
);

AOI222xp33_ASAP7_75t_L g2690 ( 
.A1(n_2650),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.C1(n_217),
.C2(n_219),
.Y(n_2690)
);

AO22x2_ASAP7_75t_L g2691 ( 
.A1(n_2636),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_2631),
.A2(n_941),
.B1(n_942),
.B2(n_946),
.Y(n_2692)
);

NAND3xp33_ASAP7_75t_SL g2693 ( 
.A(n_2666),
.B(n_220),
.C(n_221),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2647),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_R g2695 ( 
.A(n_2638),
.B(n_223),
.Y(n_2695)
);

AOI221xp5_ASAP7_75t_L g2696 ( 
.A1(n_2634),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.C(n_227),
.Y(n_2696)
);

AOI211xp5_ASAP7_75t_L g2697 ( 
.A1(n_2648),
.A2(n_229),
.B(n_231),
.C(n_232),
.Y(n_2697)
);

XNOR2x1_ASAP7_75t_L g2698 ( 
.A(n_2658),
.B(n_229),
.Y(n_2698)
);

AOI222xp33_ASAP7_75t_L g2699 ( 
.A1(n_2639),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.C1(n_238),
.C2(n_240),
.Y(n_2699)
);

INVxp67_ASAP7_75t_L g2700 ( 
.A(n_2677),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2687),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2676),
.Y(n_2702)
);

NOR2x1_ASAP7_75t_L g2703 ( 
.A(n_2680),
.B(n_2652),
.Y(n_2703)
);

NOR2x1_ASAP7_75t_L g2704 ( 
.A(n_2693),
.B(n_2660),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_2688),
.B(n_2644),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2691),
.Y(n_2706)
);

OAI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2670),
.A2(n_2642),
.B(n_2665),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2684),
.B(n_2671),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2690),
.B(n_2667),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2695),
.Y(n_2710)
);

NAND2xp33_ASAP7_75t_SL g2711 ( 
.A(n_2698),
.B(n_2664),
.Y(n_2711)
);

OR2x6_ASAP7_75t_L g2712 ( 
.A(n_2675),
.B(n_2661),
.Y(n_2712)
);

NOR2x1_ASAP7_75t_L g2713 ( 
.A(n_2685),
.B(n_2689),
.Y(n_2713)
);

OA22x2_ASAP7_75t_L g2714 ( 
.A1(n_2669),
.A2(n_2663),
.B1(n_2656),
.B2(n_2655),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2674),
.A2(n_2649),
.B1(n_235),
.B2(n_241),
.Y(n_2715)
);

AOI322xp5_ASAP7_75t_L g2716 ( 
.A1(n_2672),
.A2(n_233),
.A3(n_241),
.B1(n_242),
.B2(n_243),
.C1(n_247),
.C2(n_252),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_R g2717 ( 
.A(n_2686),
.B(n_2668),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2678),
.B(n_2673),
.Y(n_2718)
);

OAI211xp5_ASAP7_75t_SL g2719 ( 
.A1(n_2681),
.A2(n_946),
.B(n_943),
.C(n_942),
.Y(n_2719)
);

OAI21xp33_ASAP7_75t_SL g2720 ( 
.A1(n_2673),
.A2(n_265),
.B(n_269),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2682),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2683),
.B(n_271),
.Y(n_2722)
);

NAND3xp33_ASAP7_75t_L g2723 ( 
.A(n_2707),
.B(n_2696),
.C(n_2679),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2702),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2708),
.Y(n_2725)
);

BUFx3_ASAP7_75t_L g2726 ( 
.A(n_2712),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2700),
.B(n_2694),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_R g2728 ( 
.A(n_2711),
.B(n_2697),
.Y(n_2728)
);

NAND3xp33_ASAP7_75t_L g2729 ( 
.A(n_2715),
.B(n_2713),
.C(n_2706),
.Y(n_2729)
);

AOI222xp33_ASAP7_75t_L g2730 ( 
.A1(n_2705),
.A2(n_2699),
.B1(n_2692),
.B2(n_274),
.C1(n_276),
.C2(n_279),
.Y(n_2730)
);

NOR3x1_ASAP7_75t_L g2731 ( 
.A(n_2709),
.B(n_272),
.C(n_273),
.Y(n_2731)
);

BUFx2_ASAP7_75t_L g2732 ( 
.A(n_2712),
.Y(n_2732)
);

NAND4xp75_ASAP7_75t_L g2733 ( 
.A(n_2703),
.B(n_282),
.C(n_285),
.D(n_286),
.Y(n_2733)
);

OAI322xp33_ASAP7_75t_L g2734 ( 
.A1(n_2714),
.A2(n_290),
.A3(n_291),
.B1(n_298),
.B2(n_300),
.C1(n_302),
.C2(n_303),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2710),
.B(n_309),
.Y(n_2735)
);

NAND3x1_ASAP7_75t_SL g2736 ( 
.A(n_2704),
.B(n_312),
.C(n_316),
.Y(n_2736)
);

NOR3xp33_ASAP7_75t_L g2737 ( 
.A(n_2721),
.B(n_946),
.C(n_943),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_SL g2738 ( 
.A(n_2717),
.B(n_1406),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2712),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2701),
.Y(n_2740)
);

NOR3xp33_ASAP7_75t_SL g2741 ( 
.A(n_2729),
.B(n_2720),
.C(n_2722),
.Y(n_2741)
);

NOR3xp33_ASAP7_75t_SL g2742 ( 
.A(n_2723),
.B(n_2727),
.C(n_2738),
.Y(n_2742)
);

OAI221xp5_ASAP7_75t_L g2743 ( 
.A1(n_2732),
.A2(n_2718),
.B1(n_2716),
.B2(n_2719),
.C(n_903),
.Y(n_2743)
);

NAND4xp25_ASAP7_75t_L g2744 ( 
.A(n_2726),
.B(n_318),
.C(n_319),
.D(n_320),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_2728),
.A2(n_900),
.B1(n_903),
.B2(n_934),
.Y(n_2745)
);

NAND3xp33_ASAP7_75t_SL g2746 ( 
.A(n_2730),
.B(n_323),
.C(n_325),
.Y(n_2746)
);

NAND4xp25_ASAP7_75t_L g2747 ( 
.A(n_2725),
.B(n_326),
.C(n_329),
.D(n_338),
.Y(n_2747)
);

NOR3xp33_ASAP7_75t_L g2748 ( 
.A(n_2739),
.B(n_2740),
.C(n_2724),
.Y(n_2748)
);

AOI221xp5_ASAP7_75t_L g2749 ( 
.A1(n_2734),
.A2(n_903),
.B1(n_900),
.B2(n_348),
.C(n_352),
.Y(n_2749)
);

NAND3xp33_ASAP7_75t_L g2750 ( 
.A(n_2737),
.B(n_934),
.C(n_940),
.Y(n_2750)
);

OAI222xp33_ASAP7_75t_R g2751 ( 
.A1(n_2731),
.A2(n_343),
.B1(n_346),
.B2(n_354),
.C1(n_360),
.C2(n_361),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2748),
.B(n_2735),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2742),
.Y(n_2753)
);

NOR3xp33_ASAP7_75t_SL g2754 ( 
.A(n_2743),
.B(n_2733),
.C(n_2736),
.Y(n_2754)
);

CKINVDCx16_ASAP7_75t_R g2755 ( 
.A(n_2746),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_2741),
.Y(n_2756)
);

CKINVDCx12_ASAP7_75t_R g2757 ( 
.A(n_2751),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_2750),
.B(n_2735),
.Y(n_2758)
);

AND3x1_ASAP7_75t_L g2759 ( 
.A(n_2754),
.B(n_2749),
.C(n_2745),
.Y(n_2759)
);

NAND3xp33_ASAP7_75t_L g2760 ( 
.A(n_2756),
.B(n_2747),
.C(n_2744),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2752),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2758),
.Y(n_2762)
);

OAI221xp5_ASAP7_75t_L g2763 ( 
.A1(n_2753),
.A2(n_363),
.B1(n_364),
.B2(n_368),
.C(n_370),
.Y(n_2763)
);

OAI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2757),
.A2(n_1005),
.B(n_992),
.Y(n_2764)
);

INVx1_ASAP7_75t_SL g2765 ( 
.A(n_2761),
.Y(n_2765)
);

CKINVDCx20_ASAP7_75t_R g2766 ( 
.A(n_2760),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2762),
.A2(n_2755),
.B1(n_992),
.B2(n_1005),
.Y(n_2767)
);

AOI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2764),
.A2(n_947),
.B(n_940),
.Y(n_2768)
);

CKINVDCx20_ASAP7_75t_R g2769 ( 
.A(n_2766),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2765),
.Y(n_2770)
);

AOI222xp33_ASAP7_75t_L g2771 ( 
.A1(n_2770),
.A2(n_2763),
.B1(n_2759),
.B2(n_2767),
.C1(n_2768),
.C2(n_378),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2769),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2772),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2771),
.Y(n_2774)
);

OAI21xp33_ASAP7_75t_SL g2775 ( 
.A1(n_2773),
.A2(n_386),
.B(n_387),
.Y(n_2775)
);

OAI221xp5_ASAP7_75t_R g2776 ( 
.A1(n_2774),
.A2(n_388),
.B1(n_389),
.B2(n_391),
.C(n_392),
.Y(n_2776)
);

AOI221xp5_ASAP7_75t_L g2777 ( 
.A1(n_2775),
.A2(n_947),
.B1(n_940),
.B2(n_396),
.C(n_397),
.Y(n_2777)
);

AOI211xp5_ASAP7_75t_L g2778 ( 
.A1(n_2777),
.A2(n_2776),
.B(n_395),
.C(n_399),
.Y(n_2778)
);


endmodule