module fake_ariane_2036_n_1390 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_381, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_382, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1390);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1390;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_96),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_275),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_170),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_113),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_104),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_292),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_103),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_2),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_79),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_182),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_261),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_196),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_171),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_341),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_251),
.B(n_181),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_125),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_333),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_225),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_165),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_180),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_62),
.B(n_50),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_304),
.B(n_187),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_29),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_155),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_158),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_217),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_255),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_354),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_256),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_246),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_259),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_66),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_48),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_343),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_195),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_184),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_272),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_145),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_250),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_200),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_179),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_293),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_173),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_85),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_58),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_268),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_319),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_198),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_55),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_280),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_276),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_282),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_93),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_254),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_222),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_186),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_191),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_54),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_174),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_73),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_185),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_224),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_190),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_146),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_253),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_262),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_51),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_8),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_88),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_278),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_291),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_8),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_147),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_286),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_263),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_183),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_218),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_235),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_337),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_376),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_69),
.B(n_88),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_99),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_153),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_63),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_359),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_143),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_12),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_177),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_317),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_351),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_204),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_188),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_233),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_156),
.B(n_296),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_363),
.B(n_377),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_334),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_312),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_53),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_151),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_101),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_205),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_37),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_68),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_19),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_207),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_199),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_318),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_290),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_220),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_365),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_22),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_277),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_7),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_162),
.B(n_160),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_144),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_208),
.B(n_344),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_360),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_236),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_273),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_32),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_201),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_12),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_166),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_335),
.B(n_357),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_18),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_20),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_169),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_13),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_81),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_106),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_382),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_117),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_219),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_345),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_232),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_118),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_281),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_192),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_300),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_238),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_84),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_294),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_303),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_226),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_267),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_202),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_306),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_309),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_352),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_116),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_279),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_370),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_197),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_2),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_64),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_210),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_26),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_260),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_36),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_3),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_375),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_349),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_106),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_264),
.B(n_20),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_265),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_383),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_86),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_298),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_159),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_231),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_307),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_194),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_161),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_36),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_68),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_284),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_243),
.Y(n_566)
);

CKINVDCx14_ASAP7_75t_R g567 ( 
.A(n_203),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_54),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_90),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_436),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_417),
.B(n_0),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_417),
.B(n_0),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_385),
.A2(n_1),
.B(n_3),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_1),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_511),
.B(n_4),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_528),
.B(n_5),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_511),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_436),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_569),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_519),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_436),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_456),
.B(n_5),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_386),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_440),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_388),
.B(n_9),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_440),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_468),
.B(n_10),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_456),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_530),
.B(n_10),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_492),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_390),
.B(n_11),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_546),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_411),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_411),
.Y(n_599)
);

OA21x2_ASAP7_75t_L g600 ( 
.A1(n_391),
.A2(n_11),
.B(n_13),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_394),
.B(n_14),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_14),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_433),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_444),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_434),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_399),
.B(n_424),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_406),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_384),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_444),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_440),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_389),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_445),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_502),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_442),
.Y(n_615)
);

OA21x2_ASAP7_75t_L g616 ( 
.A1(n_398),
.A2(n_15),
.B(n_16),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_449),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_445),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_491),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_543),
.B(n_15),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_543),
.B(n_16),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_463),
.Y(n_622)
);

BUFx8_ASAP7_75t_SL g623 ( 
.A(n_493),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_402),
.B(n_17),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_457),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_440),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_535),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_392),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_463),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_473),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_535),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_468),
.A2(n_123),
.B(n_122),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_535),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_393),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_397),
.Y(n_636)
);

BUFx12f_ASAP7_75t_L g637 ( 
.A(n_397),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_514),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_403),
.B(n_407),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_545),
.Y(n_642)
);

OA21x2_ASAP7_75t_L g643 ( 
.A1(n_412),
.A2(n_17),
.B(n_18),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_498),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_420),
.Y(n_646)
);

AOI22x1_ASAP7_75t_SL g647 ( 
.A1(n_416),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_518),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_525),
.Y(n_649)
);

BUFx8_ASAP7_75t_SL g650 ( 
.A(n_419),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_556),
.B(n_21),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_413),
.B(n_23),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_429),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_438),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_446),
.B(n_24),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_545),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_544),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_552),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_579),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_579),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_579),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_644),
.B(n_485),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_606),
.B(n_512),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_580),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_610),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_580),
.Y(n_667)
);

AND3x2_ASAP7_75t_L g668 ( 
.A(n_591),
.B(n_395),
.C(n_387),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_578),
.B(n_446),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_606),
.B(n_529),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_580),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_580),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_610),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_547),
.Y(n_674)
);

AO21x2_ASAP7_75t_L g675 ( 
.A1(n_588),
.A2(n_553),
.B(n_430),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_570),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_587),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_607),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_655),
.B(n_558),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_584),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_570),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_587),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_627),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_627),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_627),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_570),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_570),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_584),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_589),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_604),
.B(n_561),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_608),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_581),
.B(n_498),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_589),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_589),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_589),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_641),
.B(n_547),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_609),
.B(n_567),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_612),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_613),
.Y(n_701)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_641),
.A2(n_418),
.B(n_405),
.Y(n_702)
);

BUFx6f_ASAP7_75t_SL g703 ( 
.A(n_651),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_578),
.B(n_582),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_650),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_626),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_626),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_628),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_635),
.B(n_646),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_593),
.A2(n_504),
.B1(n_523),
.B2(n_474),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_629),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_697),
.B(n_618),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_664),
.A2(n_572),
.B1(n_577),
.B2(n_575),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_675),
.B(n_666),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_701),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_663),
.B(n_637),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_704),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_674),
.B(n_654),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_622),
.Y(n_720)
);

INVxp33_ASAP7_75t_SL g721 ( 
.A(n_679),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_666),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_670),
.B(n_577),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_691),
.B(n_593),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_692),
.B(n_596),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_673),
.B(n_573),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_677),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_692),
.B(n_573),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_669),
.B(n_630),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_673),
.B(n_576),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_698),
.B(n_576),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_675),
.B(n_592),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_700),
.B(n_572),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_704),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_675),
.B(n_590),
.Y(n_735)
);

NAND2x1p5_ASAP7_75t_L g736 ( 
.A(n_700),
.B(n_620),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_709),
.B(n_585),
.C(n_590),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_592),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_710),
.A2(n_586),
.B1(n_653),
.B2(n_591),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_680),
.B(n_594),
.C(n_588),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_710),
.B(n_599),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_677),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_703),
.A2(n_621),
.B1(n_620),
.B2(n_651),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_686),
.B(n_602),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_703),
.A2(n_567),
.B1(n_601),
.B2(n_594),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_693),
.B(n_601),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_702),
.B(n_624),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_705),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_705),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_683),
.B(n_652),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_668),
.B(n_598),
.Y(n_751)
);

AND2x6_ASAP7_75t_L g752 ( 
.A(n_689),
.B(n_470),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_702),
.B(n_652),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_684),
.B(n_583),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_684),
.B(n_597),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_685),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_682),
.B(n_571),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_694),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_694),
.B(n_427),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_695),
.B(n_431),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_695),
.B(n_448),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_659),
.B(n_598),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_682),
.B(n_595),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_699),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_706),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_660),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_660),
.A2(n_447),
.B1(n_461),
.B2(n_458),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_661),
.A2(n_564),
.B1(n_471),
.B2(n_487),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_661),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_662),
.B(n_455),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_685),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_685),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_665),
.B(n_460),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_665),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_667),
.B(n_671),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_726),
.B(n_454),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_747),
.A2(n_633),
.B(n_505),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_753),
.A2(n_735),
.B(n_731),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_735),
.A2(n_688),
.B(n_687),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_SL g780 ( 
.A(n_737),
.B(n_409),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_724),
.B(n_466),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_723),
.A2(n_537),
.B1(n_499),
.B2(n_462),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_725),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_771),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_734),
.A2(n_563),
.B(n_615),
.C(n_603),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_722),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_754),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_713),
.B(n_481),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_738),
.B(n_617),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_715),
.A2(n_600),
.B(n_574),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_719),
.B(n_500),
.C(n_489),
.Y(n_791)
);

NOR2xp67_ASAP7_75t_L g792 ( 
.A(n_717),
.B(n_614),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_720),
.B(n_508),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_755),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_748),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_741),
.B(n_614),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_729),
.B(n_516),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_730),
.A2(n_638),
.B(n_648),
.C(n_625),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_714),
.A2(n_465),
.B(n_479),
.C(n_464),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_732),
.A2(n_671),
.B(n_667),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_738),
.B(n_605),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_728),
.A2(n_562),
.B1(n_486),
.B2(n_490),
.Y(n_802)
);

AOI21x1_ASAP7_75t_L g803 ( 
.A1(n_775),
.A2(n_678),
.B(n_672),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_770),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_750),
.A2(n_600),
.B(n_574),
.Y(n_805)
);

O2A1O1Ixp5_ASAP7_75t_L g806 ( 
.A1(n_746),
.A2(n_496),
.B(n_497),
.C(n_480),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_744),
.A2(n_643),
.B(n_616),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_740),
.A2(n_643),
.B(n_616),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_758),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_771),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_742),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_775),
.A2(n_696),
.B(n_681),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_SL g813 ( 
.A1(n_733),
.A2(n_507),
.B(n_510),
.C(n_506),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_742),
.A2(n_711),
.B(n_707),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_765),
.A2(n_526),
.B(n_524),
.Y(n_815)
);

BUFx2_ASAP7_75t_SL g816 ( 
.A(n_749),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_743),
.A2(n_536),
.B(n_538),
.C(n_531),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_716),
.B(n_517),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_539),
.Y(n_819)
);

AOI21x1_ASAP7_75t_L g820 ( 
.A1(n_759),
.A2(n_711),
.B(n_707),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_762),
.B(n_548),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_762),
.B(n_549),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_751),
.B(n_631),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_764),
.B(n_611),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_768),
.A2(n_658),
.B(n_657),
.C(n_640),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_745),
.B(n_568),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_757),
.A2(n_712),
.B(n_550),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_727),
.A2(n_554),
.B(n_541),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_763),
.B(n_396),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_721),
.B(n_483),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_759),
.A2(n_418),
.B(n_405),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_760),
.A2(n_559),
.B(n_560),
.C(n_555),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_767),
.B(n_739),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_774),
.B(n_605),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_771),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_772),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_752),
.B(n_400),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_760),
.B(n_647),
.C(n_645),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_752),
.B(n_404),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_752),
.B(n_408),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_761),
.A2(n_773),
.B(n_770),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_761),
.A2(n_773),
.B(n_766),
.C(n_769),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_752),
.B(n_414),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_752),
.A2(n_410),
.B(n_401),
.Y(n_844)
);

CKINVDCx10_ASAP7_75t_R g845 ( 
.A(n_756),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_725),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_735),
.A2(n_649),
.B(n_639),
.C(n_522),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_723),
.A2(n_422),
.B1(n_423),
.B2(n_415),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_726),
.B(n_425),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_723),
.B(n_619),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_747),
.A2(n_503),
.B(n_484),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_725),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_747),
.A2(n_676),
.B(n_533),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_726),
.B(n_426),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_747),
.A2(n_557),
.B(n_551),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_748),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_747),
.A2(n_432),
.B(n_428),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_771),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_747),
.A2(n_513),
.B(n_439),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_722),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_738),
.B(n_619),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_721),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_747),
.A2(n_441),
.B(n_435),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_726),
.B(n_443),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_747),
.A2(n_451),
.B(n_450),
.Y(n_865)
);

OAI321xp33_ASAP7_75t_L g866 ( 
.A1(n_737),
.A2(n_545),
.A3(n_634),
.B1(n_642),
.B2(n_632),
.C(n_629),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_747),
.A2(n_453),
.B(n_452),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_747),
.A2(n_467),
.B(n_459),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_726),
.B(n_469),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_747),
.A2(n_475),
.B(n_472),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_737),
.A2(n_478),
.B1(n_482),
.B2(n_477),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_718),
.B(n_690),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_771),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_726),
.B(n_488),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_777),
.A2(n_126),
.B(n_124),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_776),
.B(n_494),
.Y(n_876)
);

OAI21xp33_ASAP7_75t_L g877 ( 
.A1(n_781),
.A2(n_501),
.B(n_495),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_788),
.B(n_849),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_850),
.B(n_527),
.C(n_520),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_854),
.A2(n_869),
.B1(n_874),
.B2(n_864),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_792),
.B(n_532),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_851),
.A2(n_632),
.B(n_629),
.Y(n_882)
);

AO32x2_ASAP7_75t_L g883 ( 
.A1(n_831),
.A2(n_27),
.A3(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_SL g884 ( 
.A1(n_804),
.A2(n_540),
.B(n_534),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_796),
.B(n_542),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_862),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_786),
.Y(n_887)
);

AO31x2_ASAP7_75t_L g888 ( 
.A1(n_842),
.A2(n_634),
.A3(n_642),
.B(n_632),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_861),
.Y(n_889)
);

NOR2x1_ASAP7_75t_L g890 ( 
.A(n_816),
.B(n_634),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_852),
.B(n_623),
.Y(n_891)
);

OAI21x1_ASAP7_75t_L g892 ( 
.A1(n_800),
.A2(n_128),
.B(n_127),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_807),
.A2(n_130),
.B(n_129),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_783),
.B(n_623),
.Y(n_894)
);

OA21x2_ASAP7_75t_L g895 ( 
.A1(n_808),
.A2(n_566),
.B(n_565),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_805),
.A2(n_690),
.B(n_132),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_845),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_779),
.A2(n_690),
.B(n_133),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_846),
.B(n_29),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_860),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_784),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_803),
.A2(n_690),
.B(n_656),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_830),
.B(n_30),
.Y(n_903)
);

O2A1O1Ixp5_ASAP7_75t_L g904 ( 
.A1(n_780),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_904)
);

AO31x2_ASAP7_75t_L g905 ( 
.A1(n_855),
.A2(n_642),
.A3(n_34),
.B(n_31),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_857),
.A2(n_134),
.B(n_131),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_812),
.A2(n_136),
.B(n_135),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_865),
.A2(n_138),
.B(n_137),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_833),
.A2(n_37),
.B1(n_33),
.B2(n_35),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_799),
.A2(n_39),
.B1(n_35),
.B2(n_38),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_853),
.A2(n_820),
.B(n_841),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_795),
.Y(n_912)
);

AOI221x1_ASAP7_75t_L g913 ( 
.A1(n_859),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.C(n_41),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_834),
.B(n_789),
.Y(n_914)
);

AO31x2_ASAP7_75t_L g915 ( 
.A1(n_832),
.A2(n_43),
.A3(n_41),
.B(n_42),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_793),
.B(n_797),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_787),
.B(n_794),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_861),
.B(n_801),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_823),
.B(n_42),
.Y(n_919)
);

AO31x2_ASAP7_75t_L g920 ( 
.A1(n_817),
.A2(n_827),
.A3(n_828),
.B(n_826),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_847),
.A2(n_814),
.B(n_863),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_856),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_809),
.B(n_43),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_815),
.B(n_44),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_L g925 ( 
.A(n_782),
.B(n_819),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_791),
.B(n_45),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_844),
.A2(n_140),
.B(n_139),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_821),
.B(n_45),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_867),
.A2(n_142),
.B(n_141),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_823),
.B(n_46),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_824),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_848),
.A2(n_47),
.B(n_48),
.Y(n_932)
);

OAI21x1_ASAP7_75t_SL g933 ( 
.A1(n_785),
.A2(n_47),
.B(n_49),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_829),
.B(n_50),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_811),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_871),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_822),
.B(n_51),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_784),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_836),
.A2(n_56),
.B1(n_52),
.B2(n_53),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_868),
.A2(n_870),
.B(n_818),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_798),
.B(n_52),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_802),
.B(n_56),
.Y(n_942)
);

AO31x2_ASAP7_75t_L g943 ( 
.A1(n_837),
.A2(n_59),
.A3(n_57),
.B(n_58),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_838),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_806),
.A2(n_60),
.B(n_57),
.C(n_59),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_784),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_810),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_872),
.A2(n_840),
.B(n_839),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_843),
.A2(n_149),
.B(n_148),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_825),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_810),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_813),
.B(n_63),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_835),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_866),
.A2(n_152),
.B(n_150),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_835),
.A2(n_64),
.B(n_65),
.Y(n_955)
);

AO22x2_ASAP7_75t_L g956 ( 
.A1(n_858),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_873),
.B(n_67),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_776),
.B(n_70),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_778),
.A2(n_157),
.B(n_154),
.Y(n_959)
);

AO31x2_ASAP7_75t_L g960 ( 
.A1(n_831),
.A2(n_72),
.A3(n_70),
.B(n_71),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_861),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_831),
.A2(n_75),
.A3(n_73),
.B(n_74),
.Y(n_962)
);

BUFx6f_ASAP7_75t_SL g963 ( 
.A(n_795),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_831),
.A2(n_76),
.A3(n_74),
.B(n_75),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_776),
.B(n_76),
.Y(n_965)
);

AO31x2_ASAP7_75t_L g966 ( 
.A1(n_831),
.A2(n_79),
.A3(n_77),
.B(n_78),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_776),
.A2(n_80),
.B(n_77),
.C(n_78),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_784),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_790),
.A2(n_164),
.B(n_163),
.Y(n_969)
);

AOI22x1_ASAP7_75t_L g970 ( 
.A1(n_778),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_778),
.A2(n_168),
.B(n_167),
.Y(n_971)
);

OA22x2_ASAP7_75t_L g972 ( 
.A1(n_861),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_796),
.B(n_83),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_786),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_777),
.A2(n_175),
.B(n_172),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_777),
.A2(n_178),
.B(n_176),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_786),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_795),
.Y(n_978)
);

AO31x2_ASAP7_75t_L g979 ( 
.A1(n_831),
.A2(n_87),
.A3(n_85),
.B(n_86),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_776),
.B(n_87),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_776),
.B(n_89),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_845),
.Y(n_982)
);

AND2x6_ASAP7_75t_SL g983 ( 
.A(n_850),
.B(n_89),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_776),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_778),
.A2(n_193),
.B(n_189),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_776),
.B(n_91),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_831),
.A2(n_94),
.A3(n_95),
.B(n_96),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_SL g988 ( 
.A1(n_785),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.C(n_99),
.Y(n_988)
);

CKINVDCx6p67_ASAP7_75t_R g989 ( 
.A(n_845),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_776),
.B(n_97),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_850),
.B(n_98),
.C(n_100),
.Y(n_991)
);

NOR2x1_ASAP7_75t_L g992 ( 
.A(n_816),
.B(n_101),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_861),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_796),
.B(n_102),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_776),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_845),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_784),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_776),
.B(n_105),
.Y(n_998)
);

NOR2xp67_ASAP7_75t_L g999 ( 
.A(n_862),
.B(n_206),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_789),
.B(n_105),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_914),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_938),
.Y(n_1002)
);

OA21x2_ASAP7_75t_L g1003 ( 
.A1(n_911),
.A2(n_896),
.B(n_921),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_918),
.B(n_107),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_882),
.A2(n_211),
.B(n_209),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_973),
.B(n_994),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_887),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_922),
.B(n_212),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_940),
.A2(n_310),
.A3(n_381),
.B(n_380),
.Y(n_1009)
);

CKINVDCx6p67_ASAP7_75t_R g1010 ( 
.A(n_989),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_875),
.A2(n_214),
.B(n_213),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_878),
.A2(n_880),
.B(n_917),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_889),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_898),
.A2(n_216),
.B(n_215),
.Y(n_1014)
);

OAI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_936),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_958),
.A2(n_110),
.B(n_111),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_963),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_916),
.B(n_112),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_931),
.B(n_112),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_946),
.Y(n_1020)
);

NAND2x1p5_ASAP7_75t_L g1021 ( 
.A(n_978),
.B(n_221),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_900),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_R g1023 ( 
.A(n_897),
.B(n_113),
.Y(n_1023)
);

OA21x2_ASAP7_75t_L g1024 ( 
.A1(n_892),
.A2(n_227),
.B(n_223),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_908),
.A2(n_229),
.B(n_228),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_SL g1026 ( 
.A(n_894),
.B(n_114),
.Y(n_1026)
);

OA21x2_ASAP7_75t_L g1027 ( 
.A1(n_948),
.A2(n_315),
.B(n_379),
.Y(n_1027)
);

BUFx2_ASAP7_75t_SL g1028 ( 
.A(n_1000),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_961),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_912),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_903),
.A2(n_891),
.B1(n_993),
.B2(n_932),
.Y(n_1031)
);

CKINVDCx16_ASAP7_75t_R g1032 ( 
.A(n_982),
.Y(n_1032)
);

OA21x2_ASAP7_75t_L g1033 ( 
.A1(n_985),
.A2(n_314),
.B(n_378),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_953),
.B(n_230),
.Y(n_1034)
);

AO31x2_ASAP7_75t_L g1035 ( 
.A1(n_913),
.A2(n_954),
.A3(n_929),
.B(n_906),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_996),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1000),
.B(n_115),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_974),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_975),
.A2(n_316),
.B(n_374),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_919),
.Y(n_1040)
);

BUFx2_ASAP7_75t_SL g1041 ( 
.A(n_999),
.Y(n_1041)
);

OR2x6_ASAP7_75t_SL g1042 ( 
.A(n_984),
.B(n_115),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_977),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_991),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_972),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_SL g1046 ( 
.A(n_969),
.B(n_234),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_965),
.A2(n_986),
.B(n_981),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_885),
.B(n_237),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_925),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_1049)
);

INVx5_ASAP7_75t_L g1050 ( 
.A(n_901),
.Y(n_1050)
);

AO32x2_ASAP7_75t_L g1051 ( 
.A1(n_910),
.A2(n_242),
.A3(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_976),
.A2(n_248),
.B(n_249),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_907),
.A2(n_252),
.B(n_257),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_928),
.B(n_258),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_876),
.B(n_266),
.Y(n_1055)
);

XOR2xp5_ASAP7_75t_L g1056 ( 
.A(n_944),
.B(n_269),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_935),
.B(n_270),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_893),
.A2(n_271),
.B(n_274),
.Y(n_1058)
);

BUFx8_ASAP7_75t_L g1059 ( 
.A(n_930),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_956),
.A2(n_942),
.B1(n_899),
.B2(n_952),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_SL g1061 ( 
.A1(n_909),
.A2(n_283),
.B1(n_285),
.B2(n_287),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_983),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_956),
.B(n_288),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_926),
.A2(n_289),
.B(n_295),
.C(n_297),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_937),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_1065)
);

BUFx2_ASAP7_75t_SL g1066 ( 
.A(n_901),
.Y(n_1066)
);

AOI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_990),
.A2(n_305),
.B(n_308),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_947),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_SL g1069 ( 
.A(n_992),
.B(n_311),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_998),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_SL g1071 ( 
.A1(n_980),
.A2(n_323),
.B(n_324),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_888),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_941),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_888),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_949),
.A2(n_325),
.A3(n_326),
.B(n_327),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_959),
.A2(n_328),
.A3(n_330),
.B(n_331),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_336),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_890),
.B(n_373),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_SL g1079 ( 
.A1(n_970),
.A2(n_338),
.B1(n_339),
.B2(n_342),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_934),
.A2(n_346),
.B(n_347),
.C(n_348),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_884),
.B(n_350),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_968),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_968),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_927),
.A2(n_355),
.B(n_356),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_923),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_877),
.A2(n_879),
.B1(n_995),
.B2(n_895),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_988),
.B(n_372),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_997),
.B(n_361),
.Y(n_1088)
);

OAI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_939),
.A2(n_371),
.B1(n_362),
.B2(n_364),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_997),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_920),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_904),
.A2(n_366),
.B(n_367),
.Y(n_1092)
);

CKINVDCx11_ASAP7_75t_R g1093 ( 
.A(n_883),
.Y(n_1093)
);

OA21x2_ASAP7_75t_L g1094 ( 
.A1(n_945),
.A2(n_368),
.B(n_369),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_933),
.A2(n_955),
.B1(n_957),
.B2(n_951),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_950),
.Y(n_1096)
);

AOI221xp5_ASAP7_75t_SL g1097 ( 
.A1(n_967),
.A2(n_883),
.B1(n_915),
.B2(n_943),
.C(n_962),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_888),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_905),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_943),
.B(n_960),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_960),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_964),
.A2(n_966),
.B(n_979),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_964),
.A2(n_966),
.B(n_979),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_964),
.A2(n_966),
.B1(n_979),
.B2(n_987),
.Y(n_1104)
);

OAI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_987),
.A2(n_850),
.B1(n_833),
.B2(n_903),
.C(n_846),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_987),
.A2(n_800),
.B(n_911),
.Y(n_1106)
);

INVx8_ASAP7_75t_L g1107 ( 
.A(n_963),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_914),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_911),
.A2(n_800),
.B(n_902),
.Y(n_1109)
);

AOI22x1_ASAP7_75t_L g1110 ( 
.A1(n_940),
.A2(n_908),
.B1(n_898),
.B2(n_896),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_SL g1111 ( 
.A1(n_908),
.A2(n_985),
.B(n_971),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_878),
.A2(n_778),
.B(n_880),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_924),
.A2(n_721),
.B(n_776),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_914),
.B(n_931),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_911),
.A2(n_896),
.B(n_800),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_911),
.A2(n_800),
.B(n_902),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_911),
.A2(n_800),
.B(n_902),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_886),
.B(n_862),
.C(n_705),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1007),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1108),
.B(n_1040),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1012),
.B(n_1073),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_1111),
.A2(n_1100),
.B(n_1074),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1068),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_SL g1124 ( 
.A(n_1028),
.Y(n_1124)
);

OA21x2_ASAP7_75t_L g1125 ( 
.A1(n_1106),
.A2(n_1097),
.B(n_1102),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1109),
.A2(n_1117),
.B(n_1116),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1022),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1038),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1043),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1112),
.A2(n_1096),
.B(n_1018),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1010),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1015),
.A2(n_1045),
.B1(n_1105),
.B2(n_1026),
.C(n_1113),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_SL g1133 ( 
.A(n_1028),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1111),
.A2(n_1098),
.B(n_1072),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1006),
.B(n_1037),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1114),
.B(n_1004),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1114),
.B(n_1019),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1083),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1091),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1013),
.B(n_1029),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1063),
.A2(n_1060),
.B1(n_1093),
.B2(n_1016),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1107),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1063),
.A2(n_1031),
.B1(n_1061),
.B2(n_1047),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1055),
.A2(n_1025),
.B(n_1014),
.C(n_1044),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1091),
.Y(n_1145)
);

AND2x4_ASAP7_75t_SL g1146 ( 
.A(n_1020),
.B(n_1036),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1050),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1090),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1050),
.Y(n_1149)
);

AOI21xp33_ASAP7_75t_L g1150 ( 
.A1(n_1110),
.A2(n_1086),
.B(n_1101),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1085),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1030),
.B(n_1054),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1082),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1042),
.B(n_1048),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1032),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1066),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1008),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1099),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1099),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1107),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1059),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1050),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1041),
.B(n_1095),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1002),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1017),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1001),
.A2(n_1081),
.B1(n_1069),
.B2(n_1059),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1089),
.A2(n_1087),
.B1(n_1056),
.B2(n_1071),
.C(n_1104),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1021),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1118),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1057),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1034),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1062),
.B(n_1081),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1041),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1051),
.B(n_1077),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1088),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1051),
.B(n_1103),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1078),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1003),
.A2(n_1115),
.B(n_1033),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1009),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1009),
.Y(n_1180)
);

AO32x2_ASAP7_75t_L g1181 ( 
.A1(n_1051),
.A2(n_1003),
.A3(n_1046),
.B1(n_1076),
.B2(n_1005),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1064),
.A2(n_1080),
.B(n_1049),
.C(n_1067),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1092),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_SL g1184 ( 
.A(n_1005),
.B(n_1033),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1035),
.B(n_1079),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1075),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1075),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1075),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1035),
.B(n_1094),
.Y(n_1189)
);

CKINVDCx11_ASAP7_75t_R g1190 ( 
.A(n_1023),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1076),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1115),
.A2(n_1035),
.A3(n_1027),
.B(n_1053),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1011),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1039),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1052),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1084),
.B(n_1058),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1058),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1149),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1119),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1127),
.Y(n_1201)
);

AND2x2_ASAP7_75t_SL g1202 ( 
.A(n_1174),
.B(n_1141),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1135),
.B(n_1024),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1136),
.B(n_1137),
.Y(n_1204)
);

BUFx8_ASAP7_75t_L g1205 ( 
.A(n_1161),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1120),
.B(n_1024),
.Y(n_1206)
);

AND2x2_ASAP7_75t_SL g1207 ( 
.A(n_1141),
.B(n_1143),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1139),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1132),
.A2(n_1143),
.B1(n_1154),
.B2(n_1166),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1154),
.B(n_1138),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1146),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1139),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1128),
.B(n_1129),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1172),
.B(n_1151),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1148),
.B(n_1140),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1150),
.A2(n_1184),
.B(n_1179),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1156),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1121),
.B(n_1130),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1156),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1163),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1169),
.B(n_1123),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1170),
.B(n_1124),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1155),
.B(n_1166),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1155),
.B(n_1164),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1145),
.Y(n_1227)
);

NAND2x1_ASAP7_75t_L g1228 ( 
.A(n_1177),
.B(n_1168),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1145),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1158),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1160),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1171),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1132),
.A2(n_1194),
.B1(n_1167),
.B2(n_1176),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1159),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1162),
.B(n_1147),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1167),
.B(n_1122),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1133),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1133),
.B(n_1173),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1125),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1125),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1157),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1134),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1175),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1186),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1173),
.B(n_1144),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1165),
.B(n_1144),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1131),
.B(n_1190),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1131),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1187),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1185),
.B(n_1188),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1194),
.B(n_1185),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1191),
.B(n_1189),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1193),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1190),
.B(n_1181),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1207),
.A2(n_1180),
.B1(n_1197),
.B2(n_1198),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1208),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1253),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1251),
.B(n_1181),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1251),
.B(n_1178),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1200),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1244),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1201),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1246),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1249),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1223),
.B(n_1182),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1211),
.B(n_1182),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1213),
.B(n_1192),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1250),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1213),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1254),
.B(n_1181),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1250),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1203),
.B(n_1192),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1202),
.B(n_1192),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1202),
.B(n_1198),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1246),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1235),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1227),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1229),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1216),
.B(n_1183),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1230),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1234),
.B(n_1126),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1242),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1252),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1245),
.B(n_1209),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1236),
.B(n_1196),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1236),
.B(n_1195),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1270),
.B(n_1258),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1270),
.B(n_1239),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1272),
.B(n_1239),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1276),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1266),
.B(n_1248),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1272),
.B(n_1240),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1273),
.B(n_1240),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1256),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1257),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1257),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1273),
.B(n_1222),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1259),
.B(n_1219),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1263),
.B(n_1222),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1268),
.B(n_1221),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1269),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1268),
.B(n_1221),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1281),
.B(n_1217),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1271),
.B(n_1220),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1280),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1274),
.B(n_1217),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1260),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1274),
.B(n_1206),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1271),
.B(n_1220),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1262),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1261),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1261),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1264),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1267),
.B(n_1214),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1282),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1314),
.B(n_1277),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1313),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1295),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1295),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1296),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1287),
.B(n_1289),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1314),
.B(n_1277),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1296),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1299),
.B(n_1278),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1315),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1311),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1311),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1299),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1315),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1304),
.B(n_1285),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1287),
.B(n_1279),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1309),
.B(n_1285),
.Y(n_1332)
);

AND2x2_ASAP7_75t_SL g1333 ( 
.A(n_1299),
.B(n_1207),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1288),
.B(n_1283),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1312),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1298),
.B(n_1286),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1325),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1325),
.Y(n_1338)
);

AO32x1_ASAP7_75t_L g1339 ( 
.A1(n_1318),
.A2(n_1225),
.A3(n_1275),
.B1(n_1210),
.B2(n_1301),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1331),
.B(n_1289),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1316),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1329),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1333),
.A2(n_1284),
.B(n_1265),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1333),
.A2(n_1209),
.B1(n_1233),
.B2(n_1291),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1329),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1330),
.B(n_1294),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1319),
.Y(n_1347)
);

AOI21xp33_ASAP7_75t_L g1348 ( 
.A1(n_1336),
.A2(n_1302),
.B(n_1300),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1320),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1323),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1334),
.A2(n_1233),
.B1(n_1275),
.B2(n_1237),
.Y(n_1351)
);

BUFx2_ASAP7_75t_SL g1352 ( 
.A(n_1324),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1326),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1340),
.B(n_1290),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1344),
.A2(n_1330),
.B1(n_1332),
.B2(n_1336),
.C(n_1307),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1347),
.Y(n_1356)
);

CKINVDCx16_ASAP7_75t_R g1357 ( 
.A(n_1343),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1343),
.A2(n_1332),
.B1(n_1310),
.B2(n_1303),
.C(n_1317),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1351),
.A2(n_1324),
.B(n_1328),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1349),
.Y(n_1360)
);

AOI211xp5_ASAP7_75t_L g1361 ( 
.A1(n_1348),
.A2(n_1303),
.B(n_1238),
.C(n_1224),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1357),
.A2(n_1352),
.B1(n_1341),
.B2(n_1328),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1361),
.A2(n_1346),
.B(n_1350),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1356),
.Y(n_1364)
);

OAI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1355),
.A2(n_1345),
.B1(n_1337),
.B2(n_1338),
.C(n_1342),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1360),
.A2(n_1358),
.B(n_1321),
.Y(n_1366)
);

AOI322xp5_ASAP7_75t_L g1367 ( 
.A1(n_1366),
.A2(n_1292),
.A3(n_1297),
.B1(n_1293),
.B2(n_1308),
.C1(n_1306),
.C2(n_1255),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1364),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1363),
.B(n_1322),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1365),
.B(n_1353),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1362),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1364),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1368),
.Y(n_1373)
);

NOR3xp33_ASAP7_75t_L g1374 ( 
.A(n_1371),
.B(n_1359),
.C(n_1224),
.Y(n_1374)
);

NOR3xp33_ASAP7_75t_SL g1375 ( 
.A(n_1372),
.B(n_1238),
.C(n_1305),
.Y(n_1375)
);

NOR3xp33_ASAP7_75t_L g1376 ( 
.A(n_1373),
.B(n_1370),
.C(n_1247),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1375),
.Y(n_1377)
);

XNOR2xp5_ASAP7_75t_L g1378 ( 
.A(n_1377),
.B(n_1374),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1378),
.B(n_1376),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1379),
.Y(n_1380)
);

OAI31xp33_ASAP7_75t_L g1381 ( 
.A1(n_1379),
.A2(n_1369),
.A3(n_1367),
.B(n_1226),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1380),
.A2(n_1354),
.B1(n_1212),
.B2(n_1231),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1381),
.A2(n_1205),
.B(n_1241),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1382),
.A2(n_1205),
.B(n_1218),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1383),
.A2(n_1228),
.B(n_1327),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1384),
.B(n_1204),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1385),
.B(n_1199),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1387),
.A2(n_1339),
.B(n_1335),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1388),
.B(n_1386),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1389),
.A2(n_1215),
.B1(n_1232),
.B2(n_1243),
.Y(n_1390)
);


endmodule