module fake_jpeg_961_n_608 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_608);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_608;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_58),
.Y(n_187)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_59),
.Y(n_138)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_78),
.Y(n_183)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_35),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_86),
.Y(n_147)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_89),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_32),
.Y(n_95)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_123),
.Y(n_154)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_111),
.A2(n_45),
.B(n_2),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_119),
.B(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_55),
.Y(n_128)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_52),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_50),
.Y(n_174)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_46),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_127),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_128),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_41),
.B(n_20),
.C(n_26),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_130),
.B(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_41),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_136),
.B(n_141),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_37),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_37),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_142),
.B(n_155),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_40),
.B1(n_55),
.B2(n_48),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_144),
.A2(n_160),
.B1(n_178),
.B2(n_218),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_80),
.A2(n_96),
.B1(n_97),
.B2(n_92),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_149),
.A2(n_112),
.B1(n_110),
.B2(n_103),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_55),
.B1(n_25),
.B2(n_40),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_150),
.A2(n_157),
.B1(n_197),
.B2(n_200),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_106),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_25),
.B1(n_40),
.B2(n_43),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_158),
.B(n_168),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_58),
.A2(n_76),
.B1(n_48),
.B2(n_54),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_71),
.A2(n_44),
.B1(n_20),
.B2(n_50),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_195),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_104),
.A2(n_48),
.B1(n_44),
.B2(n_46),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_109),
.B(n_49),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_190),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_113),
.B(n_49),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_73),
.A2(n_29),
.B1(n_26),
.B2(n_19),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_101),
.A2(n_53),
.B1(n_52),
.B2(n_29),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_81),
.A2(n_53),
.B1(n_19),
.B2(n_45),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_62),
.B(n_1),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_63),
.B(n_1),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_98),
.B(n_121),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_210),
.B(n_213),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_118),
.B(n_2),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_126),
.B(n_3),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_127),
.B(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_214),
.B(n_217),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_70),
.B(n_5),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_94),
.A2(n_45),
.B1(n_7),
.B2(n_9),
.Y(n_218)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_220),
.Y(n_329)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_221),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_222),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_150),
.A2(n_157),
.B1(n_154),
.B2(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_223),
.A2(n_267),
.B1(n_171),
.B2(n_169),
.Y(n_299)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_224),
.Y(n_328)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_226),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_227),
.A2(n_259),
.B1(n_287),
.B2(n_173),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_129),
.B(n_75),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_228),
.Y(n_335)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_230),
.Y(n_337)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_232),
.Y(n_349)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_137),
.Y(n_235)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_237),
.Y(n_346)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_238),
.Y(n_353)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_148),
.Y(n_240)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_242),
.Y(n_348)
);

AO22x1_ASAP7_75t_SL g244 ( 
.A1(n_135),
.A2(n_102),
.B1(n_117),
.B2(n_116),
.Y(n_244)
);

AO22x1_ASAP7_75t_SL g347 ( 
.A1(n_244),
.A2(n_267),
.B1(n_228),
.B2(n_268),
.Y(n_347)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_246),
.Y(n_326)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_248),
.A2(n_286),
.B1(n_292),
.B2(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_251),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_134),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_252),
.B(n_273),
.Y(n_323)
);

BUFx4f_ASAP7_75t_SL g253 ( 
.A(n_172),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_253),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_254),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_161),
.A2(n_196),
.B1(n_184),
.B2(n_163),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_256),
.A2(n_258),
.B1(n_266),
.B2(n_272),
.Y(n_320)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_161),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_149),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_264),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_265),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_163),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_152),
.A2(n_165),
.B1(n_198),
.B2(n_178),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_199),
.B(n_13),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_147),
.B(n_18),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_269),
.B(n_282),
.Y(n_324)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

AOI222xp33_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_17),
.C2(n_18),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_274),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_160),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_134),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_192),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_164),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_275),
.B(n_277),
.Y(n_345)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_276),
.Y(n_304)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_176),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_167),
.B(n_18),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_14),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_283),
.B(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_166),
.B(n_188),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_193),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_176),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_201),
.A2(n_14),
.B1(n_15),
.B2(n_144),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_289),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_203),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_290),
.B(n_291),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_162),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_172),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_151),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_200),
.B(n_182),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_297),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_206),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_295),
.A2(n_222),
.B1(n_270),
.B2(n_220),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_206),
.A2(n_182),
.B1(n_169),
.B2(n_171),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_133),
.B1(n_140),
.B2(n_146),
.Y(n_310)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_181),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_299),
.A2(n_301),
.B1(n_308),
.B2(n_313),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_300),
.A2(n_254),
.B1(n_271),
.B2(n_232),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_233),
.A2(n_211),
.B1(n_179),
.B2(n_143),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_231),
.A2(n_173),
.B(n_162),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_303),
.A2(n_258),
.B(n_276),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_223),
.A2(n_133),
.B1(n_140),
.B2(n_143),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_305),
.A2(n_253),
.B1(n_255),
.B2(n_278),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_243),
.A2(n_179),
.B1(n_211),
.B2(n_146),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_310),
.A2(n_256),
.B1(n_244),
.B2(n_240),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_249),
.B(n_176),
.C(n_207),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_285),
.C(n_239),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_231),
.A2(n_207),
.B1(n_236),
.B2(n_281),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_233),
.A2(n_207),
.B1(n_250),
.B2(n_248),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_316),
.A2(n_322),
.B1(n_344),
.B2(n_286),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_234),
.B1(n_241),
.B2(n_272),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_339),
.A2(n_253),
.B1(n_221),
.B2(n_230),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_234),
.A2(n_287),
.B1(n_245),
.B2(n_280),
.Y(n_344)
);

AO21x2_ASAP7_75t_L g388 ( 
.A1(n_347),
.A2(n_303),
.B(n_338),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_337),
.Y(n_355)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_228),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_358),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_328),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_325),
.B(n_247),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_361),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_324),
.B(n_226),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_335),
.B(n_257),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_362),
.A2(n_319),
.B(n_349),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_246),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_342),
.C(n_340),
.Y(n_416)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_323),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_366),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_311),
.B(n_274),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_367),
.B(n_369),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_368),
.A2(n_397),
.B1(n_319),
.B2(n_329),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_244),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_377),
.Y(n_429)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_373),
.A2(n_388),
.B1(n_334),
.B2(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_314),
.C(n_333),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_376),
.C(n_346),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_229),
.C(n_289),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_298),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_343),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_378),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_379),
.B(n_381),
.Y(n_408)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_277),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_299),
.A2(n_266),
.B1(n_242),
.B2(n_291),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_326),
.Y(n_385)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_305),
.A2(n_347),
.B1(n_320),
.B2(n_301),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_302),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_393),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_389),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_307),
.Y(n_390)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_314),
.B(n_351),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_391),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_304),
.B(n_302),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_333),
.A2(n_351),
.B1(n_350),
.B2(n_317),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_394),
.A2(n_332),
.B1(n_353),
.B2(n_346),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_315),
.Y(n_395)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_395),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_315),
.B(n_327),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_396),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_336),
.B(n_354),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_398),
.A2(n_399),
.B1(n_336),
.B2(n_349),
.Y(n_421)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_381),
.A2(n_317),
.B1(n_321),
.B2(n_318),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_402),
.A2(n_404),
.B1(n_411),
.B2(n_382),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_388),
.A2(n_321),
.B1(n_342),
.B2(n_341),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_388),
.A2(n_334),
.B(n_341),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_415),
.A2(n_362),
.B(n_387),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_394),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_354),
.C(n_352),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_422),
.C(n_431),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_352),
.C(n_340),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_424),
.A2(n_435),
.B1(n_388),
.B2(n_363),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_436),
.A2(n_462),
.B(n_466),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_437),
.A2(n_441),
.B1(n_463),
.B2(n_464),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_423),
.Y(n_438)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_378),
.Y(n_439)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_439),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_407),
.A2(n_386),
.B1(n_388),
.B2(n_384),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_372),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_444),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_369),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_443),
.B(n_445),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_374),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_361),
.C(n_360),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_429),
.B(n_367),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_446),
.B(n_428),
.Y(n_483)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_448),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_424),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_451),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_377),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_428),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_395),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_455),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_461),
.C(n_467),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_423),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_407),
.A2(n_388),
.B1(n_363),
.B2(n_357),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_456),
.A2(n_458),
.B1(n_468),
.B2(n_409),
.Y(n_479)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_412),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_457),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_408),
.A2(n_370),
.B1(n_393),
.B2(n_396),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_413),
.B(n_358),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_459),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_415),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_460),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_359),
.C(n_376),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_408),
.A2(n_379),
.B(n_380),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_420),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_420),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_426),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_465),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_434),
.A2(n_385),
.B(n_371),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_417),
.C(n_403),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_433),
.A2(n_365),
.B1(n_398),
.B2(n_399),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_467),
.B(n_403),
.Y(n_470)
);

XNOR2x1_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_472),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_450),
.B(n_403),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_431),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_474),
.B(n_499),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_483),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_441),
.A2(n_433),
.B1(n_435),
.B2(n_406),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_478),
.A2(n_485),
.B1(n_455),
.B2(n_438),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_479),
.A2(n_486),
.B1(n_488),
.B2(n_449),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_416),
.C(n_422),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_487),
.C(n_494),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_437),
.A2(n_406),
.B1(n_409),
.B2(n_404),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_443),
.A2(n_410),
.B1(n_426),
.B2(n_434),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_425),
.C(n_430),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_411),
.B1(n_402),
.B2(n_427),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_425),
.C(n_430),
.Y(n_494)
);

XOR2x2_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_421),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_436),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_401),
.C(n_390),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_476),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_439),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_459),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_446),
.B(n_401),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_501),
.A2(n_512),
.B1(n_518),
.B2(n_519),
.Y(n_542)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_490),
.Y(n_503)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_479),
.A2(n_465),
.B1(n_460),
.B2(n_442),
.Y(n_504)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_491),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_505),
.B(n_520),
.Y(n_538)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_506),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_508),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_473),
.B(n_452),
.Y(n_510)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_510),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_509),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_491),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_515),
.Y(n_539)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_493),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_516),
.A2(n_498),
.B(n_471),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_481),
.B(n_444),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g530 ( 
.A(n_517),
.Y(n_530)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_492),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_478),
.A2(n_454),
.B1(n_447),
.B2(n_462),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_521),
.A2(n_525),
.B1(n_498),
.B2(n_488),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_472),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_SL g540 ( 
.A(n_522),
.B(n_475),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_474),
.B(n_466),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_524),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_470),
.B(n_468),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_469),
.A2(n_464),
.B1(n_463),
.B2(n_457),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_SL g526 ( 
.A1(n_504),
.A2(n_482),
.B(n_485),
.C(n_480),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_492),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_523),
.B(n_499),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_527),
.B(n_529),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_475),
.C(n_484),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_540),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_536),
.A2(n_544),
.B1(n_518),
.B2(n_524),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_537),
.B(n_496),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_507),
.B(n_494),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_513),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_501),
.A2(n_482),
.B1(n_489),
.B2(n_477),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_510),
.B1(n_525),
.B2(n_514),
.Y(n_546)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_546),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_537),
.A2(n_521),
.B(n_515),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_548),
.B(n_551),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_549),
.A2(n_556),
.B1(n_558),
.B2(n_541),
.Y(n_567)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_550),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_534),
.B(n_513),
.C(n_511),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_542),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_552),
.B(n_554),
.Y(n_569)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_539),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_561),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_538),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_544),
.A2(n_506),
.B1(n_503),
.B2(n_495),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_557),
.B(n_559),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_536),
.A2(n_533),
.B1(n_532),
.B2(n_539),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_543),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_560),
.B(n_526),
.Y(n_572)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_528),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_555),
.B(n_535),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_563),
.B(n_566),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_560),
.A2(n_532),
.B(n_533),
.Y(n_564)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_564),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_535),
.Y(n_566)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_558),
.A2(n_526),
.B1(n_531),
.B2(n_483),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_568),
.A2(n_570),
.B1(n_572),
.B2(n_574),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_547),
.B(n_432),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_560),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_575),
.B(n_556),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_577),
.B(n_579),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_551),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_557),
.C(n_555),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_582),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_529),
.C(n_527),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_502),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_584),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_509),
.C(n_502),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_573),
.B(n_432),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_586),
.B(n_562),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_580),
.A2(n_569),
.B(n_581),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_587),
.A2(n_588),
.B(n_564),
.Y(n_597)
);

NAND2x1_ASAP7_75t_L g588 ( 
.A(n_578),
.B(n_568),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_576),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_589),
.B(n_592),
.Y(n_596)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_585),
.Y(n_592)
);

INVxp33_ASAP7_75t_L g599 ( 
.A(n_594),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_590),
.B(n_569),
.C(n_581),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_595),
.B(n_582),
.C(n_432),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_597),
.A2(n_598),
.B(n_584),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_591),
.A2(n_572),
.B(n_583),
.Y(n_598)
);

OAI321xp33_ASAP7_75t_L g600 ( 
.A1(n_596),
.A2(n_588),
.A3(n_526),
.B1(n_448),
.B2(n_590),
.C(n_593),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_600),
.A2(n_601),
.B(n_602),
.Y(n_604)
);

AOI321xp33_ASAP7_75t_L g603 ( 
.A1(n_601),
.A2(n_599),
.A3(n_405),
.B1(n_355),
.B2(n_383),
.C(n_332),
.Y(n_603)
);

AO21x1_ASAP7_75t_L g605 ( 
.A1(n_603),
.A2(n_405),
.B(n_400),
.Y(n_605)
);

BUFx24_ASAP7_75t_SL g606 ( 
.A(n_605),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_606),
.A2(n_604),
.B1(n_331),
.B2(n_329),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_331),
.Y(n_608)
);


endmodule