module fake_jpeg_17799_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_0),
.B(n_8),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_42),
.B(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_0),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_52),
.B(n_56),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_55),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_1),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_39),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_68),
.B(n_81),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_33),
.B1(n_28),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_72),
.A2(n_74),
.B1(n_82),
.B2(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_33),
.B1(n_28),
.B2(n_20),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_31),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_33),
.B1(n_31),
.B2(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_87),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_85),
.A2(n_102),
.B1(n_6),
.B2(n_12),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_27),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_35),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_29),
.B1(n_59),
.B2(n_37),
.Y(n_115)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_37),
.B(n_10),
.Y(n_123)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_31),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_24),
.Y(n_105)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_26),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_22),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_112),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_36),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_29),
.B(n_23),
.C(n_22),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_36),
.C(n_21),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_117),
.C(n_76),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_77),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_36),
.C(n_37),
.Y(n_117)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_37),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_138),
.B1(n_86),
.B2(n_80),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_142),
.B(n_137),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_70),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_86),
.B1(n_80),
.B2(n_78),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_5),
.B1(n_13),
.B2(n_12),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_147),
.B1(n_108),
.B2(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_135),
.Y(n_150)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_77),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_76),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_95),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_15),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_2),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_3),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_92),
.B1(n_102),
.B2(n_93),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_104),
.B(n_92),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_164),
.B(n_171),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_156),
.B1(n_178),
.B2(n_134),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_177),
.B1(n_158),
.B2(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_75),
.B1(n_94),
.B2(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_162),
.B(n_172),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_118),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_104),
.B(n_79),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_116),
.B(n_123),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_117),
.C(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_129),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_146),
.B1(n_144),
.B2(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_180),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_118),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_184),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_113),
.A3(n_120),
.B1(n_132),
.B2(n_126),
.C1(n_139),
.C2(n_136),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_136),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_188),
.B1(n_199),
.B2(n_180),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_135),
.B1(n_133),
.B2(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_191),
.Y(n_216)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_109),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_139),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_203),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_167),
.C(n_182),
.Y(n_221)
);

AO22x1_ASAP7_75t_L g198 ( 
.A1(n_157),
.A2(n_164),
.B1(n_158),
.B2(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_160),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_167),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_175),
.Y(n_203)
);

NOR4xp25_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_166),
.C(n_155),
.D(n_149),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_188),
.A3(n_187),
.B1(n_203),
.B2(n_194),
.C1(n_198),
.C2(n_186),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_173),
.B1(n_171),
.B2(n_159),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_197),
.B1(n_185),
.B2(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_178),
.A3(n_152),
.B1(n_149),
.B2(n_162),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_213),
.B(n_215),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_212),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_150),
.B(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_174),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_151),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_221),
.C(n_224),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_223),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_167),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_207),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_209),
.C(n_204),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_230),
.B1(n_215),
.B2(n_216),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_184),
.B1(n_185),
.B2(n_199),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_214),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_222),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_218),
.B(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_193),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_198),
.C(n_190),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_224),
.C(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_247),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_234),
.B(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_217),
.C(n_220),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_211),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_239),
.C(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_250),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_206),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_225),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_253),
.B(n_213),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_257),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_260),
.B(n_263),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_252),
.A3(n_253),
.B1(n_235),
.B2(n_208),
.C1(n_231),
.C2(n_241),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_228),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_226),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_265),
.C(n_259),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_234),
.B(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_268),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_226),
.A3(n_235),
.B1(n_237),
.B2(n_242),
.C1(n_258),
.C2(n_261),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_269),
.B(n_258),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_226),
.C(n_237),
.Y(n_273)
);


endmodule