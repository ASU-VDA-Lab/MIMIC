module fake_jpeg_1801_n_404 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_404);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_404;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_52),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_61),
.Y(n_94)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_25),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_71),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_81),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

NAND2x1_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_39),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_76),
.Y(n_123)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_38),
.B1(n_17),
.B2(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_85),
.A2(n_91),
.B1(n_108),
.B2(n_117),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_86),
.A2(n_90),
.B1(n_112),
.B2(n_4),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_37),
.B1(n_34),
.B2(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_43),
.A2(n_17),
.B1(n_36),
.B2(n_39),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_30),
.B1(n_35),
.B2(n_22),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_97),
.A2(n_76),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_34),
.B1(n_39),
.B2(n_35),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_104),
.A2(n_120),
.B1(n_9),
.B2(n_89),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_45),
.A2(n_39),
.B1(n_34),
.B2(n_16),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_127),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_30),
.B1(n_18),
.B2(n_26),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_68),
.B1(n_62),
.B2(n_54),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_40),
.B1(n_19),
.B2(n_26),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_118),
.A2(n_124),
.B1(n_131),
.B2(n_134),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_26),
.B1(n_40),
.B2(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_132),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_40),
.B1(n_26),
.B2(n_2),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_49),
.A2(n_0),
.B(n_1),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_80),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_0),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_136),
.Y(n_194)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_60),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_142),
.Y(n_195)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_51),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_141),
.B(n_144),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_60),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_51),
.B(n_64),
.C(n_44),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_149),
.Y(n_209)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_77),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_148),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_88),
.B(n_81),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_78),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_151),
.B(n_152),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_14),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_2),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_76),
.C(n_44),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_106),
.C(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_156),
.B(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_3),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_158),
.A2(n_185),
.B1(n_157),
.B2(n_153),
.Y(n_224)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

CKINVDCx12_ASAP7_75t_R g161 ( 
.A(n_87),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_100),
.B(n_12),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_163),
.B(n_169),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_176),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_6),
.C(n_8),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_6),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_167),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_8),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_8),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_8),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_172),
.B(n_181),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_123),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_180),
.Y(n_196)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_89),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_186),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g186 ( 
.A(n_129),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_104),
.B1(n_106),
.B2(n_116),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_192),
.A2(n_216),
.B(n_193),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_137),
.A2(n_109),
.B1(n_114),
.B2(n_116),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_178),
.B1(n_170),
.B2(n_160),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_137),
.A2(n_114),
.B1(n_99),
.B2(n_128),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_224),
.B1(n_167),
.B2(n_182),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_122),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_214),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_92),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_103),
.B(n_120),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_143),
.B(n_130),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_221),
.B(n_154),
.C(n_156),
.D(n_180),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_139),
.B(n_126),
.C(n_103),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.C(n_176),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_9),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_146),
.B(n_105),
.C(n_9),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_173),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_136),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_266),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_155),
.B(n_176),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_240),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_217),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_250),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_243),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_138),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_244),
.C(n_246),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_184),
.B1(n_158),
.B2(n_181),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_238),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_145),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_239),
.B(n_242),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_177),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_147),
.C(n_140),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_175),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_253),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_159),
.B1(n_162),
.B2(n_224),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_215),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_210),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_196),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_216),
.B1(n_218),
.B2(n_202),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_262),
.B1(n_225),
.B2(n_238),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_204),
.A2(n_194),
.B1(n_205),
.B2(n_199),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_258),
.A2(n_188),
.B1(n_225),
.B2(n_187),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_227),
.B(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_264),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_193),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_199),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_198),
.B(n_189),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_269),
.A2(n_279),
.B(n_298),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_205),
.B1(n_200),
.B2(n_211),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_271),
.A2(n_284),
.B1(n_260),
.B2(n_240),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_286),
.Y(n_311)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_189),
.CI(n_194),
.CON(n_279),
.SN(n_279)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_243),
.B(n_201),
.CI(n_226),
.CON(n_282),
.SN(n_282)
);

AOI221xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_289),
.B1(n_240),
.B2(n_248),
.C(n_264),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_201),
.C(n_226),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_291),
.C(n_295),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_235),
.A2(n_200),
.B1(n_187),
.B2(n_188),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_285),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_233),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_246),
.C(n_253),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_230),
.B(n_254),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_236),
.C(n_247),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_249),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_234),
.B(n_257),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_292),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_299),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_251),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_300),
.B(n_304),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_292),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_301),
.Y(n_343)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_307),
.C(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_287),
.B(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_270),
.A2(n_289),
.B1(n_267),
.B2(n_279),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_267),
.B1(n_273),
.B2(n_298),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_278),
.B1(n_291),
.B2(n_282),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_232),
.Y(n_310)
);

AOI221xp5_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_316),
.B1(n_318),
.B2(n_320),
.C(n_321),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_276),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_313),
.A2(n_317),
.B(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_270),
.A2(n_241),
.B1(n_252),
.B2(n_255),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_283),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_273),
.B(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_331),
.C(n_334),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_313),
.B1(n_322),
.B2(n_323),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_277),
.B(n_269),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_345),
.B(n_302),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_278),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_332),
.A2(n_333),
.B1(n_337),
.B2(n_342),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_271),
.B1(n_284),
.B2(n_281),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_281),
.C(n_282),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_294),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_324),
.C(n_332),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_268),
.B1(n_285),
.B2(n_319),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_320),
.C(n_315),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_344),
.C(n_318),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_310),
.B1(n_305),
.B2(n_314),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_311),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_326),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_351),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_325),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_356),
.Y(n_365)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_353),
.B(n_340),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_344),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_352),
.A2(n_354),
.B1(n_357),
.B2(n_362),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_345),
.A2(n_306),
.B(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_339),
.C(n_334),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_329),
.C(n_330),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_343),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_359),
.B(n_360),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_360),
.A2(n_348),
.B1(n_353),
.B2(n_352),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_336),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_370),
.C(n_355),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_362),
.A2(n_336),
.B1(n_333),
.B2(n_337),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_374),
.Y(n_378)
);

AO21x1_ASAP7_75t_L g379 ( 
.A1(n_369),
.A2(n_349),
.B(n_354),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_341),
.B(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_363),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_375),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_358),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_368),
.B(n_367),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_382),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_355),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_377),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_385),
.B(n_386),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_364),
.Y(n_386)
);

INVx11_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_389),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_375),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_391),
.B(n_365),
.C(n_384),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_380),
.B(n_365),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_393),
.A2(n_388),
.B1(n_389),
.B2(n_373),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_387),
.A2(n_386),
.B(n_378),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_396),
.A2(n_394),
.B(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_397),
.B(n_398),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_395),
.A2(n_370),
.B(n_378),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_400),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_401),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_395),
.Y(n_404)
);


endmodule