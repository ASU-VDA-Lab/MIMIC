module fake_jpeg_9257_n_132 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_SL g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_33),
.B(n_13),
.Y(n_49)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_12),
.B1(n_18),
.B2(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_47),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_16),
.B1(n_12),
.B2(n_18),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_52),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_53),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_27),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_37),
.B(n_6),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_50),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_32),
.A3(n_31),
.B1(n_22),
.B2(n_8),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_9),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_32),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_32),
.C(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_10),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_71),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_47),
.B1(n_50),
.B2(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_84),
.B(n_74),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_7),
.C(n_8),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_7),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_67),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_68),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_60),
.C(n_69),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_68),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_97),
.C(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_99),
.B(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_109),
.C(n_89),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_86),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_88),
.B1(n_76),
.B2(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_79),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_101),
.A3(n_103),
.B1(n_102),
.B2(n_106),
.C(n_97),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_110),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_115),
.C(n_85),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_94),
.C(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_125),
.B(n_124),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_129),
.C(n_128),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule