module fake_jpeg_19328_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_6),
.B(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_52),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_50),
.Y(n_129)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx12f_ASAP7_75t_SL g55 ( 
.A(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_87),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_59),
.Y(n_123)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_76),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_13),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_82),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_88),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_38),
.B(n_15),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_13),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_42),
.Y(n_128)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_34),
.B1(n_19),
.B2(n_21),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_19),
.B1(n_22),
.B2(n_36),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_103),
.A2(n_107),
.B1(n_132),
.B2(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_104),
.B(n_112),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_50),
.A2(n_26),
.B1(n_41),
.B2(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_41),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_114),
.B(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_47),
.B(n_37),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_82),
.A2(n_63),
.B1(n_64),
.B2(n_26),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_76),
.B(n_18),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_83),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_42),
.B1(n_18),
.B2(n_23),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_80),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_48),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_144),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_49),
.A2(n_22),
.B1(n_36),
.B2(n_25),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_59),
.B1(n_1),
.B2(n_3),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_53),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_152),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_146),
.B(n_159),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_22),
.B1(n_36),
.B2(n_43),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_147),
.A2(n_169),
.B1(n_176),
.B2(n_143),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_97),
.A2(n_43),
.B1(n_29),
.B2(n_33),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_61),
.B1(n_91),
.B2(n_86),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_150),
.A2(n_164),
.B1(n_180),
.B2(n_182),
.Y(n_216)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_56),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_45),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_175),
.B(n_132),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_113),
.A2(n_33),
.B(n_39),
.C(n_35),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_161),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_79),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_79),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_173),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_29),
.B(n_39),
.C(n_35),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_166),
.Y(n_214)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_97),
.A2(n_13),
.B1(n_12),
.B2(n_89),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_102),
.B(n_45),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_72),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_75),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_174),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_110),
.B(n_70),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_105),
.B(n_66),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_184),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_129),
.B(n_0),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_0),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_189),
.Y(n_207)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_122),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

BUFx24_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_107),
.B(n_134),
.C(n_138),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_200),
.B1(n_201),
.B2(n_180),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_196),
.A2(n_197),
.B(n_204),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_96),
.B(n_138),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_131),
.B1(n_130),
.B2(n_120),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_120),
.B1(n_93),
.B2(n_140),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_116),
.B(n_93),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_109),
.B(n_111),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_205),
.A2(n_10),
.B(n_195),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_109),
.B(n_117),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_145),
.B(n_171),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_141),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_220),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_116),
.B1(n_143),
.B2(n_125),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_190),
.B1(n_166),
.B2(n_165),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_175),
.B1(n_183),
.B2(n_155),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_125),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_148),
.B(n_100),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_175),
.Y(n_238)
);

AO22x2_ASAP7_75t_SL g224 ( 
.A1(n_150),
.A2(n_100),
.B1(n_99),
.B2(n_5),
.Y(n_224)
);

AO21x2_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_182),
.B(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_99),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_151),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_229),
.A2(n_245),
.B1(n_255),
.B2(n_259),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_230),
.A2(n_239),
.B1(n_241),
.B2(n_244),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_156),
.B1(n_158),
.B2(n_161),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_234),
.B1(n_247),
.B2(n_205),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_158),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_207),
.B(n_206),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_163),
.B1(n_152),
.B2(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_238),
.B(n_232),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_189),
.B1(n_157),
.B2(n_154),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_185),
.B1(n_160),
.B2(n_159),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_185),
.B1(n_186),
.B2(n_146),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_248),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_188),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_153),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_251),
.A2(n_257),
.B1(n_226),
.B2(n_227),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_191),
.A2(n_181),
.B1(n_183),
.B2(n_177),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_196),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_195),
.A2(n_3),
.B1(n_10),
.B2(n_213),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_10),
.C(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_260),
.C(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_212),
.B(n_199),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_10),
.C(n_193),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_261),
.A2(n_284),
.B1(n_286),
.B2(n_288),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_262),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_265),
.A2(n_268),
.B1(n_273),
.B2(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_193),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_267),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_212),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_215),
.B1(n_212),
.B2(n_224),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_206),
.B(n_200),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_255),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_279),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_215),
.C(n_220),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_260),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_280),
.B(n_287),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_229),
.A2(n_207),
.B1(n_224),
.B2(n_225),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_198),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_236),
.A2(n_224),
.B1(n_227),
.B2(n_226),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_246),
.B1(n_221),
.B2(n_257),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_240),
.B(n_253),
.C(n_234),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_294),
.A2(n_303),
.B(n_304),
.Y(n_329)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_297),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_302),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_230),
.B(n_248),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_231),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_307),
.A2(n_308),
.B1(n_310),
.B2(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_309),
.A2(n_312),
.B1(n_314),
.B2(n_191),
.Y(n_336)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_230),
.B1(n_241),
.B2(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_315),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_261),
.B1(n_274),
.B2(n_230),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_319),
.B1(n_321),
.B2(n_327),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_274),
.B1(n_230),
.B2(n_285),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_278),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_328),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_239),
.B1(n_280),
.B2(n_253),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_265),
.B(n_254),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_290),
.B(n_292),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_266),
.C(n_279),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_326),
.C(n_313),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_267),
.C(n_277),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_306),
.A2(n_264),
.B1(n_247),
.B2(n_271),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_287),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_300),
.B(n_253),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_194),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_264),
.B(n_271),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g350 ( 
.A(n_332),
.B(n_303),
.C(n_304),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_310),
.A2(n_263),
.B1(n_221),
.B2(n_209),
.Y(n_334)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

NAND2x1_ASAP7_75t_SL g338 ( 
.A(n_317),
.B(n_305),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_338),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_339),
.A2(n_347),
.B1(n_332),
.B2(n_321),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_343),
.C(n_353),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_325),
.B(n_308),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_352),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_303),
.C(n_301),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_295),
.Y(n_345)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_292),
.B1(n_302),
.B2(n_291),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_293),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_348),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_314),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_349),
.Y(n_355)
);

AO21x1_ASAP7_75t_L g359 ( 
.A1(n_350),
.A2(n_329),
.B(n_322),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_326),
.B(n_194),
.Y(n_352)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_356),
.Y(n_378)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_331),
.C(n_320),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_362),
.B(n_365),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_366),
.Y(n_370)
);

AO22x1_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_329),
.B1(n_331),
.B2(n_319),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_327),
.C(n_333),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

AO22x1_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_323),
.B1(n_333),
.B2(n_330),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_369),
.A2(n_344),
.B1(n_346),
.B2(n_339),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_353),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

INVx11_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_376),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_367),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_337),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_340),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_363),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_371),
.B(n_362),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_372),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_359),
.B(n_358),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_382),
.B(n_380),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_386),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_378),
.A2(n_354),
.B1(n_365),
.B2(n_355),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_360),
.C(n_366),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_387),
.B(n_388),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_360),
.C(n_364),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_396),
.C(n_388),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_384),
.B(n_375),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_393),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_389),
.A2(n_370),
.B(n_380),
.Y(n_394)
);

NOR2x1_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_395),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_355),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_397),
.B(n_399),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_381),
.C(n_383),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_374),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_398),
.A2(n_393),
.B(n_383),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_401),
.A2(n_403),
.B(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_364),
.C(n_369),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_406),
.A2(n_405),
.B(n_368),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_369),
.C(n_328),
.Y(n_408)
);

FAx1_ASAP7_75t_SL g409 ( 
.A(n_408),
.B(n_337),
.CI(n_395),
.CON(n_409),
.SN(n_409)
);


endmodule