module real_aes_5584_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_1025, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_1028, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_1027, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_1026, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_1024, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_1025;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_1028;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_1027;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_1026;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_1024;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_287;
wire n_792;
wire n_673;
wire n_357;
wire n_386;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_994;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_976;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_973;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_1013;
wire n_1017;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_363;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_288;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_1003;
wire n_1000;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_0), .A2(n_435), .B(n_438), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_1), .A2(n_140), .B1(n_328), .B2(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g463 ( .A(n_2), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_3), .A2(n_96), .B1(n_420), .B2(n_510), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_4), .A2(n_6), .B1(n_367), .B2(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_5), .Y(n_767) );
AND2x4_ASAP7_75t_L g778 ( .A(n_5), .B(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g784 ( .A(n_5), .B(n_260), .Y(n_784) );
AOI221x1_ASAP7_75t_L g542 ( .A1(n_7), .A2(n_73), .B1(n_437), .B2(n_543), .C(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g715 ( .A(n_8), .Y(n_715) );
AO22x1_ASAP7_75t_L g782 ( .A1(n_9), .A2(n_12), .B1(n_783), .B2(n_785), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_10), .A2(n_165), .B1(n_421), .B2(n_476), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_11), .A2(n_153), .B1(n_369), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_13), .A2(n_196), .B1(n_775), .B2(n_790), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_14), .A2(n_136), .B1(n_364), .B2(n_502), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_15), .A2(n_225), .B1(n_425), .B2(n_426), .Y(n_681) );
INVx1_ASAP7_75t_L g702 ( .A(n_16), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_17), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_18), .A2(n_119), .B1(n_425), .B2(n_652), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_19), .A2(n_127), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_20), .A2(n_81), .B1(n_313), .B2(n_317), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_21), .A2(n_252), .B1(n_441), .B2(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_22), .B(n_545), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_23), .A2(n_82), .B1(n_417), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_24), .A2(n_152), .B1(n_443), .B2(n_445), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_25), .Y(n_560) );
INVx1_ASAP7_75t_L g755 ( .A(n_26), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_27), .B(n_617), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_28), .A2(n_232), .B1(n_277), .B2(n_299), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_29), .A2(n_61), .B1(n_417), .B2(n_482), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_30), .A2(n_104), .B1(n_385), .B2(n_387), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_31), .A2(n_263), .B1(n_652), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g574 ( .A(n_32), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_33), .A2(n_259), .B1(n_415), .B2(n_416), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_34), .A2(n_71), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_35), .A2(n_164), .B1(n_617), .B2(n_669), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_36), .A2(n_160), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g505 ( .A(n_37), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_38), .A2(n_87), .B1(n_367), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_39), .A2(n_264), .B1(n_385), .B2(n_527), .Y(n_750) );
INVx1_ASAP7_75t_L g296 ( .A(n_40), .Y(n_296) );
INVxp67_ASAP7_75t_L g336 ( .A(n_40), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_40), .B(n_202), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_41), .A2(n_44), .B1(n_430), .B2(n_713), .C(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g514 ( .A(n_42), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_43), .A2(n_223), .B1(n_498), .B2(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g466 ( .A(n_45), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_46), .A2(n_49), .B1(n_373), .B2(n_375), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_47), .A2(n_64), .B1(n_369), .B2(n_423), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_48), .A2(n_216), .B1(n_415), .B2(n_416), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_50), .B(n_443), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_51), .B(n_281), .Y(n_291) );
INVx1_ASAP7_75t_L g522 ( .A(n_52), .Y(n_522) );
INVx1_ASAP7_75t_L g454 ( .A(n_53), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_54), .A2(n_170), .B1(n_456), .B2(n_610), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_55), .A2(n_401), .B(n_403), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_56), .A2(n_111), .B1(n_725), .B2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_57), .A2(n_122), .B1(n_373), .B2(n_495), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_58), .A2(n_178), .B1(n_785), .B2(n_801), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_59), .A2(n_262), .B1(n_426), .B2(n_479), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_60), .A2(n_155), .B1(n_415), .B2(n_580), .Y(n_727) );
INVx2_ASAP7_75t_L g765 ( .A(n_62), .Y(n_765) );
INVx1_ASAP7_75t_L g777 ( .A(n_63), .Y(n_777) );
AND2x4_ASAP7_75t_L g781 ( .A(n_63), .B(n_765), .Y(n_781) );
INVx1_ASAP7_75t_SL g789 ( .A(n_63), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_65), .A2(n_187), .B1(n_387), .B2(n_395), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_66), .A2(n_251), .B1(n_381), .B2(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_67), .A2(n_209), .B1(n_510), .B2(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g460 ( .A(n_68), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_69), .A2(n_185), .B1(n_783), .B2(n_802), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_70), .A2(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g641 ( .A(n_72), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_74), .A2(n_207), .B1(n_369), .B2(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_75), .A2(n_109), .B1(n_497), .B2(n_499), .Y(n_496) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_76), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_77), .A2(n_228), .B1(n_420), .B2(n_510), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_78), .A2(n_126), .B1(n_420), .B2(n_479), .Y(n_728) );
INVx1_ASAP7_75t_L g447 ( .A(n_79), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_80), .B(n_338), .Y(n_337) );
XOR2x2_ASAP7_75t_L g606 ( .A(n_83), .B(n_607), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_83), .A2(n_167), .B1(n_775), .B2(n_780), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_84), .A2(n_100), .B1(n_671), .B2(n_673), .Y(n_670) );
AO22x2_ASAP7_75t_L g501 ( .A1(n_85), .A2(n_174), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx1_ASAP7_75t_SL g541 ( .A(n_86), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_86), .B(n_569), .C(n_570), .Y(n_568) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_88), .B(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_89), .A2(n_195), .B1(n_785), .B2(n_801), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_90), .A2(n_180), .B1(n_783), .B2(n_785), .Y(n_810) );
INVx1_ASAP7_75t_L g282 ( .A(n_91), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_91), .B(n_200), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_92), .A2(n_231), .B1(n_527), .B2(n_528), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_93), .A2(n_242), .B1(n_598), .B2(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g457 ( .A(n_94), .Y(n_457) );
AOI33xp33_ASAP7_75t_R g625 ( .A1(n_95), .A2(n_230), .A3(n_278), .B1(n_318), .B2(n_626), .B3(n_1026), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_97), .A2(n_189), .B1(n_362), .B2(n_364), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_98), .A2(n_240), .B1(n_362), .B2(n_622), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_99), .Y(n_562) );
INVx1_ASAP7_75t_L g710 ( .A(n_101), .Y(n_710) );
OAI222xp33_ASAP7_75t_L g721 ( .A1(n_101), .A2(n_722), .B1(n_727), .B2(n_728), .C1(n_1027), .C2(n_1028), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_101), .B(n_728), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_102), .A2(n_172), .B1(n_775), .B2(n_798), .Y(n_797) );
AOI222xp33_ASAP7_75t_L g992 ( .A1(n_102), .A2(n_993), .B1(n_1009), .B2(n_1013), .C1(n_1017), .C2(n_1019), .Y(n_992) );
XOR2xp5_ASAP7_75t_L g993 ( .A(n_102), .B(n_994), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_103), .A2(n_212), .B1(n_381), .B2(n_476), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_105), .A2(n_255), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_106), .A2(n_121), .B1(n_775), .B2(n_790), .Y(n_811) );
INVx1_ASAP7_75t_L g358 ( .A(n_107), .Y(n_358) );
INVx1_ASAP7_75t_L g589 ( .A(n_108), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_110), .A2(n_341), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g346 ( .A(n_112), .Y(n_346) );
INVx1_ASAP7_75t_L g644 ( .A(n_113), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_114), .A2(n_344), .B(n_345), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_115), .A2(n_142), .B1(n_314), .B2(n_325), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_116), .A2(n_257), .B1(n_313), .B2(n_314), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_117), .A2(n_213), .B1(n_364), .B2(n_415), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_118), .A2(n_149), .B1(n_367), .B2(n_369), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_120), .A2(n_239), .B1(n_479), .B2(n_652), .Y(n_651) );
AOI22x1_ASAP7_75t_L g629 ( .A1(n_123), .A2(n_630), .B1(n_631), .B2(n_653), .Y(n_629) );
INVx1_ASAP7_75t_L g653 ( .A(n_123), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_123), .A2(n_139), .B1(n_798), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_124), .A2(n_233), .B1(n_369), .B2(n_423), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_125), .A2(n_204), .B1(n_395), .B2(n_397), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_128), .A2(n_184), .B1(n_445), .B2(n_543), .Y(n_1001) );
AO22x1_ASAP7_75t_L g720 ( .A1(n_129), .A2(n_131), .B1(n_423), .B2(n_426), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_130), .A2(n_186), .B1(n_317), .B2(n_325), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_132), .A2(n_138), .B1(n_415), .B2(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_133), .A2(n_249), .B1(n_775), .B2(n_790), .Y(n_817) );
CKINVDCx16_ASAP7_75t_R g703 ( .A(n_134), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_135), .A2(n_151), .B1(n_303), .B2(n_309), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_137), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_141), .A2(n_156), .B1(n_430), .B2(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_143), .A2(n_250), .B1(n_415), .B2(n_580), .Y(n_1007) );
INVx1_ASAP7_75t_L g516 ( .A(n_144), .Y(n_516) );
INVx1_ASAP7_75t_L g439 ( .A(n_145), .Y(n_439) );
INVx1_ASAP7_75t_L g511 ( .A(n_146), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_147), .A2(n_635), .B(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_148), .A2(n_220), .B1(n_385), .B2(n_598), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_150), .A2(n_163), .B1(n_478), .B2(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_154), .A2(n_246), .B1(n_788), .B2(n_790), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_157), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_158), .A2(n_198), .B1(n_379), .B2(n_381), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_159), .A2(n_241), .B1(n_445), .B2(n_617), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_161), .A2(n_169), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_162), .A2(n_215), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_166), .A2(n_430), .B(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_168), .A2(n_218), .B1(n_369), .B2(n_423), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_171), .A2(n_214), .B1(n_793), .B2(n_801), .Y(n_822) );
AOI22x1_ASAP7_75t_L g658 ( .A1(n_173), .A2(n_659), .B1(n_660), .B2(n_682), .Y(n_658) );
INVx1_ASAP7_75t_L g682 ( .A(n_173), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_173), .A2(n_659), .B1(n_660), .B2(n_682), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_175), .A2(n_203), .B1(n_385), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g665 ( .A(n_176), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_177), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_179), .B(n_441), .Y(n_440) );
AO221x2_ASAP7_75t_L g774 ( .A1(n_181), .A2(n_227), .B1(n_775), .B2(n_780), .C(n_782), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_182), .A2(n_266), .B1(n_425), .B2(n_426), .Y(n_424) );
OA22x2_ASAP7_75t_L g286 ( .A1(n_183), .A2(n_202), .B1(n_281), .B2(n_285), .Y(n_286) );
INVx1_ASAP7_75t_L g322 ( .A(n_183), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_188), .A2(n_254), .B1(n_801), .B2(n_802), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_190), .Y(n_555) );
AO22x2_ASAP7_75t_L g448 ( .A1(n_191), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_191), .Y(n_449) );
AND2x2_ASAP7_75t_L g544 ( .A(n_192), .B(n_545), .Y(n_544) );
NAND2xp33_ASAP7_75t_L g696 ( .A(n_193), .B(n_635), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_194), .A2(n_247), .B1(n_421), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_197), .A2(n_211), .B1(n_420), .B2(n_510), .Y(n_578) );
INVx1_ASAP7_75t_L g591 ( .A(n_199), .Y(n_591) );
INVx1_ASAP7_75t_L g298 ( .A(n_200), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_200), .B(n_320), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_201), .A2(n_226), .B1(n_341), .B2(n_342), .Y(n_340) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_202), .A2(n_221), .B(n_324), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_205), .A2(n_219), .B1(n_367), .B2(n_369), .Y(n_648) );
XNOR2x2_ASAP7_75t_SL g273 ( .A(n_206), .B(n_274), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_208), .A2(n_236), .B1(n_277), .B2(n_367), .Y(n_540) );
INVx1_ASAP7_75t_L g740 ( .A(n_210), .Y(n_740) );
INVx1_ASAP7_75t_L g584 ( .A(n_217), .Y(n_584) );
INVx1_ASAP7_75t_L g284 ( .A(n_221), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_221), .B(n_253), .Y(n_352) );
INVx1_ASAP7_75t_L g585 ( .A(n_222), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_224), .A2(n_245), .B1(n_476), .B2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g594 ( .A(n_229), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_234), .A2(n_248), .B1(n_362), .B2(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g642 ( .A(n_235), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_237), .B(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g637 ( .A(n_238), .Y(n_637) );
INVx1_ASAP7_75t_L g404 ( .A(n_243), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_244), .A2(n_258), .B1(n_430), .B2(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_253), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g519 ( .A(n_256), .Y(n_519) );
INVx1_ASAP7_75t_L g779 ( .A(n_260), .Y(n_779) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_260), .Y(n_1021) );
INVx1_ASAP7_75t_L g520 ( .A(n_261), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_265), .A2(n_1014), .B1(n_1015), .B2(n_1016), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_265), .Y(n_1014) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_759), .B(n_768), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_531), .Y(n_268) );
INVx1_ASAP7_75t_L g760 ( .A(n_269), .Y(n_760) );
AO22x1_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_271), .B1(n_409), .B2(n_530), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_355), .B1(n_407), .B2(n_408), .Y(n_271) );
INVx2_ASAP7_75t_L g407 ( .A(n_272), .Y(n_407) );
BUFx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_326), .Y(n_274) );
NAND4xp25_ASAP7_75t_L g275 ( .A(n_276), .B(n_302), .C(n_312), .D(n_316), .Y(n_275) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_287), .Y(n_277) );
AND2x4_ASAP7_75t_L g299 ( .A(n_278), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g328 ( .A(n_278), .B(n_307), .Y(n_328) );
AND2x2_ASAP7_75t_L g341 ( .A(n_278), .B(n_310), .Y(n_341) );
AND2x4_ASAP7_75t_L g368 ( .A(n_278), .B(n_315), .Y(n_368) );
AND2x2_ASAP7_75t_L g374 ( .A(n_278), .B(n_287), .Y(n_374) );
AND2x2_ASAP7_75t_L g386 ( .A(n_278), .B(n_307), .Y(n_386) );
AND2x2_ASAP7_75t_L g392 ( .A(n_278), .B(n_310), .Y(n_392) );
AND2x2_ASAP7_75t_L g427 ( .A(n_278), .B(n_287), .Y(n_427) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_286), .Y(n_278) );
INVx1_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
NAND2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g285 ( .A(n_281), .Y(n_285) );
INVx3_ASAP7_75t_L g290 ( .A(n_281), .Y(n_290) );
NAND2xp33_ASAP7_75t_L g297 ( .A(n_281), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_282), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_284), .A2(n_324), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g306 ( .A(n_286), .Y(n_306) );
AND2x2_ASAP7_75t_L g334 ( .A(n_286), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g339 ( .A(n_286), .B(n_305), .Y(n_339) );
AND2x4_ASAP7_75t_L g313 ( .A(n_287), .B(n_304), .Y(n_313) );
AND2x4_ASAP7_75t_L g317 ( .A(n_287), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g377 ( .A(n_287), .B(n_318), .Y(n_377) );
AND2x4_ASAP7_75t_L g380 ( .A(n_287), .B(n_304), .Y(n_380) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_287), .Y(n_626) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .Y(n_287) );
OR2x2_ASAP7_75t_L g301 ( .A(n_288), .B(n_293), .Y(n_301) );
AND2x4_ASAP7_75t_L g307 ( .A(n_288), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_288), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_290), .B(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_291), .B(n_319), .C(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x4_ASAP7_75t_L g325 ( .A(n_300), .B(n_318), .Y(n_325) );
AND2x4_ASAP7_75t_L g370 ( .A(n_300), .B(n_318), .Y(n_370) );
AND2x4_ASAP7_75t_L g382 ( .A(n_300), .B(n_304), .Y(n_382) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g315 ( .A(n_301), .Y(n_315) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
AND2x4_ASAP7_75t_L g309 ( .A(n_304), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g314 ( .A(n_304), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g363 ( .A(n_304), .B(n_307), .Y(n_363) );
AND2x2_ASAP7_75t_L g365 ( .A(n_304), .B(n_310), .Y(n_365) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x4_ASAP7_75t_L g344 ( .A(n_307), .B(n_339), .Y(n_344) );
AND2x4_ASAP7_75t_L g396 ( .A(n_307), .B(n_339), .Y(n_396) );
AND2x4_ASAP7_75t_L g310 ( .A(n_308), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g338 ( .A(n_310), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g342 ( .A(n_310), .B(n_318), .Y(n_342) );
AND2x4_ASAP7_75t_L g388 ( .A(n_310), .B(n_318), .Y(n_388) );
AND2x4_ASAP7_75t_L g402 ( .A(n_310), .B(n_339), .Y(n_402) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND4xp25_ASAP7_75t_L g326 ( .A(n_327), .B(n_337), .C(n_340), .D(n_343), .Y(n_326) );
INVx2_ASAP7_75t_L g563 ( .A(n_328), .Y(n_563) );
INVx4_ASAP7_75t_L g556 ( .A(n_329), .Y(n_556) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_334), .Y(n_329) );
AND2x4_ASAP7_75t_L g399 ( .A(n_330), .B(n_334), .Y(n_399) );
AND2x2_ASAP7_75t_L g470 ( .A(n_330), .B(n_334), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g349 ( .A(n_332), .Y(n_349) );
INVx2_ASAP7_75t_L g558 ( .A(n_342), .Y(n_558) );
INVx2_ASAP7_75t_L g561 ( .A(n_344), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx2_ASAP7_75t_L g441 ( .A(n_347), .Y(n_441) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_347), .Y(n_472) );
INVx2_ASAP7_75t_SL g599 ( .A(n_347), .Y(n_599) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_347), .Y(n_756) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g406 ( .A(n_348), .Y(n_406) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B(n_353), .Y(n_348) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_350), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
XNOR2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NOR4xp75_ASAP7_75t_L g359 ( .A(n_360), .B(n_371), .C(n_383), .D(n_393), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_366), .Y(n_360) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_363), .Y(n_415) );
INVx3_ASAP7_75t_L g483 ( .A(n_363), .Y(n_483) );
BUFx2_ASAP7_75t_SL g503 ( .A(n_364), .Y(n_503) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
BUFx5_ASAP7_75t_L g580 ( .A(n_365), .Y(n_580) );
BUFx3_ASAP7_75t_L g622 ( .A(n_365), .Y(n_622) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_368), .Y(n_423) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_368), .Y(n_498) );
BUFx12f_ASAP7_75t_L g692 ( .A(n_368), .Y(n_692) );
BUFx3_ASAP7_75t_L g499 ( .A(n_369), .Y(n_499) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx6_ASAP7_75t_L g486 ( .A(n_370), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_378), .Y(n_371) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx4f_ASAP7_75t_L g478 ( .A(n_374), .Y(n_478) );
BUFx2_ASAP7_75t_L g495 ( .A(n_375), .Y(n_495) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx4_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
INVx4_ASAP7_75t_L g479 ( .A(n_376), .Y(n_479) );
INVx2_ASAP7_75t_L g694 ( .A(n_376), .Y(n_694) );
INVx2_ASAP7_75t_SL g746 ( .A(n_376), .Y(n_746) );
INVx8_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
BUFx12f_ASAP7_75t_L g476 ( .A(n_380), .Y(n_476) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_382), .Y(n_510) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_382), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_389), .Y(n_383) );
INVx3_ASAP7_75t_L g458 ( .A(n_385), .Y(n_458) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g433 ( .A(n_386), .Y(n_433) );
BUFx3_ASAP7_75t_L g724 ( .A(n_386), .Y(n_724) );
INVx3_ASAP7_75t_L g464 ( .A(n_387), .Y(n_464) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g446 ( .A(n_388), .Y(n_446) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_388), .Y(n_669) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g437 ( .A(n_391), .Y(n_437) );
INVx2_ASAP7_75t_L g596 ( .A(n_391), .Y(n_596) );
INVx3_ASAP7_75t_SL g635 ( .A(n_391), .Y(n_635) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx3_ASAP7_75t_L g468 ( .A(n_392), .Y(n_468) );
INVx2_ASAP7_75t_L g615 ( .A(n_392), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_400), .Y(n_393) );
INVx2_ASAP7_75t_L g672 ( .A(n_395), .Y(n_672) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_396), .Y(n_430) );
BUFx3_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
INVx4_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_398), .A2(n_439), .B(n_440), .Y(n_438) );
INVx2_ASAP7_75t_L g598 ( .A(n_398), .Y(n_598) );
INVx3_ASAP7_75t_L g646 ( .A(n_398), .Y(n_646) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_398), .A2(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_L g725 ( .A(n_398), .Y(n_725) );
INVx5_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx4f_ASAP7_75t_L g527 ( .A(n_399), .Y(n_527) );
BUFx2_ASAP7_75t_L g612 ( .A(n_399), .Y(n_612) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
BUFx8_ASAP7_75t_SL g543 ( .A(n_402), .Y(n_543) );
INVx2_ASAP7_75t_L g590 ( .A(n_402), .Y(n_590) );
BUFx3_ASAP7_75t_L g617 ( .A(n_402), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx4_ASAP7_75t_L g528 ( .A(n_405), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_405), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g1003 ( .A(n_405), .Y(n_1003) );
INVx4_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g546 ( .A(n_406), .Y(n_546) );
INVx2_ASAP7_75t_L g530 ( .A(n_409), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_489), .B1(n_490), .B2(n_529), .Y(n_409) );
INVx1_ASAP7_75t_L g529 ( .A(n_410), .Y(n_529) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_448), .B1(n_487), .B2(n_488), .Y(n_410) );
INVx1_ASAP7_75t_L g487 ( .A(n_411), .Y(n_487) );
XOR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_447), .Y(n_411) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_428), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_419), .C(n_422), .D(n_424), .Y(n_413) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx8_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_427), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_434), .C(n_442), .Y(n_428) );
INVx4_ASAP7_75t_L g515 ( .A(n_430), .Y(n_515) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_432), .Y(n_517) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_432), .A2(n_644), .B(n_645), .Y(n_643) );
INVx2_ASAP7_75t_L g1000 ( .A(n_432), .Y(n_1000) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g587 ( .A(n_433), .Y(n_587) );
INVx2_ASAP7_75t_L g675 ( .A(n_433), .Y(n_675) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g638 ( .A(n_441), .Y(n_638) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g668 ( .A(n_444), .Y(n_668) );
INVx1_ASAP7_75t_L g592 ( .A(n_445), .Y(n_592) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_446), .A2(n_461), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g610 ( .A(n_446), .Y(n_610) );
INVx2_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_473), .Y(n_451) );
NOR3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_459), .C(n_465), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B1(n_457), .B2(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_463), .B2(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_469), .Y(n_465) );
INVx2_ASAP7_75t_L g713 ( .A(n_467), .Y(n_713) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g525 ( .A(n_468), .Y(n_525) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_480), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_476), .Y(n_507) );
BUFx12f_ASAP7_75t_L g678 ( .A(n_476), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_484), .Y(n_480) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g502 ( .A(n_483), .Y(n_502) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx5_ASAP7_75t_L g620 ( .A(n_486), .Y(n_620) );
INVx1_ASAP7_75t_L g719 ( .A(n_486), .Y(n_719) );
INVx2_ASAP7_75t_L g744 ( .A(n_486), .Y(n_744) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .C(n_512), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
OAI22x1_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_506), .B1(n_508), .B2(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR3xp33_ASAP7_75t_SL g512 ( .A(n_513), .B(n_518), .C(n_521), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_515), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_515), .A2(n_592), .B1(n_641), .B2(n_642), .Y(n_640) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_526), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_532), .A2(n_760), .B(n_761), .Y(n_759) );
XNOR2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_655), .Y(n_532) );
XNOR2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_602), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_571), .B1(n_600), .B2(n_601), .Y(n_534) );
INVx1_ASAP7_75t_L g600 ( .A(n_535), .Y(n_600) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2x1_ASAP7_75t_L g537 ( .A(n_538), .B(n_564), .Y(n_537) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .C(n_551), .Y(n_538) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_542), .B2(n_1024), .Y(n_539) );
INVx1_ASAP7_75t_L g569 ( .A(n_540), .Y(n_569) );
NOR2xp67_ASAP7_75t_L g547 ( .A(n_541), .B(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_541), .A2(n_552), .B1(n_553), .B2(n_1025), .Y(n_551) );
INVx1_ASAP7_75t_L g566 ( .A(n_542), .Y(n_566) );
INVx4_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_548), .B(n_565), .C(n_568), .Y(n_564) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g570 ( .A(n_552), .Y(n_570) );
INVx1_ASAP7_75t_L g567 ( .A(n_553), .Y(n_567) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVxp67_ASAP7_75t_L g601 ( .A(n_571), .Y(n_601) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
XNOR2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_582), .Y(n_575) );
AND4x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .C(n_579), .D(n_581), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_588), .C(n_593), .Y(n_582) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_591), .B2(n_592), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_597), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_627), .B(n_654), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_606), .B(n_629), .Y(n_654) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_618), .Y(n_607) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .C(n_613), .D(n_616), .Y(n_608) );
BUFx3_ASAP7_75t_L g663 ( .A(n_614), .Y(n_663) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g998 ( .A(n_615), .Y(n_998) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .C(n_623), .D(n_625), .Y(n_618) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_647), .Y(n_631) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_640), .C(n_643), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_634), .B(n_639), .Y(n_633) );
NOR2xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_638), .B(n_702), .Y(n_701) );
AND4x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .C(n_650), .D(n_651), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_706), .B2(n_758), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_683), .B1(n_704), .B2(n_705), .Y(n_657) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_676), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_667), .C(n_670), .Y(n_661) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND4xp25_ASAP7_75t_SL g676 ( .A(n_677), .B(n_679), .C(n_680), .D(n_681), .Y(n_676) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g705 ( .A(n_684), .Y(n_705) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XNOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_703), .Y(n_685) );
NAND4xp75_ASAP7_75t_L g686 ( .A(n_687), .B(n_690), .C(n_695), .D(n_698), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_SL g758 ( .A(n_706), .Y(n_758) );
OA22x2_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_736), .B2(n_757), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_709), .B(n_729), .Y(n_708) );
AOI21x1_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_721), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_716), .Y(n_711) );
BUFx2_ASAP7_75t_L g730 ( .A(n_712), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVxp67_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g734 ( .A(n_718), .B(n_727), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_720), .Y(n_735) );
INVx1_ASAP7_75t_L g733 ( .A(n_722), .Y(n_733) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .Y(n_722) );
NAND4xp75_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .C(n_734), .D(n_735), .Y(n_729) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g757 ( .A(n_736), .Y(n_757) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
XNOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_749), .Y(n_741) );
NAND4xp25_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .C(n_747), .D(n_748), .Y(n_742) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .C(n_752), .D(n_753), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
BUFx4_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .C(n_767), .Y(n_762) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_763), .B(n_1011), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_763), .B(n_1012), .Y(n_1018) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_763), .A2(n_767), .B(n_789), .Y(n_1022) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AO21x1_ASAP7_75t_L g1020 ( .A1(n_764), .A2(n_1021), .B(n_1022), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g776 ( .A(n_765), .B(n_777), .Y(n_776) );
AND3x4_ASAP7_75t_L g788 ( .A(n_765), .B(n_778), .C(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_766), .B(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_767), .Y(n_1012) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_990), .B(n_992), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_917), .C(n_955), .Y(n_769) );
OAI221xp5_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_875), .B1(n_876), .B2(n_881), .C(n_901), .Y(n_770) );
NOR4xp25_ASAP7_75t_L g771 ( .A(n_772), .B(n_846), .C(n_860), .D(n_868), .Y(n_771) );
OAI211xp5_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_794), .B(n_812), .C(n_839), .Y(n_772) );
INVx1_ASAP7_75t_L g844 ( .A(n_773), .Y(n_844) );
NOR2x1_ASAP7_75t_L g943 ( .A(n_773), .B(n_849), .Y(n_943) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_786), .Y(n_773) );
INVx1_ASAP7_75t_L g830 ( .A(n_774), .Y(n_830) );
AND2x2_ASAP7_75t_L g859 ( .A(n_774), .B(n_823), .Y(n_859) );
AND2x2_ASAP7_75t_L g865 ( .A(n_774), .B(n_786), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_774), .B(n_820), .Y(n_953) );
OAI321xp33_ASAP7_75t_L g974 ( .A1(n_774), .A2(n_857), .A3(n_949), .B1(n_975), .B2(n_976), .C(n_978), .Y(n_974) );
AND2x2_ASAP7_75t_L g988 ( .A(n_774), .B(n_819), .Y(n_988) );
INVx3_ASAP7_75t_L g879 ( .A(n_775), .Y(n_879) );
AND2x4_ASAP7_75t_L g775 ( .A(n_776), .B(n_778), .Y(n_775) );
AND2x4_ASAP7_75t_L g783 ( .A(n_776), .B(n_784), .Y(n_783) );
AND2x2_ASAP7_75t_L g792 ( .A(n_776), .B(n_784), .Y(n_792) );
AND2x2_ASAP7_75t_L g801 ( .A(n_776), .B(n_784), .Y(n_801) );
AND2x4_ASAP7_75t_L g780 ( .A(n_778), .B(n_781), .Y(n_780) );
AND2x4_ASAP7_75t_L g790 ( .A(n_778), .B(n_781), .Y(n_790) );
AND2x2_ASAP7_75t_L g785 ( .A(n_781), .B(n_784), .Y(n_785) );
AND2x2_ASAP7_75t_L g793 ( .A(n_781), .B(n_784), .Y(n_793) );
AND2x4_ASAP7_75t_L g802 ( .A(n_781), .B(n_784), .Y(n_802) );
INVx1_ASAP7_75t_L g823 ( .A(n_786), .Y(n_823) );
AND2x2_ASAP7_75t_L g835 ( .A(n_786), .B(n_820), .Y(n_835) );
AND2x2_ASAP7_75t_L g854 ( .A(n_786), .B(n_830), .Y(n_854) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_791), .Y(n_786) );
INVx2_ASAP7_75t_SL g799 ( .A(n_790), .Y(n_799) );
INVx1_ASAP7_75t_L g971 ( .A(n_794), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_803), .Y(n_794) );
AND2x2_ASAP7_75t_L g831 ( .A(n_795), .B(n_808), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_795), .B(n_833), .Y(n_855) );
AND2x2_ASAP7_75t_L g867 ( .A(n_795), .B(n_857), .Y(n_867) );
OR2x2_ASAP7_75t_L g893 ( .A(n_795), .B(n_894), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_795), .B(n_815), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_795), .B(n_875), .Y(n_969) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_795), .B(n_874), .Y(n_985) );
INVx4_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g884 ( .A(n_796), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g890 ( .A(n_796), .B(n_809), .Y(n_890) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_796), .B(n_854), .C(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g907 ( .A(n_796), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_796), .B(n_876), .Y(n_929) );
AND2x2_ASAP7_75t_L g932 ( .A(n_796), .B(n_857), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_796), .B(n_886), .Y(n_977) );
NOR3xp33_ASAP7_75t_SL g979 ( .A(n_796), .B(n_910), .C(n_946), .Y(n_979) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_800), .Y(n_796) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OAI332xp33_ASAP7_75t_L g944 ( .A1(n_804), .A2(n_889), .A3(n_945), .B1(n_948), .B2(n_949), .B3(n_950), .C1(n_951), .C2(n_954), .Y(n_944) );
OAI222xp33_ASAP7_75t_SL g961 ( .A1(n_804), .A2(n_819), .B1(n_874), .B2(n_962), .C1(n_966), .C2(n_967), .Y(n_961) );
OR2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
INVx4_ASAP7_75t_L g828 ( .A(n_805), .Y(n_828) );
OR2x2_ASAP7_75t_L g874 ( .A(n_805), .B(n_809), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_805), .B(n_838), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_805), .B(n_815), .Y(n_896) );
AND2x2_ASAP7_75t_L g899 ( .A(n_805), .B(n_808), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_805), .B(n_838), .Y(n_910) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx2_ASAP7_75t_L g833 ( .A(n_808), .Y(n_833) );
OR2x2_ASAP7_75t_L g886 ( .A(n_808), .B(n_828), .Y(n_886) );
INVxp67_ASAP7_75t_L g894 ( .A(n_808), .Y(n_894) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
O2A1O1Ixp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_824), .B(n_831), .C(n_832), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_818), .Y(n_813) );
AND2x2_ASAP7_75t_L g862 ( .A(n_814), .B(n_858), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_814), .B(n_923), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_814), .B(n_853), .Y(n_936) );
AND2x2_ASAP7_75t_L g989 ( .A(n_814), .B(n_885), .Y(n_989) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g838 ( .A(n_815), .Y(n_838) );
AND2x2_ASAP7_75t_L g845 ( .A(n_815), .B(n_819), .Y(n_845) );
INVx3_ASAP7_75t_L g850 ( .A(n_815), .Y(n_850) );
AOI211xp5_ASAP7_75t_L g881 ( .A1(n_815), .A2(n_882), .B(n_887), .C(n_897), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_815), .B(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_815), .B(n_899), .Y(n_966) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx1_ASAP7_75t_L g923 ( .A(n_818), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_823), .Y(n_818) );
AND2x2_ASAP7_75t_L g852 ( .A(n_819), .B(n_844), .Y(n_852) );
AND2x2_ASAP7_75t_L g864 ( .A(n_819), .B(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_819), .B(n_854), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_819), .B(n_905), .Y(n_904) );
AND2x2_ASAP7_75t_L g911 ( .A(n_819), .B(n_859), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_819), .B(n_943), .Y(n_942) );
CKINVDCx6p67_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_820), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g853 ( .A(n_820), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g858 ( .A(n_820), .B(n_859), .Y(n_858) );
AND2x2_ASAP7_75t_L g873 ( .A(n_820), .B(n_844), .Y(n_873) );
AND2x2_ASAP7_75t_L g915 ( .A(n_820), .B(n_849), .Y(n_915) );
AND2x2_ASAP7_75t_L g959 ( .A(n_820), .B(n_905), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_820), .B(n_823), .Y(n_965) );
AND2x2_ASAP7_75t_L g972 ( .A(n_820), .B(n_823), .Y(n_972) );
AND2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_823), .B(n_892), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_829), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_825), .B(n_914), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g956 ( .A1(n_825), .A2(n_957), .B1(n_959), .B2(n_960), .C(n_961), .Y(n_956) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_826), .Y(n_960) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g837 ( .A(n_827), .Y(n_837) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g857 ( .A(n_828), .Y(n_857) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_830), .A2(n_848), .B1(n_919), .B2(n_921), .C(n_924), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_831), .A2(n_938), .B1(n_939), .B2(n_941), .C(n_944), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_831), .B(n_935), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx3_ASAP7_75t_SL g848 ( .A(n_833), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_833), .B(n_875), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_833), .B(n_876), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g950 ( .A(n_835), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g842 ( .A(n_837), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_838), .B(n_964), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_840), .B(n_942), .Y(n_941) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g935 ( .A(n_842), .Y(n_935) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
AND2x2_ASAP7_75t_L g914 ( .A(n_844), .B(n_915), .Y(n_914) );
INVxp67_ASAP7_75t_L g948 ( .A(n_845), .Y(n_948) );
OAI22xp33_ASAP7_75t_SL g846 ( .A1(n_847), .A2(n_851), .B1(n_855), .B2(n_856), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_848), .A2(n_971), .B1(n_972), .B2(n_973), .C(n_974), .Y(n_970) );
NOR2x1_ASAP7_75t_L g870 ( .A(n_849), .B(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_849), .B(n_920), .Y(n_919) );
AND2x2_ASAP7_75t_L g938 ( .A(n_849), .B(n_900), .Y(n_938) );
INVx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AND2x2_ASAP7_75t_L g905 ( .A(n_850), .B(n_865), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g986 ( .A(n_852), .Y(n_986) );
INVx1_ASAP7_75t_L g888 ( .A(n_853), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g987 ( .A1(n_853), .A2(n_988), .B(n_989), .Y(n_987) );
INVx1_ASAP7_75t_L g946 ( .A(n_854), .Y(n_946) );
INVx1_ASAP7_75t_L g902 ( .A(n_855), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_L g912 ( .A1(n_857), .A2(n_863), .B(n_913), .C(n_916), .Y(n_912) );
INVx1_ASAP7_75t_L g967 ( .A(n_858), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_859), .B(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_859), .B(n_915), .Y(n_927) );
INVx1_ASAP7_75t_L g947 ( .A(n_859), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_863), .B(n_866), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_865), .B(n_915), .Y(n_958) );
INVx1_ASAP7_75t_L g975 ( .A(n_865), .Y(n_975) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
AOI21xp33_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_872), .B(n_874), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g900 ( .A(n_871), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_872), .B(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_876), .Y(n_875) );
OAI221xp5_ASAP7_75t_SL g917 ( .A1(n_876), .A2(n_918), .B1(n_928), .B2(n_930), .C(n_937), .Y(n_917) );
OAI221xp5_ASAP7_75t_SL g955 ( .A1(n_876), .A2(n_956), .B1(n_968), .B2(n_970), .C(n_980), .Y(n_955) );
AND2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_880), .Y(n_876) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_878), .Y(n_991) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVxp67_ASAP7_75t_SL g882 ( .A(n_883), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_884), .A2(n_921), .B1(n_981), .B2(n_982), .C(n_983), .Y(n_980) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_891), .B2(n_893), .C(n_895), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
INVx1_ASAP7_75t_L g920 ( .A(n_899), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_899), .B(n_926), .Y(n_925) );
AOI211xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B(n_906), .C(n_912), .Y(n_901) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_903), .A2(n_931), .B(n_933), .Y(n_930) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_911), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_916), .Y(n_982) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVxp67_ASAP7_75t_SL g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_936), .Y(n_933) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g981 ( .A(n_936), .Y(n_981) );
INVxp67_ASAP7_75t_SL g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g973 ( .A(n_942), .Y(n_973) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVxp67_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVxp67_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI21xp5_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_986), .B(n_987), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_991), .Y(n_990) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_994), .Y(n_1015) );
OR2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_1004), .Y(n_994) );
NAND4xp25_ASAP7_75t_L g995 ( .A(n_996), .B(n_999), .C(n_1001), .D(n_1002), .Y(n_995) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
NAND4xp25_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .C(n_1007), .D(n_1008), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1015), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
endmodule