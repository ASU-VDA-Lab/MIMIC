module fake_netlist_1_2339_n_27 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_7;
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
BUFx10_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
OAI22xp33_ASAP7_75t_SL g10 ( .A1(n_2), .A2(n_0), .B1(n_6), .B2(n_3), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx2_ASAP7_75t_SL g12 ( .A(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_9), .B(n_0), .Y(n_14) );
OAI21x1_ASAP7_75t_L g15 ( .A1(n_7), .A2(n_1), .B(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_8), .B(n_12), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_8), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_18), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_17), .Y(n_22) );
NOR3xp33_ASAP7_75t_L g23 ( .A(n_21), .B(n_10), .C(n_16), .Y(n_23) );
OAI211xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_16), .B(n_12), .C(n_20), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_14), .B1(n_15), .B2(n_24), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
XNOR2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_15), .Y(n_27) );
endmodule