module real_jpeg_33905_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_0),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_0),
.Y(n_366)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_0),
.Y(n_384)
);

INVx2_ASAP7_75t_R g87 ( 
.A(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_1),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_1),
.B(n_364),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_14),
.B1(n_203),
.B2(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_41),
.Y(n_40)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_3),
.B(n_134),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_4),
.B(n_177),
.Y(n_569)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_5),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_5),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_5),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_5),
.B(n_501),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_9),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_9),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_9),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_9),
.B(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_9),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_12),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_12),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_77),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_12),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_28),
.Y(n_197)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_13),
.Y(n_155)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

NAND2x1_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_14),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_14),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_14),
.B(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_14),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_14),
.B(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_14),
.B(n_517),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_15),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_16),
.B(n_33),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_16),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_16),
.B(n_151),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_16),
.B(n_245),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_16),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_16),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_16),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_16),
.B(n_513),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_17),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_567),
.C(n_570),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_179),
.Y(n_19)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.C(n_175),
.Y(n_20)
);

NOR4xp25_ASAP7_75t_L g573 ( 
.A(n_21),
.B(n_113),
.C(n_175),
.D(n_571),
.Y(n_573)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_22),
.B(n_177),
.Y(n_568)
);

AO21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_71),
.B(n_112),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_71),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_51),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_50),
.Y(n_24)
);

CKINVDCx11_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.C(n_36),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_27),
.A2(n_36),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_27),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_27),
.A2(n_55),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_30),
.Y(n_405)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_30),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_32),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

XOR2x2_ASAP7_75t_L g120 ( 
.A(n_31),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_32),
.B(n_122),
.C(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_35),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_R g44 ( 
.A1(n_36),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_44),
.B2(n_49),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_63),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_40),
.A2(n_49),
.B1(n_75),
.B2(n_76),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_42),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_42),
.Y(n_151)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_45),
.A2(n_46),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_45),
.A2(n_46),
.B1(n_157),
.B2(n_158),
.Y(n_346)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_46),
.B(n_147),
.C(n_157),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_46),
.B(n_288),
.C(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_47),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_48),
.B(n_258),
.C(n_261),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_48),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_61),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_62),
.C(n_66),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

NAND2x1_ASAP7_75t_SL g122 ( 
.A(n_58),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_58),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_58),
.B(n_381),
.Y(n_380)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g249 ( 
.A(n_60),
.Y(n_249)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_62),
.A2(n_63),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_62),
.B(n_236),
.C(n_240),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_62),
.A2(n_63),
.B1(n_240),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_65),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_65),
.Y(n_459)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_132),
.C(n_135),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_66),
.A2(n_67),
.B1(n_135),
.B2(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_70),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_108),
.C(n_109),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_72),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_93),
.C(n_106),
.Y(n_72)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_73),
.B(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_80),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_81),
.C(n_86),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_76),
.B1(n_139),
.B2(n_145),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_75),
.B(n_132),
.C(n_143),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_75),
.A2(n_76),
.B1(n_313),
.B2(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_76),
.B(n_309),
.C(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_79),
.Y(n_447)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_79),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_85),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_87),
.B(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_93),
.B(n_106),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_102),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_98),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_99),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_99),
.A2(n_163),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_99),
.B(n_148),
.C(n_273),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_99),
.B(n_148),
.C(n_273),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_101),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_101),
.Y(n_287)
);

XOR2x2_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_108),
.B(n_109),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g567 ( 
.A1(n_113),
.A2(n_568),
.B(n_569),
.Y(n_567)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_173),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_115),
.B(n_173),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_164),
.C(n_171),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_117),
.B(n_547),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_146),
.C(n_161),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_118),
.B(n_550),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_131),
.C(n_138),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_120),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_126),
.A2(n_127),
.B1(n_231),
.B2(n_234),
.Y(n_230)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_127),
.B(n_227),
.C(n_234),
.Y(n_275)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_131),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_132),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_132),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_132),
.B(n_198),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_132),
.A2(n_144),
.B1(n_198),
.B2(n_199),
.Y(n_449)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_133),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_134),
.Y(n_525)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_135),
.Y(n_267)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_138),
.Y(n_336)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_146),
.B(n_161),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_147),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_148),
.B(n_150),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_148),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_148),
.B(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_148),
.B(n_439),
.Y(n_475)
);

INVx8_ASAP7_75t_L g471 ( 
.A(n_149),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_152),
.B(n_244),
.C(n_248),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_152),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_152),
.A2(n_244),
.B1(n_254),
.B2(n_375),
.Y(n_374)
);

OR2x2_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_155),
.Y(n_264)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_164),
.B(n_171),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_165),
.B(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_168),
.B(n_169),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI31xp33_ASAP7_75t_L g570 ( 
.A1(n_180),
.A2(n_568),
.A3(n_571),
.B(n_573),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_544),
.B(n_564),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_423),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_349),
.B(n_419),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g423 ( 
.A(n_184),
.B(n_424),
.C(n_542),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_290),
.B1(n_327),
.B2(n_330),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_186),
.B(n_291),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_251),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_188),
.B(n_268),
.C(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_209),
.C(n_224),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_190),
.A2(n_191),
.B1(n_210),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_201),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_205),
.C(n_208),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.C(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_193),
.A2(n_198),
.B1(n_199),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_200),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_206),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_210),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_217),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_211),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_211),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_216),
.B(n_218),
.Y(n_301)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_223),
.Y(n_499)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_225),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_235),
.C(n_243),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_226),
.B(n_243),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2x2_ASAP7_75t_L g385 ( 
.A(n_235),
.B(n_386),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_239),
.Y(n_442)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_248),
.B(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_250),
.B(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_250),
.B(n_528),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_268),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_252),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_253),
.B(n_257),
.C(n_265),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_263),
.Y(n_529)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_279),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_280),
.C(n_289),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.C(n_276),
.Y(n_269)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_273),
.B(n_315),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_289),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_319),
.C(n_323),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_292),
.B(n_353),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_303),
.B(n_318),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_298),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_299),
.Y(n_357)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OA21x2_ASAP7_75t_SL g376 ( 
.A1(n_300),
.A2(n_377),
.B(n_380),
.Y(n_376)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_305),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_308),
.B(n_314),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_309),
.B(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_311),
.Y(n_501)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_354),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_331),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_328),
.B(n_331),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_332),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_339),
.B2(n_348),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_334),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_347),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_344),
.B2(n_345),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_342),
.B(n_555),
.C(n_556),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_344),
.Y(n_556)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g555 ( 
.A(n_347),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_348),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_387),
.B(n_418),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_351),
.B(n_543),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_352),
.B(n_355),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.C(n_385),
.Y(n_355)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_373),
.C(n_376),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.C(n_367),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_360),
.A2(n_361),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_362),
.A2(n_363),
.B1(n_367),
.B2(n_368),
.Y(n_435)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_365),
.B(n_457),
.Y(n_521)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx12f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_376),
.Y(n_394)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_390),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_392),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_388),
.B(n_392),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_416),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_416),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_399),
.C(n_414),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_399),
.A2(n_414),
.B1(n_415),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_406),
.C(n_409),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_400),
.A2(n_401),
.B1(n_409),
.B2(n_410),
.Y(n_483)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_406),
.B(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B(n_422),
.Y(n_419)
);

AO21x1_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_450),
.B(n_541),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_426),
.B(n_428),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_433),
.C(n_436),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_430),
.B(n_539),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_433),
.B(n_436),
.Y(n_539)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_443),
.C(n_448),
.Y(n_436)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_437),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_441),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_443),
.A2(n_448),
.B1(n_449),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_443),
.Y(n_487)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_535),
.B(n_540),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_490),
.B(n_534),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_476),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_453),
.B(n_476),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_467),
.C(n_475),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_454),
.B(n_503),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_464),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_460),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_464),
.C(n_480),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_460),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_467),
.A2(n_468),
.B1(n_475),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_469),
.A2(n_472),
.B1(n_473),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_469),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_475),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_484),
.B1(n_488),
.B2(n_489),
.Y(n_476)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_477),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_481),
.B2(n_482),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_479),
.B(n_489),
.C(n_537),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_484),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_505),
.B(n_533),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_502),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_502),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_496),
.C(n_500),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_494),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_496),
.B(n_500),
.Y(n_509)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_519),
.B(n_532),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_510),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_510),
.Y(n_532)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_515),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_511),
.A2(n_512),
.B1(n_515),
.B2(n_516),
.Y(n_530)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_526),
.B(n_531),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_530),
.Y(n_531)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_538),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_538),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_557),
.Y(n_544)
);

AOI21x1_ASAP7_75t_SL g564 ( 
.A1(n_545),
.A2(n_565),
.B(n_566),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_548),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_548),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_551),
.C(n_553),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_551),
.Y(n_559)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_559),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_560),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_SL g565 ( 
.A(n_558),
.B(n_560),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_562),
.C(n_563),
.Y(n_560)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);


endmodule