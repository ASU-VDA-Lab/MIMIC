module fake_jpeg_16922_n_248 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_37),
.Y(n_39)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_44),
.B1(n_49),
.B2(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_36),
.B1(n_24),
.B2(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_26),
.B1(n_28),
.B2(n_15),
.Y(n_49)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_55),
.B(n_56),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_29),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_70),
.B(n_50),
.C(n_35),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_34),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_29),
.C(n_19),
.Y(n_71)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_51),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_81),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_44),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_45),
.B1(n_70),
.B2(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_47),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_27),
.B1(n_23),
.B2(n_19),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_50),
.B(n_38),
.C(n_49),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_93),
.B(n_89),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_50),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_45),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_53),
.B(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_38),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_62),
.C(n_58),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_116),
.C(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_67),
.B1(n_54),
.B2(n_50),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_118),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_122),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_54),
.B1(n_45),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_119),
.B1(n_120),
.B2(n_82),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_65),
.B1(n_59),
.B2(n_62),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_65),
.B1(n_35),
.B2(n_23),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_18),
.B1(n_17),
.B2(n_27),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_81),
.B1(n_77),
.B2(n_15),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_21),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_92),
.B(n_83),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_21),
.A3(n_18),
.B1(n_17),
.B2(n_23),
.Y(n_126)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.C(n_17),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_18),
.C(n_17),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_95),
.B1(n_104),
.B2(n_113),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_131),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_136),
.B(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_142),
.B1(n_144),
.B2(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_87),
.B1(n_91),
.B2(n_97),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_94),
.B(n_84),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_97),
.B1(n_99),
.B2(n_94),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_84),
.C(n_78),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_95),
.C(n_8),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_97),
.B1(n_78),
.B2(n_82),
.Y(n_148)
);

FAx1_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_118),
.CI(n_107),
.CON(n_161),
.SN(n_161)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_78),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_154),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_6),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_116),
.B(n_118),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_152),
.B(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_144),
.B(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_167),
.C(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_95),
.C(n_8),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_5),
.C(n_12),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_5),
.C(n_12),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_176),
.C(n_9),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_4),
.C(n_11),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_152),
.B1(n_153),
.B2(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_188),
.B1(n_190),
.B2(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_191),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_148),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_162),
.C(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_134),
.B1(n_145),
.B2(n_137),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_149),
.B1(n_130),
.B2(n_151),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_131),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_149),
.B1(n_9),
.B2(n_3),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_158),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_203),
.Y(n_209)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_161),
.C(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_161),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_174),
.B(n_156),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_205),
.A2(n_198),
.B1(n_193),
.B2(n_202),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_164),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_177),
.C(n_168),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.C(n_185),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_165),
.C(n_175),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_214),
.C(n_200),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_205),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_199),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_197),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_184),
.B1(n_182),
.B2(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_197),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_226),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_214),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_208),
.B1(n_155),
.B2(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_184),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_155),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_207),
.B(n_206),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_169),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_170),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_209),
.B(n_176),
.C(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_233),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_235),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_3),
.B(n_11),
.C(n_13),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_221),
.B1(n_220),
.B2(n_222),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_229),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_3),
.C(n_13),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_0),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_242),
.A3(n_243),
.B1(n_236),
.B2(n_238),
.C1(n_2),
.C2(n_0),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_1),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_1),
.Y(n_248)
);


endmodule