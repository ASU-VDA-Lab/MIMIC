module real_jpeg_6429_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_1),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_122),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_45),
.B1(n_119),
.B2(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_27),
.C(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_84),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_96),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_69),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_6),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_7),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_34),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_9),
.A2(n_43),
.B1(n_86),
.B2(n_89),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_9),
.A2(n_43),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

XNOR2x2_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_154),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_152),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_90),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_90),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_56),
.C(n_66),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_15),
.A2(n_16),
.B1(n_56),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_28),
.B(n_38),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_24),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_25),
.Y(n_169)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_28),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_93)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx5_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_47)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_33),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_33),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_39),
.B(n_96),
.Y(n_162)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_42),
.Y(n_146)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_56),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_66),
.B(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_75),
.B(n_82),
.Y(n_66)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_75),
.A2(n_82),
.B(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_85),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_76),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_129),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_101),
.B2(n_102),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_94),
.A2(n_158),
.B(n_162),
.Y(n_157)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_116),
.B(n_123),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_114),
.Y(n_105)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_119),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_142),
.A3(n_143),
.B1(n_147),
.B2(n_150),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_139),
.B(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_184),
.B(n_190),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_173),
.B(n_205),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_170),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_157),
.A2(n_163),
.B1(n_164),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_195),
.B(n_204),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_182),
.B(n_194),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_193),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_202),
.Y(n_204)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);


endmodule