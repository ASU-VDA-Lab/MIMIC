module fake_jpeg_1089_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_3),
.B(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_14),
.A2(n_6),
.B1(n_10),
.B2(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_8),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_8),
.B(n_6),
.C(n_10),
.D(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_13),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_22),
.B(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_23),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_26),
.B1(n_28),
.B2(n_7),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_35),
.C(n_15),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_37),
.C(n_11),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.C(n_11),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_1),
.Y(n_39)
);


endmodule