module fake_jpeg_828_n_220 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_220);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_53),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_76),
.B1(n_74),
.B2(n_64),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_67),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_99),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_76),
.B1(n_77),
.B2(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_97),
.B1(n_54),
.B2(n_52),
.Y(n_101)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_62),
.B1(n_75),
.B2(n_57),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_109),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_96),
.B1(n_63),
.B2(n_67),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_59),
.B(n_55),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_105),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_64),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_75),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_113),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_70),
.B1(n_58),
.B2(n_59),
.Y(n_111)
);

OAI22x1_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_96),
.B1(n_71),
.B2(n_69),
.Y(n_134)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_66),
.B1(n_73),
.B2(n_70),
.Y(n_115)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_134),
.B1(n_10),
.B2(n_11),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_62),
.A3(n_73),
.B1(n_52),
.B2(n_77),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_8),
.B(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_50),
.C(n_49),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_111),
.Y(n_143)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_145),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_104),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_153),
.C(n_156),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_101),
.B1(n_117),
.B2(n_115),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_152),
.B1(n_161),
.B2(n_14),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_4),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_115),
.B1(n_6),
.B2(n_7),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_44),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_43),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_158),
.B(n_17),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_5),
.B(n_7),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_8),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_34),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_164),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_131),
.B(n_128),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_134),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_120),
.B(n_13),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_12),
.B(n_13),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_12),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_15),
.B(n_17),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_23),
.B(n_30),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_184),
.C(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_184),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_173),
.A2(n_157),
.B1(n_160),
.B2(n_156),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_177),
.B1(n_172),
.B2(n_181),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_148),
.C(n_24),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_178),
.C(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_170),
.B1(n_165),
.B2(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

AOI31xp67_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_202),
.A3(n_204),
.B(n_193),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_168),
.C(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_176),
.B1(n_174),
.B2(n_181),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_168),
.C(n_175),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_188),
.C(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_195),
.C(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_21),
.C(n_28),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_192),
.CI(n_193),
.CON(n_208),
.SN(n_208)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_208),
.A2(n_209),
.B(n_204),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_211),
.B(n_206),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_206),
.C(n_207),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_215),
.B(n_208),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_20),
.B(n_26),
.C(n_33),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_19),
.B(n_18),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_18),
.Y(n_220)
);


endmodule