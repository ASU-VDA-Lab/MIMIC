module fake_netlist_6_870_n_1652 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1652);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1652;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_63),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_5),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_72),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_74),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_115),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_64),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_53),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_19),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_49),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_51),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_94),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_120),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_56),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_107),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_150),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_24),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_162),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_102),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_133),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_46),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_96),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_1),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_26),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_12),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_3),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_108),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_77),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_13),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_124),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_33),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_34),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_101),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_49),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_30),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_122),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_155),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_24),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_114),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_144),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_105),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_160),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_97),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_141),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_45),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_13),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_55),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_28),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_43),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_60),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_151),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_167),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_38),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_145),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_38),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_111),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_157),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_73),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_67),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_165),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_118),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_9),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_68),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_76),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_136),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_121),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_21),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_41),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_103),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_42),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_28),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_149),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_46),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_86),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_50),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_128),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_18),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_21),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_11),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_35),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_78),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_3),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_129),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_26),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_39),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_83),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_31),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_87),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_55),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_66),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_15),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_109),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_91),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_71),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_132),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_104),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_36),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_93),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_48),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_79),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_4),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_58),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_32),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_202),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_204),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_2),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_243),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_210),
.B(n_6),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_228),
.B(n_7),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_187),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_175),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_262),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_228),
.B(n_7),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_199),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_208),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_203),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_205),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_179),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_210),
.B(n_8),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_211),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_262),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_212),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_201),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_215),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_201),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_216),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_201),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_219),
.B(n_8),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_201),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_233),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_201),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_285),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_218),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_226),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_226),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_231),
.B(n_11),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_226),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_313),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_224),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_225),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_266),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_232),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_244),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_247),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_249),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_251),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_226),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_174),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_253),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_231),
.B(n_14),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_175),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_226),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_264),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_254),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_219),
.B(n_14),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_246),
.B(n_16),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_270),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_254),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_271),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_254),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_254),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_301),
.B(n_16),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_254),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_185),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_176),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_190),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_206),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_192),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_213),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_272),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_206),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_273),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_222),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_274),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_246),
.B(n_17),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_276),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_238),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_278),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_185),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_259),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_261),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_315),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_340),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_345),
.B(n_315),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_332),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_342),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_343),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_344),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_328),
.A2(n_230),
.B(n_180),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_355),
.B(n_169),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_333),
.A2(n_230),
.B(n_180),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_R g429 ( 
.A(n_329),
.B(n_280),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_348),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_345),
.B(n_169),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_350),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_359),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_359),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_363),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_393),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_172),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_352),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_358),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_354),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_361),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_362),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_368),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_335),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_369),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

AND2x2_ASAP7_75t_SL g454 ( 
.A(n_379),
.B(n_268),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_336),
.A2(n_279),
.B(n_268),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_371),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_372),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_393),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_397),
.B(n_170),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_336),
.A2(n_341),
.B(n_337),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_383),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_401),
.B(n_236),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_401),
.B(n_236),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_373),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_374),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_375),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_389),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_337),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_386),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_388),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_346),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_325),
.B(n_240),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_382),
.B(n_293),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_346),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_432),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_454),
.A2(n_330),
.B1(n_347),
.B2(n_384),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_279),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_356),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_314),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_L g493 ( 
.A1(n_436),
.A2(n_326),
.B1(n_405),
.B2(n_220),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_400),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_454),
.B(n_470),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_334),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_421),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_465),
.A2(n_385),
.B1(n_331),
.B2(n_339),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_470),
.A2(n_404),
.B1(n_408),
.B2(n_402),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_432),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_464),
.B(n_314),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_465),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_441),
.B(n_426),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_436),
.B(n_406),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_419),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_416),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_450),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_476),
.B(n_172),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_476),
.B(n_172),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_172),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_465),
.A2(n_365),
.B1(n_392),
.B2(n_380),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_443),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_426),
.B(n_334),
.Y(n_522)
);

INVx4_ASAP7_75t_SL g523 ( 
.A(n_441),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_415),
.A2(n_370),
.B1(n_294),
.B2(n_260),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_417),
.B(n_380),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_478),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_443),
.Y(n_528)
);

INVx4_ASAP7_75t_SL g529 ( 
.A(n_441),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_465),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_441),
.B(n_485),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_476),
.B(n_172),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_424),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_423),
.B(n_409),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_486),
.B(n_184),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_429),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_441),
.B(n_349),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_441),
.B(n_477),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_443),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_477),
.B(n_349),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_412),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_477),
.B(n_240),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_484),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_395),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_439),
.B(n_440),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_430),
.B(n_327),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_484),
.B(n_184),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_418),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_418),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_424),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_481),
.B(n_338),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_413),
.B(n_267),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_487),
.B(n_184),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_463),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_463),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_420),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g565 ( 
.A(n_433),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_442),
.B(n_184),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_424),
.B(n_184),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_439),
.B(n_440),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_439),
.B(n_177),
.Y(n_572)
);

INVx4_ASAP7_75t_SL g573 ( 
.A(n_487),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_439),
.B(n_235),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_487),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_445),
.A2(n_239),
.B1(n_299),
.B2(n_237),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_440),
.B(n_248),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_422),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_446),
.B(n_391),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_444),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_447),
.B(n_377),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_448),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_425),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_424),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_451),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_460),
.B(n_395),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_463),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_425),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_427),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_461),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_463),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_471),
.A2(n_234),
.B1(n_275),
.B2(n_209),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_427),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_458),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_472),
.B(n_183),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_435),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_455),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_428),
.B(n_396),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_428),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_473),
.B(n_193),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_482),
.B(n_411),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_483),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_437),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_437),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_483),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_458),
.A2(n_367),
.B1(n_195),
.B2(n_191),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_438),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_480),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_480),
.B(n_197),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_438),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_449),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_452),
.B(n_396),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_479),
.B(n_200),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_453),
.B(n_295),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_456),
.B(n_398),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_457),
.B(n_411),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_459),
.B(n_398),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_496),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_490),
.B(n_263),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_548),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_548),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_602),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_536),
.B(n_182),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_495),
.B(n_494),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_522),
.B(n_462),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_522),
.B(n_462),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_498),
.B(n_196),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_585),
.B(n_290),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_530),
.A2(n_296),
.B1(n_305),
.B2(n_300),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_581),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_500),
.B(n_466),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_508),
.B(n_263),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_508),
.B(n_263),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_530),
.A2(n_292),
.B1(n_258),
.B2(n_242),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_466),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_488),
.Y(n_638)
);

OAI22xp33_ASAP7_75t_L g639 ( 
.A1(n_558),
.A2(n_324),
.B1(n_297),
.B2(n_286),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_207),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_580),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_599),
.Y(n_642)
);

A2O1A1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_489),
.A2(n_399),
.B(n_410),
.C(n_407),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_531),
.B(n_263),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_580),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_490),
.B(n_263),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_510),
.B(n_170),
.Y(n_648)
);

AND2x2_ASAP7_75t_SL g649 ( 
.A(n_518),
.B(n_223),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_604),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_536),
.B(n_467),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_510),
.B(n_227),
.C(n_245),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_504),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g654 ( 
.A(n_556),
.B(n_399),
.C(n_410),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_600),
.B(n_250),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_598),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_609),
.B(n_467),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_468),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_619),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_594),
.B(n_468),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_594),
.B(n_475),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_606),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_565),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_597),
.B(n_252),
.Y(n_664)
);

BUFx5_ASAP7_75t_L g665 ( 
.A(n_568),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_497),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_506),
.A2(n_568),
.B1(n_555),
.B2(n_533),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_600),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_509),
.B(n_269),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_595),
.B(n_171),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_597),
.B(n_277),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_607),
.B(n_287),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_612),
.B(n_289),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_600),
.B(n_316),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_537),
.B(n_317),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_499),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_595),
.B(n_171),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_526),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_539),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_601),
.B(n_173),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_490),
.A2(n_302),
.B1(n_321),
.B2(n_319),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_572),
.B(n_574),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_577),
.B(n_173),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_521),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_497),
.B(n_501),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_497),
.B(n_178),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_601),
.B(n_181),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_534),
.B(n_403),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_541),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_490),
.B(n_181),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_590),
.B(n_186),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_492),
.A2(n_491),
.B1(n_557),
.B2(n_556),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_544),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_497),
.B(n_501),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_553),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_492),
.B(n_188),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_553),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_554),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_191),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_501),
.B(n_523),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_554),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_616),
.B(n_195),
.Y(n_703)
);

NOR2x1p5_ASAP7_75t_L g704 ( 
.A(n_551),
.B(n_189),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_555),
.B(n_304),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_561),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_558),
.B(n_403),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_561),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_584),
.B(n_304),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_564),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_565),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_567),
.B(n_307),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_598),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_564),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_507),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_501),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_491),
.A2(n_307),
.B1(n_309),
.B2(n_321),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_584),
.B(n_311),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_608),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_613),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_608),
.B(n_319),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_571),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_517),
.A2(n_323),
.B1(n_320),
.B2(n_318),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_578),
.B(n_214),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_523),
.B(n_217),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_491),
.A2(n_283),
.B1(n_229),
.B2(n_241),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_491),
.A2(n_284),
.B1(n_255),
.B2(n_256),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_579),
.A2(n_288),
.B1(n_257),
.B2(n_265),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_576),
.B(n_323),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_583),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_517),
.A2(n_320),
.B1(n_318),
.B2(n_312),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_558),
.A2(n_312),
.B1(n_310),
.B2(n_308),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_583),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_588),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_588),
.B(n_291),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_529),
.B(n_298),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_529),
.B(n_282),
.Y(n_737)
);

BUFx6f_ASAP7_75t_SL g738 ( 
.A(n_507),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_589),
.B(n_593),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_589),
.B(n_281),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_535),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_596),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_596),
.B(n_605),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_605),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_535),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_549),
.B(n_306),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_517),
.B(n_306),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_503),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_579),
.A2(n_303),
.B1(n_198),
.B2(n_194),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_636),
.B(n_723),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_623),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_SL g752 ( 
.A1(n_634),
.A2(n_532),
.B(n_515),
.C(n_516),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_660),
.A2(n_569),
.B(n_538),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_622),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_640),
.B(n_532),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_646),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_640),
.B(n_517),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_648),
.B(n_513),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_689),
.B(n_502),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_626),
.A2(n_648),
.B1(n_649),
.B2(n_624),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_627),
.B(n_517),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_670),
.A2(n_680),
.B(n_687),
.C(n_677),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_643),
.A2(n_610),
.B(n_493),
.C(n_545),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_676),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_634),
.A2(n_575),
.B(n_546),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_670),
.A2(n_617),
.B(n_614),
.C(n_525),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_628),
.B(n_649),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_668),
.A2(n_547),
.B(n_560),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_667),
.B(n_613),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_667),
.A2(n_613),
.B1(n_592),
.B2(n_542),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_620),
.B(n_563),
.Y(n_771)
);

OAI21xp33_ASAP7_75t_L g772 ( 
.A1(n_629),
.A2(n_303),
.B(n_505),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_623),
.A2(n_570),
.B(n_566),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_646),
.A2(n_566),
.B(n_552),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_677),
.A2(n_527),
.B(n_512),
.C(n_520),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_646),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_679),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_633),
.A2(n_566),
.B(n_552),
.Y(n_778)
);

OAI321xp33_ASAP7_75t_L g779 ( 
.A1(n_732),
.A2(n_514),
.A3(n_18),
.B1(n_22),
.B2(n_23),
.C(n_25),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_688),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_656),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_665),
.A2(n_615),
.B1(n_519),
.B2(n_587),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_674),
.A2(n_519),
.B(n_543),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_672),
.A2(n_519),
.B(n_587),
.C(n_528),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_707),
.B(n_562),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_674),
.A2(n_562),
.B(n_543),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_642),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_641),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_629),
.B(n_528),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_741),
.B(n_528),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_663),
.B(n_540),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_745),
.B(n_543),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_721),
.B(n_507),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_680),
.B(n_587),
.C(n_562),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_721),
.B(n_511),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_720),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_693),
.A2(n_524),
.B1(n_550),
.B2(n_591),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_662),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_720),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_665),
.B(n_615),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_672),
.A2(n_615),
.B1(n_550),
.B2(n_559),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_632),
.B(n_511),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_685),
.A2(n_573),
.B(n_559),
.Y(n_803)
);

OA22x2_ASAP7_75t_L g804 ( 
.A1(n_749),
.A2(n_511),
.B1(n_582),
.B2(n_23),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_661),
.A2(n_559),
.B(n_582),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_695),
.A2(n_559),
.B(n_65),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_695),
.A2(n_716),
.B(n_664),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_665),
.A2(n_61),
.B1(n_161),
.B2(n_159),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_665),
.B(n_637),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_665),
.B(n_651),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_659),
.B(n_17),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_690),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_671),
.A2(n_666),
.B(n_739),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_635),
.A2(n_164),
.B(n_152),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_665),
.B(n_22),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_635),
.A2(n_147),
.B(n_140),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_657),
.B(n_27),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_707),
.B(n_139),
.Y(n_818)
);

AO21x1_ASAP7_75t_L g819 ( 
.A1(n_669),
.A2(n_29),
.B(n_30),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_666),
.A2(n_134),
.B(n_130),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_645),
.Y(n_821)
);

BUFx4f_ASAP7_75t_L g822 ( 
.A(n_678),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_687),
.A2(n_126),
.B1(n_125),
.B2(n_123),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_743),
.A2(n_106),
.B(n_99),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_700),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_700),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_712),
.A2(n_98),
.B1(n_92),
.B2(n_88),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_712),
.A2(n_75),
.B1(n_69),
.B2(n_44),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_658),
.B(n_40),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_625),
.B(n_43),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_644),
.A2(n_44),
.B(n_47),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_696),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_713),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_701),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_683),
.B(n_48),
.Y(n_835)
);

CKINVDCx8_ASAP7_75t_R g836 ( 
.A(n_711),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_644),
.A2(n_51),
.B(n_52),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_669),
.A2(n_54),
.B(n_57),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_650),
.B(n_59),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_723),
.A2(n_731),
.B1(n_729),
.B2(n_707),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_652),
.B(n_719),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_705),
.A2(n_709),
.B1(n_718),
.B2(n_697),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_703),
.B(n_694),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_728),
.B(n_654),
.C(n_727),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_699),
.B(n_702),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_706),
.A2(n_714),
.B(n_722),
.C(n_733),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_621),
.A2(n_647),
.B(n_691),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_698),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_734),
.B(n_708),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_710),
.B(n_744),
.Y(n_850)
);

NOR2x1_ASAP7_75t_R g851 ( 
.A(n_715),
.B(n_686),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_630),
.B(n_692),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_675),
.A2(n_725),
.B(n_737),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_736),
.A2(n_742),
.B(n_730),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_630),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_638),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_748),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_681),
.A2(n_731),
.B1(n_726),
.B2(n_747),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_746),
.A2(n_686),
.B1(n_724),
.B2(n_740),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_639),
.B(n_717),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_735),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_704),
.B(n_673),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_653),
.A2(n_684),
.B(n_655),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_655),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_738),
.A2(n_495),
.B1(n_640),
.B2(n_626),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_640),
.B(n_648),
.Y(n_866)
);

CKINVDCx8_ASAP7_75t_R g867 ( 
.A(n_663),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_624),
.B(n_693),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_668),
.A2(n_508),
.B(n_594),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_646),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_689),
.B(n_620),
.Y(n_871)
);

OAI21xp33_ASAP7_75t_L g872 ( 
.A1(n_640),
.A2(n_648),
.B(n_629),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_646),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_640),
.A2(n_495),
.B1(n_626),
.B2(n_648),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_667),
.A2(n_626),
.B1(n_495),
.B2(n_640),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_646),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_640),
.A2(n_648),
.B(n_677),
.C(n_670),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_640),
.A2(n_648),
.B(n_677),
.C(n_670),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_640),
.A2(n_495),
.B1(n_626),
.B2(n_648),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_682),
.B(n_640),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_624),
.B(n_693),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_688),
.B(n_581),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_682),
.B(n_640),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_640),
.A2(n_495),
.B1(n_626),
.B2(n_648),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_682),
.B(n_640),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_667),
.A2(n_508),
.B(n_626),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_682),
.B(n_640),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_682),
.B(n_640),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_624),
.B(n_693),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_682),
.B(n_640),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_636),
.A2(n_631),
.B1(n_649),
.B2(n_667),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_682),
.B(n_640),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_667),
.A2(n_626),
.B1(n_495),
.B2(n_640),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_663),
.B(n_585),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_640),
.B(n_648),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_636),
.A2(n_631),
.B1(n_649),
.B2(n_667),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_622),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_640),
.A2(n_648),
.B(n_677),
.C(n_670),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_764),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_780),
.B(n_880),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_788),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_756),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_833),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_894),
.B(n_802),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_754),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_842),
.A2(n_893),
.B(n_875),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_783),
.A2(n_753),
.B(n_807),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_836),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_813),
.A2(n_752),
.B(n_886),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_866),
.B(n_895),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_872),
.A2(n_891),
.B(n_896),
.C(n_884),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_756),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_886),
.A2(n_885),
.B(n_883),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_867),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_887),
.B(n_888),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_890),
.A2(n_892),
.B(n_853),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_793),
.B(n_795),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_755),
.A2(n_809),
.B(n_778),
.Y(n_920)
);

AOI21xp33_ASAP7_75t_L g921 ( 
.A1(n_750),
.A2(n_860),
.B(n_758),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_874),
.B(n_879),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_781),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_756),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_863),
.A2(n_774),
.B(n_869),
.Y(n_925)
);

BUFx6f_ASAP7_75t_SL g926 ( 
.A(n_821),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_760),
.B(n_865),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_SL g928 ( 
.A(n_891),
.B(n_896),
.Y(n_928)
);

AND2x2_ASAP7_75t_SL g929 ( 
.A(n_825),
.B(n_767),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_818),
.B(n_798),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_882),
.B(n_780),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_785),
.B(n_871),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_810),
.A2(n_789),
.B(n_800),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_861),
.B(n_766),
.Y(n_934)
);

AO31x2_ASAP7_75t_L g935 ( 
.A1(n_775),
.A2(n_819),
.A3(n_846),
.B(n_770),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_785),
.B(n_871),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_818),
.B(n_864),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_776),
.B(n_870),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_843),
.B(n_817),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_829),
.B(n_859),
.Y(n_941)
);

AOI21xp33_ASAP7_75t_L g942 ( 
.A1(n_840),
.A2(n_858),
.B(n_844),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_815),
.A2(n_757),
.B(n_840),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_759),
.B(n_811),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_897),
.B(n_835),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_768),
.A2(n_784),
.B(n_773),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_776),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_759),
.B(n_868),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_889),
.B(n_881),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_856),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_772),
.B(n_812),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_870),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_769),
.A2(n_761),
.B1(n_751),
.B2(n_782),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_845),
.A2(n_797),
.B(n_805),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_870),
.B(n_876),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_777),
.B(n_841),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_751),
.B(n_834),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_822),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_803),
.A2(n_792),
.B(n_790),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_794),
.A2(n_850),
.B(n_849),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_814),
.A2(n_816),
.B(n_763),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_857),
.B(n_771),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_771),
.B(n_852),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_855),
.B(n_822),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_873),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_830),
.B(n_839),
.C(n_838),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_814),
.A2(n_816),
.B(n_831),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_873),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_876),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_801),
.A2(n_862),
.B(n_848),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_862),
.B(n_804),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_832),
.B(n_796),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_832),
.A2(n_837),
.B(n_820),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_791),
.B(n_796),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_799),
.B(n_834),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_799),
.B(n_834),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_824),
.A2(n_806),
.B(n_808),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_779),
.A2(n_826),
.B1(n_828),
.B2(n_823),
.C(n_827),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_804),
.A2(n_851),
.B(n_779),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_866),
.B(n_895),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_847),
.A2(n_668),
.B(n_762),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_866),
.B(n_895),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_780),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_787),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_877),
.B(n_878),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_882),
.B(n_780),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_756),
.Y(n_993)
);

OAI21x1_ASAP7_75t_SL g994 ( 
.A1(n_814),
.A2(n_816),
.B(n_819),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_866),
.B(n_895),
.Y(n_995)
);

OAI21x1_ASAP7_75t_SL g996 ( 
.A1(n_814),
.A2(n_816),
.B(n_819),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_866),
.A2(n_895),
.B(n_877),
.C(n_878),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_866),
.A2(n_895),
.B(n_877),
.C(n_878),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_836),
.B(n_416),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_866),
.B(n_895),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_754),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_866),
.B(n_895),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_764),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_756),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_866),
.B(n_895),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_875),
.A2(n_893),
.A3(n_878),
.B(n_877),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_1010)
);

INVx3_ASAP7_75t_SL g1011 ( 
.A(n_759),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_882),
.B(n_780),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_788),
.Y(n_1013)
);

OR2x2_ASAP7_75t_SL g1014 ( 
.A(n_844),
.B(n_417),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_866),
.B(n_895),
.Y(n_1015)
);

OAI22x1_ASAP7_75t_L g1016 ( 
.A1(n_860),
.A2(n_895),
.B1(n_866),
.B2(n_795),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_836),
.B(n_565),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_833),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_866),
.A2(n_895),
.B1(n_872),
.B2(n_878),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_877),
.A2(n_898),
.B(n_878),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_866),
.B(n_895),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_756),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_847),
.A2(n_668),
.B(n_762),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_756),
.B(n_646),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_765),
.A2(n_854),
.B(n_786),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_764),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_900),
.B(n_912),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_902),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_931),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_932),
.B(n_936),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_903),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_SL g1034 ( 
.A(n_914),
.B(n_968),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_981),
.A2(n_1022),
.B1(n_1015),
.B2(n_1008),
.Y(n_1035)
);

NAND2x2_ASAP7_75t_L g1036 ( 
.A(n_902),
.B(n_958),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_944),
.B(n_981),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1022),
.B(n_992),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_932),
.B(n_936),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_916),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_SL g1041 ( 
.A(n_921),
.B(n_997),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_SL g1042 ( 
.A1(n_990),
.A2(n_942),
.B(n_982),
.C(n_988),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_986),
.B(n_995),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1000),
.B(n_1003),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_917),
.B(n_1020),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1013),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_1016),
.A2(n_928),
.B1(n_966),
.B2(n_929),
.Y(n_1047)
);

CKINVDCx6p67_ASAP7_75t_R g1048 ( 
.A(n_926),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_997),
.B(n_998),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_998),
.B(n_922),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_915),
.B(n_940),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_918),
.A2(n_920),
.B(n_961),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_961),
.A2(n_991),
.B(n_904),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_929),
.A2(n_1001),
.B1(n_1018),
.B2(n_1005),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_919),
.B(n_915),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_903),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_903),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1012),
.B(n_948),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_913),
.A2(n_978),
.B1(n_990),
.B2(n_908),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_956),
.B(n_1017),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_937),
.B(n_930),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_903),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1011),
.B(n_948),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_934),
.B(n_949),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1002),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_914),
.B(n_968),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_938),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_938),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1011),
.B(n_987),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_927),
.A2(n_1021),
.B1(n_971),
.B2(n_908),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_910),
.B(n_923),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_999),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_945),
.B(n_956),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_913),
.B(n_927),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1021),
.A2(n_967),
.B1(n_994),
.B2(n_996),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_999),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_906),
.B(n_963),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_941),
.A2(n_987),
.B1(n_943),
.B2(n_951),
.C(n_1006),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_899),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_L g1080 ( 
.A(n_989),
.B(n_950),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_962),
.B(n_1009),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1028),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_972),
.Y(n_1083)
);

OAI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_937),
.A2(n_930),
.B1(n_975),
.B2(n_976),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_947),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_SL g1086 ( 
.A(n_969),
.B(n_957),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1009),
.B(n_979),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_926),
.Y(n_1088)
);

AO21x1_ASAP7_75t_L g1089 ( 
.A1(n_953),
.A2(n_983),
.B(n_1024),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_905),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_937),
.B(n_930),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_970),
.A2(n_974),
.B1(n_964),
.B2(n_957),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_974),
.B(n_969),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_965),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_924),
.B(n_993),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_1014),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_970),
.A2(n_960),
.B1(n_911),
.B2(n_947),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1019),
.A2(n_977),
.B1(n_1023),
.B2(n_1009),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1009),
.B(n_993),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_L g1100 ( 
.A(n_965),
.B(n_1007),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_965),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1023),
.B(n_952),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_939),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_939),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_924),
.B(n_952),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_1025),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1025),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_965),
.B(n_1007),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1007),
.B(n_955),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_935),
.B(n_1007),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_973),
.B(n_925),
.Y(n_1111)
);

AND2x6_ASAP7_75t_L g1112 ( 
.A(n_935),
.B(n_954),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_959),
.B(n_946),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_935),
.B(n_933),
.Y(n_1114)
);

BUFx8_ASAP7_75t_L g1115 ( 
.A(n_901),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_980),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_984),
.B(n_985),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1004),
.A2(n_1010),
.B1(n_1026),
.B2(n_1027),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_909),
.B(n_900),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_903),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_903),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_944),
.B(n_882),
.Y(n_1122)
);

BUFx2_ASAP7_75t_SL g1123 ( 
.A(n_926),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_907),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_932),
.B(n_936),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_903),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_987),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_SL g1128 ( 
.A(n_910),
.B(n_836),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_907),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_981),
.B(n_1022),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_932),
.B(n_936),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_944),
.B(n_882),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_932),
.B(n_936),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_981),
.A2(n_866),
.B(n_895),
.C(n_878),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_981),
.A2(n_1022),
.B1(n_986),
.B2(n_995),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_932),
.B(n_936),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_999),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_899),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_981),
.B(n_1022),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_981),
.A2(n_895),
.B1(n_866),
.B2(n_1022),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_987),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_981),
.A2(n_1022),
.B1(n_986),
.B2(n_995),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_L g1143 ( 
.A(n_997),
.B(n_762),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_981),
.B(n_1022),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_SL g1145 ( 
.A(n_902),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_944),
.B(n_882),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_931),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_932),
.B(n_936),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_981),
.B(n_1022),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_944),
.B(n_882),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_932),
.B(n_936),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_937),
.B(n_930),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_931),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_902),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_937),
.B(n_930),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_944),
.B(n_882),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1065),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1110),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1140),
.B(n_1139),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1110),
.Y(n_1160)
);

AOI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1134),
.A2(n_1143),
.B(n_1135),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1087),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1061),
.B(n_1091),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1092),
.B(n_1099),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1115),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1127),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1124),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1115),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1141),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1129),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1054),
.A2(n_1047),
.B1(n_1041),
.B2(n_1035),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1092),
.B(n_1119),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1173)
);

BUFx2_ASAP7_75t_R g1174 ( 
.A(n_1090),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1035),
.A2(n_1135),
.B1(n_1142),
.B2(n_1041),
.Y(n_1175)
);

AO21x1_ASAP7_75t_L g1176 ( 
.A1(n_1059),
.A2(n_1053),
.B(n_1074),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1154),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_1082),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1081),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1059),
.A2(n_1130),
.B1(n_1096),
.B2(n_1074),
.Y(n_1180)
);

INVxp33_ASAP7_75t_L g1181 ( 
.A(n_1069),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_SL g1182 ( 
.A(n_1079),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1114),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1038),
.B(n_1037),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1114),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1097),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1130),
.A2(n_1044),
.B1(n_1043),
.B2(n_1073),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1096),
.A2(n_1053),
.B1(n_1060),
.B2(n_1045),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1138),
.Y(n_1189)
);

INVx8_ASAP7_75t_L g1190 ( 
.A(n_1033),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1031),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_1145),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1044),
.A2(n_1029),
.B1(n_1058),
.B2(n_1045),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1031),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1147),
.B(n_1153),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1063),
.A2(n_1049),
.B1(n_1122),
.B2(n_1146),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1040),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1147),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1049),
.A2(n_1156),
.B1(n_1132),
.B2(n_1150),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1050),
.A2(n_1078),
.B1(n_1070),
.B2(n_1098),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1050),
.A2(n_1064),
.B1(n_1153),
.B2(n_1077),
.Y(n_1201)
);

AO21x2_ASAP7_75t_L g1202 ( 
.A1(n_1052),
.A2(n_1117),
.B(n_1089),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1085),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1145),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1033),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1083),
.Y(n_1206)
);

BUFx8_ASAP7_75t_L g1207 ( 
.A(n_1061),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1084),
.A2(n_1091),
.B1(n_1155),
.B2(n_1152),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1093),
.B(n_1109),
.Y(n_1209)
);

BUFx8_ASAP7_75t_L g1210 ( 
.A(n_1032),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1046),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1048),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1093),
.B(n_1155),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1108),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1152),
.A2(n_1155),
.B1(n_1055),
.B2(n_1051),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1097),
.A2(n_1075),
.B(n_1118),
.Y(n_1216)
);

CKINVDCx6p67_ASAP7_75t_R g1217 ( 
.A(n_1123),
.Y(n_1217)
);

AO21x1_ASAP7_75t_SL g1218 ( 
.A1(n_1051),
.A2(n_1042),
.B(n_1104),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1105),
.B(n_1102),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1072),
.A2(n_1076),
.B1(n_1137),
.B2(n_1152),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1080),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_1113),
.A2(n_1086),
.B(n_1111),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1107),
.B(n_1068),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1112),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1057),
.B(n_1121),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1032),
.B(n_1151),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1103),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1068),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1066),
.Y(n_1229)
);

OAI21xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1106),
.A2(n_1121),
.B(n_1126),
.Y(n_1230)
);

CKINVDCx16_ASAP7_75t_R g1231 ( 
.A(n_1039),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1066),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1039),
.B(n_1136),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1030),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1125),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1112),
.A2(n_1095),
.B(n_1133),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1112),
.A2(n_1100),
.B(n_1034),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1112),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1131),
.Y(n_1239)
);

CKINVDCx12_ASAP7_75t_R g1240 ( 
.A(n_1128),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1095),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1036),
.A2(n_1071),
.B1(n_1133),
.B2(n_1131),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1088),
.A2(n_1101),
.B1(n_1067),
.B2(n_1148),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1056),
.A2(n_1062),
.B1(n_1094),
.B2(n_1120),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1101),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1056),
.A2(n_1120),
.B1(n_1062),
.B2(n_1094),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1094),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1120),
.Y(n_1248)
);

BUFx2_ASAP7_75t_SL g1249 ( 
.A(n_1033),
.Y(n_1249)
);

BUFx2_ASAP7_75t_R g1250 ( 
.A(n_1090),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1154),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1140),
.A2(n_895),
.B1(n_866),
.B2(n_981),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1059),
.A2(n_895),
.B(n_866),
.Y(n_1253)
);

BUFx2_ASAP7_75t_R g1254 ( 
.A(n_1090),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1081),
.B(n_1074),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1127),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1140),
.B(n_981),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1040),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1145),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1115),
.Y(n_1260)
);

BUFx2_ASAP7_75t_R g1261 ( 
.A(n_1090),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1140),
.B(n_981),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1110),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1088),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1255),
.B(n_1179),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1181),
.B(n_1159),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1177),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1255),
.B(n_1158),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1158),
.B(n_1160),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1236),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1186),
.Y(n_1271)
);

INVxp33_ASAP7_75t_L g1272 ( 
.A(n_1182),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1197),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1191),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1253),
.A2(n_1161),
.B(n_1176),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1213),
.B(n_1163),
.Y(n_1276)
);

CKINVDCx14_ASAP7_75t_R g1277 ( 
.A(n_1197),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1236),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1173),
.B(n_1184),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1236),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1224),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1263),
.B(n_1175),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1252),
.A2(n_1171),
.B1(n_1196),
.B2(n_1199),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1162),
.B(n_1164),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1176),
.A2(n_1183),
.A3(n_1185),
.B(n_1238),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1198),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1162),
.B(n_1164),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1224),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1166),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1258),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_L g1291 ( 
.A(n_1190),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1222),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1216),
.A2(n_1172),
.B(n_1168),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1177),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1172),
.B(n_1238),
.Y(n_1295)
);

NAND2x1_ASAP7_75t_L g1296 ( 
.A(n_1224),
.B(n_1165),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1202),
.A2(n_1193),
.B(n_1187),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1203),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1195),
.B(n_1188),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1256),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1169),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1202),
.A2(n_1222),
.B(n_1237),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1206),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1216),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1219),
.Y(n_1305)
);

AO21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1200),
.A2(n_1208),
.B(n_1215),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1202),
.B(n_1216),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1194),
.B(n_1214),
.Y(n_1308)
);

NAND2xp33_ASAP7_75t_R g1309 ( 
.A(n_1204),
.B(n_1165),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1157),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1230),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1237),
.A2(n_1262),
.B(n_1257),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1167),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1170),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1190),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1180),
.B(n_1201),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1223),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1184),
.B(n_1165),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1227),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1237),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1218),
.B(n_1223),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1258),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1189),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1218),
.B(n_1163),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1228),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1163),
.B(n_1209),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1225),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1225),
.B(n_1209),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1168),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1168),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1247),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1296),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1281),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1281),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1285),
.B(n_1260),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1285),
.B(n_1260),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1285),
.B(n_1248),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1288),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1270),
.B(n_1213),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1285),
.B(n_1278),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1285),
.B(n_1248),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1265),
.B(n_1243),
.Y(n_1342)
);

OAI211xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1283),
.A2(n_1178),
.B(n_1220),
.C(n_1221),
.Y(n_1343)
);

AND2x4_ASAP7_75t_SL g1344 ( 
.A(n_1295),
.B(n_1213),
.Y(n_1344)
);

NOR2x1_ASAP7_75t_L g1345 ( 
.A(n_1312),
.B(n_1249),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1265),
.B(n_1241),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1311),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1280),
.B(n_1209),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1316),
.B(n_1232),
.Y(n_1349)
);

NOR2x1p5_ASAP7_75t_L g1350 ( 
.A(n_1316),
.B(n_1259),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1299),
.A2(n_1231),
.B1(n_1259),
.B2(n_1217),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1311),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1280),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1268),
.B(n_1232),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1288),
.Y(n_1355)
);

OAI33xp33_ASAP7_75t_L g1356 ( 
.A1(n_1308),
.A2(n_1242),
.A3(n_1204),
.B1(n_1245),
.B2(n_1226),
.B3(n_1240),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1304),
.B(n_1234),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1324),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1284),
.B(n_1239),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1324),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1300),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1306),
.A2(n_1207),
.B1(n_1233),
.B2(n_1210),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1312),
.B(n_1235),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1312),
.B(n_1307),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_SL g1365 ( 
.A(n_1282),
.B(n_1205),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1302),
.B(n_1233),
.Y(n_1366)
);

NOR2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1322),
.B(n_1217),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1287),
.B(n_1229),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1300),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1343),
.B(n_1275),
.C(n_1266),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1358),
.B(n_1295),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1346),
.B(n_1274),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1338),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1346),
.B(n_1286),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1358),
.B(n_1295),
.Y(n_1375)
);

AOI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1356),
.A2(n_1279),
.B1(n_1289),
.B2(n_1301),
.C(n_1323),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1351),
.B(n_1272),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1351),
.B(n_1276),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1354),
.B(n_1305),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1362),
.B(n_1276),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1349),
.A2(n_1277),
.B(n_1282),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1350),
.A2(n_1273),
.B1(n_1290),
.B2(n_1318),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1347),
.B(n_1276),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1350),
.A2(n_1273),
.B1(n_1290),
.B2(n_1295),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1347),
.B(n_1322),
.Y(n_1385)
);

OAI21xp33_ASAP7_75t_L g1386 ( 
.A1(n_1349),
.A2(n_1347),
.B(n_1342),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1345),
.A2(n_1330),
.B(n_1329),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1360),
.B(n_1366),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1360),
.B(n_1321),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1360),
.B(n_1268),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1347),
.A2(n_1309),
.B1(n_1326),
.B2(n_1291),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1369),
.B(n_1317),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1359),
.B(n_1240),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1366),
.B(n_1320),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1369),
.B(n_1303),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1344),
.A2(n_1306),
.B(n_1328),
.Y(n_1396)
);

NOR3xp33_ASAP7_75t_L g1397 ( 
.A(n_1356),
.B(n_1315),
.C(n_1308),
.Y(n_1397)
);

NOR3xp33_ASAP7_75t_L g1398 ( 
.A(n_1345),
.B(n_1315),
.C(n_1229),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1361),
.B(n_1271),
.Y(n_1399)
);

AOI211xp5_ASAP7_75t_L g1400 ( 
.A1(n_1335),
.A2(n_1294),
.B(n_1267),
.C(n_1313),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1357),
.B(n_1298),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1365),
.A2(n_1327),
.B1(n_1297),
.B2(n_1331),
.C(n_1314),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1357),
.B(n_1319),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_SL g1404 ( 
.A(n_1352),
.B(n_1314),
.C(n_1310),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1366),
.B(n_1292),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1335),
.B(n_1310),
.C(n_1207),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1352),
.A2(n_1267),
.B1(n_1294),
.B2(n_1251),
.C(n_1211),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1348),
.A2(n_1207),
.B1(n_1328),
.B2(n_1297),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1368),
.B(n_1269),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1348),
.A2(n_1297),
.B1(n_1210),
.B2(n_1327),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1373),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1373),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1388),
.B(n_1340),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1403),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1388),
.B(n_1340),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1405),
.B(n_1340),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1394),
.B(n_1333),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1405),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1409),
.B(n_1372),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1374),
.B(n_1333),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1401),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1392),
.B(n_1333),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1371),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1390),
.B(n_1336),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1395),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1399),
.Y(n_1426)
);

AND2x4_ASAP7_75t_SL g1427 ( 
.A(n_1398),
.B(n_1339),
.Y(n_1427)
);

AOI33xp33_ASAP7_75t_L g1428 ( 
.A1(n_1376),
.A2(n_1336),
.A3(n_1364),
.B1(n_1337),
.B2(n_1341),
.B3(n_1363),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1383),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1389),
.B(n_1352),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1371),
.Y(n_1431)
);

AND2x4_ASAP7_75t_SL g1432 ( 
.A(n_1375),
.B(n_1339),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1386),
.B(n_1337),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1386),
.B(n_1337),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1370),
.B(n_1341),
.C(n_1325),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1379),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1387),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1404),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1402),
.B(n_1341),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1407),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1437),
.B(n_1338),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1439),
.B(n_1365),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1418),
.B(n_1400),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1418),
.B(n_1400),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1432),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1439),
.B(n_1365),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1437),
.B(n_1421),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1411),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1411),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1438),
.B(n_1365),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1334),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1416),
.B(n_1353),
.Y(n_1452)
);

OR3x2_ASAP7_75t_L g1453 ( 
.A(n_1428),
.B(n_1367),
.C(n_1250),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1413),
.B(n_1353),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1412),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1412),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1414),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1427),
.B(n_1332),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1438),
.B(n_1355),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1414),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1413),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1413),
.B(n_1353),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1415),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1426),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1421),
.B(n_1355),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1426),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1440),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1415),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1425),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1432),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1415),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1417),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1461),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1461),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1458),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1448),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1467),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1435),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1442),
.B(n_1433),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1442),
.B(n_1440),
.Y(n_1481)
);

OAI32xp33_ASAP7_75t_L g1482 ( 
.A1(n_1442),
.A2(n_1434),
.A3(n_1433),
.B1(n_1435),
.B2(n_1429),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1430),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1446),
.B(n_1429),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1427),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1446),
.A2(n_1434),
.B1(n_1381),
.B2(n_1370),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1443),
.B(n_1430),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1446),
.B(n_1419),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1449),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1443),
.B(n_1430),
.Y(n_1491)
);

NAND2x2_ASAP7_75t_L g1492 ( 
.A(n_1445),
.B(n_1367),
.Y(n_1492)
);

A2O1A1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1453),
.A2(n_1381),
.B(n_1377),
.C(n_1396),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1445),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1455),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1419),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1469),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1455),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1455),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1455),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1472),
.B(n_1420),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1453),
.A2(n_1396),
.B1(n_1406),
.B2(n_1384),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1470),
.A2(n_1406),
.B1(n_1408),
.B2(n_1410),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1472),
.B(n_1420),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1447),
.B(n_1422),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1447),
.B(n_1425),
.Y(n_1509)
);

AND2x2_ASAP7_75t_SL g1510 ( 
.A(n_1450),
.B(n_1397),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1470),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1456),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1431),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1450),
.B(n_1436),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_1469),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1480),
.B(n_1464),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1500),
.B(n_1461),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1498),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1473),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1500),
.B(n_1461),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1476),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1489),
.B(n_1459),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1510),
.B(n_1466),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1487),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1494),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1514),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1481),
.B(n_1466),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1478),
.A2(n_1391),
.B1(n_1382),
.B2(n_1378),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1486),
.B(n_1450),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1474),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1507),
.B(n_1463),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1489),
.B(n_1459),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1490),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1507),
.B(n_1463),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1512),
.B(n_1463),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1493),
.A2(n_1431),
.B1(n_1385),
.B2(n_1423),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1508),
.B(n_1459),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1494),
.B(n_1463),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_SL g1542 ( 
.A(n_1493),
.B(n_1174),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1483),
.B(n_1457),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1474),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1514),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1512),
.B(n_1468),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1495),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1441),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1488),
.B(n_1457),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1496),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1545),
.B(n_1488),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1541),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1523),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1523),
.Y(n_1557)
);

AOI321xp33_ASAP7_75t_L g1558 ( 
.A1(n_1532),
.A2(n_1482),
.A3(n_1504),
.B1(n_1484),
.B2(n_1505),
.C(n_1478),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1491),
.Y(n_1559)
);

OAI31xp33_ASAP7_75t_L g1560 ( 
.A1(n_1542),
.A2(n_1511),
.A3(n_1479),
.B(n_1485),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1531),
.A2(n_1492),
.B1(n_1539),
.B2(n_1526),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1528),
.B(n_1518),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1542),
.A2(n_1511),
.B(n_1479),
.C(n_1515),
.Y(n_1563)
);

AO22x2_ASAP7_75t_L g1564 ( 
.A1(n_1520),
.A2(n_1475),
.B1(n_1485),
.B2(n_1513),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1531),
.A2(n_1492),
.B1(n_1485),
.B2(n_1475),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1524),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1530),
.A2(n_1509),
.B(n_1441),
.Y(n_1567)
);

AOI322xp5_ASAP7_75t_L g1568 ( 
.A1(n_1520),
.A2(n_1468),
.A3(n_1471),
.B1(n_1462),
.B2(n_1454),
.C1(n_1452),
.C2(n_1451),
.Y(n_1568)
);

AND2x2_ASAP7_75t_SL g1569 ( 
.A(n_1516),
.B(n_1291),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1517),
.B(n_1503),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1527),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1524),
.A2(n_1535),
.B1(n_1540),
.B2(n_1475),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1535),
.B(n_1212),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1527),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1506),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1536),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1541),
.B(n_1458),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1564),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1552),
.B(n_1573),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1558),
.B(n_1540),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1573),
.B(n_1541),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1566),
.B(n_1550),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1556),
.B(n_1547),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1554),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1557),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1536),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1561),
.B(n_1212),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1559),
.B(n_1548),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1555),
.B(n_1548),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1565),
.B(n_1264),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1571),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1563),
.A2(n_1522),
.B(n_1519),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1564),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1576),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1574),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1553),
.B(n_1547),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1587),
.A2(n_1572),
.B(n_1574),
.Y(n_1598)
);

O2A1O1Ixp5_ASAP7_75t_L g1599 ( 
.A1(n_1580),
.A2(n_1577),
.B(n_1553),
.C(n_1575),
.Y(n_1599)
);

OAI211xp5_ASAP7_75t_L g1600 ( 
.A1(n_1586),
.A2(n_1560),
.B(n_1568),
.C(n_1577),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1594),
.A2(n_1567),
.B1(n_1570),
.B2(n_1551),
.C(n_1519),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1593),
.A2(n_1569),
.B(n_1549),
.Y(n_1602)
);

NAND4xp25_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1549),
.C(n_1538),
.D(n_1522),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1581),
.B(n_1569),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1578),
.Y(n_1605)
);

AOI222xp33_ASAP7_75t_L g1606 ( 
.A1(n_1594),
.A2(n_1546),
.B1(n_1534),
.B2(n_1538),
.C1(n_1537),
.C2(n_1551),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1578),
.A2(n_1546),
.B1(n_1534),
.B2(n_1537),
.C(n_1544),
.Y(n_1607)
);

NAND4xp75_ASAP7_75t_L g1608 ( 
.A(n_1596),
.B(n_1590),
.C(n_1579),
.D(n_1581),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1591),
.A2(n_1583),
.B1(n_1590),
.B2(n_1597),
.Y(n_1609)
);

AOI211xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1589),
.A2(n_1544),
.B(n_1521),
.C(n_1525),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1605),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_L g1612 ( 
.A(n_1608),
.B(n_1588),
.C(n_1592),
.Y(n_1612)
);

XOR2xp5_ASAP7_75t_L g1613 ( 
.A(n_1609),
.B(n_1582),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1604),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1598),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1600),
.A2(n_1583),
.B1(n_1597),
.B2(n_1582),
.Y(n_1616)
);

AOI211x1_ASAP7_75t_L g1617 ( 
.A1(n_1602),
.A2(n_1595),
.B(n_1585),
.C(n_1584),
.Y(n_1617)
);

NOR4xp25_ASAP7_75t_L g1618 ( 
.A(n_1601),
.B(n_1595),
.C(n_1585),
.D(n_1584),
.Y(n_1618)
);

NOR2x1_ASAP7_75t_L g1619 ( 
.A(n_1603),
.B(n_1521),
.Y(n_1619)
);

AND4x1_ASAP7_75t_L g1620 ( 
.A(n_1599),
.B(n_1606),
.C(n_1610),
.D(n_1607),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_L g1621 ( 
.A(n_1608),
.B(n_1521),
.Y(n_1621)
);

NAND4xp25_ASAP7_75t_L g1622 ( 
.A(n_1616),
.B(n_1544),
.C(n_1525),
.D(n_1533),
.Y(n_1622)
);

OA211x2_ASAP7_75t_L g1623 ( 
.A1(n_1615),
.A2(n_1393),
.B(n_1465),
.C(n_1380),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1620),
.A2(n_1533),
.B(n_1525),
.Y(n_1624)
);

NAND4xp25_ASAP7_75t_SL g1625 ( 
.A(n_1612),
.B(n_1533),
.C(n_1261),
.D(n_1254),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1614),
.Y(n_1626)
);

OR3x1_ASAP7_75t_L g1627 ( 
.A(n_1625),
.B(n_1622),
.C(n_1611),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1626),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1624),
.A2(n_1613),
.B1(n_1621),
.B2(n_1618),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1623),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1626),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1626),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1631),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1628),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1632),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1629),
.B(n_1264),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1629),
.B(n_1619),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1637),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1633),
.Y(n_1639)
);

NOR2xp67_ASAP7_75t_SL g1640 ( 
.A(n_1634),
.B(n_1630),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1639),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1641),
.B(n_1635),
.Y(n_1642)
);

AOI221x1_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1640),
.B1(n_1638),
.B2(n_1636),
.C(n_1627),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1642),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1644),
.B(n_1617),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1643),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1645),
.A2(n_1211),
.B(n_1499),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1646),
.A2(n_1502),
.B1(n_1501),
.B2(n_1471),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1647),
.A2(n_1251),
.B(n_1192),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1649),
.B(n_1648),
.C(n_1192),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_R g1651 ( 
.A1(n_1650),
.A2(n_1192),
.B1(n_1190),
.B2(n_1244),
.C(n_1246),
.Y(n_1651)
);

OAI31xp33_ASAP7_75t_L g1652 ( 
.A1(n_1651),
.A2(n_1205),
.A3(n_1460),
.B(n_1456),
.Y(n_1652)
);


endmodule