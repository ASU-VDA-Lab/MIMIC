module fake_aes_2552_n_667 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_667);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_667;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_19), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_44), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_21), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_58), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_41), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_4), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_63), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_38), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_31), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_42), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_55), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_22), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_33), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_40), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_32), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_39), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_13), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_16), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_64), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_68), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
NOR2xp67_ASAP7_75t_L g100 ( .A(n_6), .B(n_65), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_23), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_69), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_61), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_28), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_60), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_26), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_25), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_56), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_15), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_9), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_70), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_54), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_67), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_9), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_20), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_30), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_53), .Y(n_121) );
AND2x6_ASAP7_75t_L g122 ( .A(n_121), .B(n_24), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g123 ( .A(n_121), .B(n_0), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_121), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_83), .B(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_75), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_111), .B(n_1), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_102), .B(n_1), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_94), .B(n_2), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_102), .B(n_2), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_95), .B(n_3), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_87), .Y(n_146) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_88), .A2(n_35), .B(n_66), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_94), .B(n_3), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_95), .B(n_4), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_90), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_91), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_91), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_92), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_101), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_128), .B(n_103), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_135), .A2(n_80), .B1(n_118), .B2(n_113), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_128), .B(n_117), .Y(n_164) );
INVx2_ASAP7_75t_SL g165 ( .A(n_143), .Y(n_165) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_135), .B(n_101), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_129), .A2(n_109), .B(n_115), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_129), .B(n_80), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_135), .A2(n_120), .B1(n_85), .B2(n_112), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
NOR2x1p5_ASAP7_75t_L g171 ( .A(n_127), .B(n_117), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_143), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
OAI221xp5_ASAP7_75t_L g175 ( .A1(n_131), .A2(n_97), .B1(n_105), .B2(n_106), .C(n_109), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_131), .B(n_99), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_134), .B(n_114), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_134), .B(n_114), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_136), .B(n_120), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_136), .B(n_137), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_137), .B(n_96), .Y(n_183) );
NAND3xp33_ASAP7_75t_L g184 ( .A(n_132), .B(n_116), .C(n_98), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_139), .A2(n_76), .B1(n_108), .B2(n_107), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_139), .B(n_77), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_141), .B(n_85), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_141), .B(n_104), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_150), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_148), .A2(n_81), .B1(n_78), .B2(n_93), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_130), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_144), .B(n_119), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_124), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_130), .Y(n_194) );
NOR2xp33_ASAP7_75t_SL g195 ( .A(n_122), .B(n_100), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_143), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_144), .B(n_5), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_124), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_149), .B(n_36), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_149), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_153), .B(n_7), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_153), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_154), .B(n_8), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_154), .A2(n_155), .B1(n_160), .B2(n_156), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_122), .B(n_45), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_155), .B(n_10), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_160), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_125), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_122), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g212 ( .A(n_133), .B(n_12), .C(n_14), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_123), .A2(n_14), .B(n_15), .C(n_18), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_142), .B(n_34), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_142), .B(n_37), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_145), .B(n_43), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_125), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_145), .B(n_47), .Y(n_219) );
NOR2xp67_ASAP7_75t_L g220 ( .A(n_146), .B(n_48), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_208), .B(n_146), .Y(n_221) );
INVx5_ASAP7_75t_L g222 ( .A(n_210), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_200), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_166), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_189), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_181), .B(n_157), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_213), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_182), .A2(n_152), .B(n_157), .C(n_125), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_187), .B(n_138), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_173), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_164), .B(n_122), .Y(n_235) );
AND3x2_ASAP7_75t_SL g236 ( .A(n_189), .B(n_126), .C(n_122), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_165), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_179), .B(n_122), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_185), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_166), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_176), .B(n_122), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_210), .Y(n_242) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_206), .B(n_147), .Y(n_243) );
AOI211xp5_ASAP7_75t_L g244 ( .A1(n_175), .A2(n_126), .B(n_130), .C(n_151), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_173), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_180), .B(n_151), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_171), .B(n_151), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_193), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g249 ( .A(n_211), .B(n_161), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_162), .B(n_151), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_168), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_210), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_170), .A2(n_161), .B(n_159), .C(n_158), .Y(n_254) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_205), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_168), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_174), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_185), .B(n_201), .Y(n_258) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_192), .B(n_147), .Y(n_259) );
BUFx4f_ASAP7_75t_L g260 ( .A(n_217), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_169), .A2(n_147), .B1(n_159), .B2(n_158), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_190), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_192), .B(n_161), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_165), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_163), .B(n_147), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_203), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_167), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_178), .B(n_161), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_174), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_214), .B(n_202), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_218), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_218), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_178), .B(n_161), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_204), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_191), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_172), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_207), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_191), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_212), .Y(n_281) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_172), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_242), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_224), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_281), .B(n_195), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g286 ( .A(n_244), .B(n_206), .C(n_184), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_239), .Y(n_287) );
O2A1O1Ixp5_ASAP7_75t_L g288 ( .A1(n_267), .A2(n_183), .B(n_188), .C(n_186), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_235), .A2(n_196), .B(n_215), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_252), .B(n_183), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_238), .A2(n_196), .B(n_216), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_225), .B(n_188), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_256), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_242), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_226), .B(n_240), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_226), .B(n_186), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_252), .Y(n_297) );
AO21x1_ASAP7_75t_L g298 ( .A1(n_249), .A2(n_199), .B(n_219), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_227), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_276), .B(n_220), .Y(n_300) );
AND2x6_ASAP7_75t_L g301 ( .A(n_241), .B(n_194), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_233), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_241), .A2(n_199), .B(n_194), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_223), .Y(n_304) );
INVx8_ASAP7_75t_L g305 ( .A(n_258), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g306 ( .A1(n_226), .A2(n_159), .B1(n_158), .B2(n_51), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_262), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_241), .A2(n_159), .B(n_158), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_234), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_240), .B(n_49), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_240), .B(n_255), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_260), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_247), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_269), .A2(n_260), .B1(n_258), .B2(n_279), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_242), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_247), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_260), .A2(n_158), .B(n_159), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_231), .B(n_71), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_242), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_230), .A2(n_50), .B(n_52), .C(n_57), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_251), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_263), .B(n_62), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_247), .B(n_258), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_221), .B(n_228), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_272), .B(n_274), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_243), .A2(n_259), .B(n_246), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_258), .A2(n_229), .B1(n_272), .B2(n_249), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_326), .B(n_229), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_305), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_328), .A2(n_261), .B(n_270), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_284), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_298), .A2(n_278), .B(n_243), .Y(n_336) );
AO31x2_ASAP7_75t_L g337 ( .A1(n_327), .A2(n_230), .A3(n_254), .B(n_250), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_311), .B(n_273), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_323), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_315), .B(n_263), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_323), .Y(n_342) );
AO21x2_ASAP7_75t_L g343 ( .A1(n_327), .A2(n_254), .B(n_275), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_311), .B(n_253), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_283), .Y(n_347) );
NAND2x1_ASAP7_75t_L g348 ( .A(n_283), .B(n_278), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_329), .A2(n_278), .B(n_275), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_322), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_283), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_302), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_287), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_320), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_331), .B(n_311), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_332), .B(n_325), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_331), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_350), .B(n_293), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_335), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_346), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_330), .B(n_325), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_330), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_338), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_346), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_345), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_350), .B(n_296), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_342), .B(n_295), .Y(n_376) );
AO31x2_ASAP7_75t_L g377 ( .A1(n_338), .A2(n_314), .A3(n_285), .B(n_303), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_342), .B(n_295), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_346), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_357), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_346), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_353), .B(n_310), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_363), .B(n_355), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_381), .B(n_341), .C(n_299), .D(n_285), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_363), .B(n_355), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_381), .A2(n_227), .B(n_341), .C(n_324), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_384), .A2(n_305), .B1(n_329), .B2(n_325), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_371), .B(n_306), .C(n_318), .Y(n_390) );
INVx3_ASAP7_75t_SL g391 ( .A(n_362), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_360), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_361), .A2(n_268), .B1(n_305), .B2(n_310), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_361), .A2(n_268), .B1(n_310), .B2(n_297), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_368), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_373), .B(n_287), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_361), .A2(n_344), .B1(n_339), .B2(n_296), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_383), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_382), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_359), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_379), .A2(n_336), .B(n_349), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_321), .B(n_312), .C(n_349), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_384), .A2(n_339), .B1(n_344), .B2(n_296), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_379), .A2(n_336), .B(n_349), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_359), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_359), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_364), .B(n_292), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_369), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_369), .B(n_332), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_382), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_372), .B(n_337), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_369), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
NOR4xp75_ASAP7_75t_L g421 ( .A(n_389), .B(n_364), .C(n_374), .D(n_300), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_414), .B(n_375), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_385), .B(n_375), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_413), .B(n_377), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_395), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_385), .B(n_374), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_418), .B(n_370), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_400), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_418), .B(n_377), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_406), .B(n_377), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_387), .B(n_367), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_397), .B(n_377), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_417), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
AND2x4_ASAP7_75t_SL g435 ( .A(n_403), .B(n_362), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_387), .B(n_367), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_400), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_406), .B(n_377), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_411), .B(n_377), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_404), .B(n_378), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_415), .B(n_377), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_401), .B(n_379), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_419), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_419), .B(n_378), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_386), .B(n_378), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_407), .B(n_376), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_407), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_396), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_391), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_407), .B(n_376), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_407), .B(n_376), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_392), .B(n_337), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_416), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_394), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
NOR2x1p5_ASAP7_75t_SL g462 ( .A(n_417), .B(n_347), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_410), .B(n_380), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_393), .B(n_362), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_410), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_388), .A2(n_336), .B(n_286), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_410), .B(n_380), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_393), .B(n_362), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_391), .B(n_412), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_448), .B(n_391), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_452), .B(n_409), .Y(n_472) );
OAI31xp33_ASAP7_75t_L g473 ( .A1(n_449), .A2(n_408), .A3(n_390), .B(n_265), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_443), .B(n_399), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_422), .B(n_412), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_434), .B(n_402), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_445), .B(n_402), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_428), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_460), .B(n_343), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_428), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_457), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_437), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_448), .B(n_446), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_431), .B(n_380), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_454), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_423), .B(n_440), .Y(n_488) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_453), .B(n_420), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_466), .B(n_272), .C(n_265), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_470), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_445), .B(n_366), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_444), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_425), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_436), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_427), .B(n_366), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_444), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_461), .B(n_426), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_447), .Y(n_500) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_435), .A2(n_265), .A3(n_312), .B(n_313), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_458), .Y(n_503) );
INVxp67_ASAP7_75t_L g504 ( .A(n_432), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_433), .B(n_370), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_435), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_450), .B(n_337), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_459), .B(n_370), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_450), .B(n_337), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_455), .B(n_366), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_464), .B(n_343), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_432), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_455), .Y(n_515) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_451), .B(n_370), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_456), .Y(n_517) );
OAI31xp33_ASAP7_75t_L g518 ( .A1(n_468), .A2(n_317), .A3(n_307), .B(n_290), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_456), .B(n_417), .Y(n_519) );
NAND2xp33_ASAP7_75t_L g520 ( .A(n_433), .B(n_417), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_424), .A2(n_288), .B1(n_308), .B2(n_273), .C(n_274), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_429), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_457), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_427), .B(n_382), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_427), .B(n_382), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_424), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_451), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
AOI211x1_ASAP7_75t_L g529 ( .A1(n_496), .A2(n_421), .B(n_465), .C(n_439), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_485), .B(n_438), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_522), .B(n_438), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_517), .B(n_433), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_491), .B(n_430), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_515), .B(n_467), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_522), .B(n_430), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_526), .B(n_439), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_488), .B(n_429), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_499), .B(n_467), .Y(n_538) );
NOR2xp33_ASAP7_75t_SL g539 ( .A(n_507), .B(n_433), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_506), .B(n_463), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_476), .B(n_463), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_504), .B(n_442), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_494), .B(n_442), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_495), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_487), .B(n_469), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_489), .B(n_469), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_482), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_479), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_481), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_504), .B(n_462), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_503), .B(n_343), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_471), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_483), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_484), .Y(n_554) );
NOR4xp25_ASAP7_75t_L g555 ( .A(n_475), .B(n_358), .C(n_352), .D(n_351), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_477), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_528), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_527), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_478), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_474), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_527), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_474), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_514), .B(n_462), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_513), .B(n_519), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_514), .B(n_337), .Y(n_566) );
INVxp33_ASAP7_75t_L g567 ( .A(n_516), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_480), .B(n_337), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_472), .B(n_343), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_480), .B(n_382), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_520), .A2(n_382), .B(n_348), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_493), .Y(n_572) );
AOI21xp33_ASAP7_75t_SL g573 ( .A1(n_518), .A2(n_236), .B(n_334), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_490), .A2(n_272), .B(n_319), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_474), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_493), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_512), .B(n_510), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_497), .B(n_334), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_498), .Y(n_579) );
NAND4xp25_ASAP7_75t_SL g580 ( .A(n_552), .B(n_501), .C(n_473), .D(n_508), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_573), .B(n_521), .C(n_509), .Y(n_581) );
OAI22xp33_ASAP7_75t_SL g582 ( .A1(n_532), .A2(n_511), .B1(n_492), .B2(n_512), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_544), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_550), .B(n_520), .C(n_505), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_560), .B(n_486), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_564), .B(n_523), .C(n_482), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_548), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_572), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_545), .B(n_523), .C(n_502), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_569), .A2(n_525), .B1(n_524), .B2(n_500), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_532), .B(n_334), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_577), .B(n_333), .Y(n_592) );
NAND5xp2_ASAP7_75t_L g593 ( .A(n_539), .B(n_236), .C(n_289), .D(n_291), .E(n_301), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_574), .B(n_334), .C(n_348), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_549), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_545), .B(n_356), .C(n_346), .Y(n_596) );
OA22x2_ASAP7_75t_L g597 ( .A1(n_563), .A2(n_333), .B1(n_347), .B2(n_354), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_561), .B(n_358), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g599 ( .A(n_533), .B(n_358), .C(n_351), .D(n_354), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_333), .Y(n_600) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_569), .A2(n_301), .B1(n_354), .B2(n_352), .C1(n_351), .C2(n_274), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_557), .B(n_352), .C(n_273), .Y(n_602) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_575), .B(n_346), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_565), .B(n_356), .Y(n_604) );
OAI321xp33_ASAP7_75t_L g605 ( .A1(n_566), .A2(n_356), .A3(n_264), .B1(n_242), .B2(n_257), .C(n_245), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_553), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_558), .B(n_546), .C(n_568), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_556), .B(n_356), .Y(n_608) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_546), .B(n_356), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_537), .B(n_356), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_572), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_565), .B(n_316), .Y(n_613) );
NAND2xp33_ASAP7_75t_L g614 ( .A(n_531), .B(n_301), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_583), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_588), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_580), .A2(n_534), .B1(n_538), .B2(n_541), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_587), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_607), .B(n_534), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_581), .A2(n_555), .B(n_567), .Y(n_620) );
NOR4xp75_ASAP7_75t_L g621 ( .A(n_592), .B(n_535), .C(n_540), .D(n_536), .Y(n_621) );
OAI21xp33_ASAP7_75t_SL g622 ( .A1(n_597), .A2(n_567), .B(n_576), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_598), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_585), .B(n_534), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_595), .B(n_542), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_606), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_591), .A2(n_571), .B(n_543), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_597), .A2(n_547), .B(n_570), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_603), .A2(n_562), .B(n_559), .Y(n_629) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_609), .A2(n_579), .B(n_547), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_590), .A2(n_529), .B1(n_578), .B2(n_551), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_610), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_586), .B(n_584), .C(n_589), .Y(n_633) );
AOI32xp33_ASAP7_75t_L g634 ( .A1(n_612), .A2(n_551), .A3(n_253), .B1(n_237), .B2(n_266), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_582), .B(n_222), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_592), .A2(n_253), .B1(n_264), .B2(n_222), .C(n_245), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_617), .A2(n_599), .B1(n_614), .B2(n_611), .Y(n_637) );
AND3x4_ASAP7_75t_L g638 ( .A(n_621), .B(n_594), .C(n_602), .Y(n_638) );
AND3x4_ASAP7_75t_L g639 ( .A(n_622), .B(n_593), .C(n_601), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g640 ( .A(n_633), .B(n_620), .C(n_634), .Y(n_640) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_619), .B(n_596), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_629), .A2(n_600), .B(n_605), .C(n_613), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_631), .A2(n_608), .B1(n_593), .B2(n_604), .C(n_264), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_625), .A2(n_264), .B1(n_222), .B2(n_282), .C(n_257), .Y(n_644) );
NAND2xp33_ASAP7_75t_SL g645 ( .A(n_630), .B(n_264), .Y(n_645) );
NOR2xp67_ASAP7_75t_L g646 ( .A(n_628), .B(n_222), .Y(n_646) );
AND3x4_ASAP7_75t_L g647 ( .A(n_624), .B(n_266), .C(n_237), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_615), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_618), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_640), .A2(n_635), .B(n_628), .C(n_623), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_648), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_645), .A2(n_616), .B1(n_627), .B2(n_632), .C(n_626), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_649), .B(n_636), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_641), .Y(n_654) );
OAI31xp33_ASAP7_75t_SL g655 ( .A1(n_643), .A2(n_301), .A3(n_282), .B(n_222), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_638), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_656), .B(n_644), .C(n_642), .Y(n_657) );
AOI321xp33_ASAP7_75t_L g658 ( .A1(n_654), .A2(n_637), .A3(n_639), .B1(n_647), .B2(n_646), .C(n_232), .Y(n_658) );
NOR4xp25_ASAP7_75t_L g659 ( .A(n_650), .B(n_232), .C(n_271), .D(n_277), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_652), .A2(n_301), .B(n_277), .C(n_280), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_657), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_658), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_659), .A2(n_655), .B1(n_653), .B2(n_651), .C(n_282), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_661), .A2(n_655), .B1(n_660), .B2(n_271), .Y(n_664) );
OR2x6_ASAP7_75t_L g665 ( .A(n_662), .B(n_280), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_665), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_663), .B(n_664), .Y(n_667) );
endmodule