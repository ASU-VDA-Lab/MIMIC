module real_aes_17940_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_848, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_848;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g115 ( .A(n_0), .B(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_1), .A2(n_4), .B1(n_148), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_2), .A2(n_43), .B1(n_155), .B2(n_191), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_3), .A2(n_24), .B1(n_191), .B2(n_233), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_5), .A2(n_16), .B1(n_145), .B2(n_222), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_6), .A2(n_62), .B1(n_205), .B2(n_235), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_7), .A2(n_17), .B1(n_155), .B2(n_176), .Y(n_627) );
INVx1_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_9), .A2(n_479), .B(n_836), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_10), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_11), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_12), .A2(n_18), .B1(n_204), .B2(n_207), .Y(n_203) );
BUFx2_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
OR2x2_ASAP7_75t_L g474 ( .A(n_13), .B(n_37), .Y(n_474) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_14), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_15), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_19), .A2(n_101), .B1(n_145), .B2(n_148), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_20), .A2(n_38), .B1(n_180), .B2(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_21), .B(n_146), .Y(n_177) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_22), .A2(n_58), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_23), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_25), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_26), .B(n_152), .Y(n_547) );
INVx4_ASAP7_75t_R g595 ( .A(n_27), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_28), .A2(n_48), .B1(n_193), .B2(n_194), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_29), .A2(n_55), .B1(n_145), .B2(n_194), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_30), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_31), .B(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_32), .Y(n_256) );
INVx1_ASAP7_75t_L g526 ( .A(n_33), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_34), .B(n_191), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_SL g538 ( .A1(n_35), .A2(n_151), .B(n_155), .C(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_36), .A2(n_56), .B1(n_155), .B2(n_194), .Y(n_515) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_39), .A2(n_88), .B1(n_155), .B2(n_232), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_40), .Y(n_844) );
XOR2x2_ASAP7_75t_L g829 ( .A(n_41), .B(n_830), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_42), .A2(n_46), .B1(n_155), .B2(n_176), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_44), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_45), .A2(n_60), .B1(n_145), .B2(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_47), .A2(n_74), .B1(n_831), .B2(n_832), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_47), .Y(n_832) );
INVx1_ASAP7_75t_L g550 ( .A(n_49), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_50), .B(n_155), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_51), .Y(n_567) );
INVx2_ASAP7_75t_L g487 ( .A(n_52), .Y(n_487) );
INVx1_ASAP7_75t_L g111 ( .A(n_53), .Y(n_111) );
BUFx3_ASAP7_75t_L g496 ( .A(n_53), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_54), .A2(n_124), .B(n_475), .Y(n_123) );
AOI31xp33_ASAP7_75t_L g475 ( .A1(n_54), .A2(n_476), .A3(n_478), .B(n_479), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_57), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_59), .A2(n_89), .B1(n_155), .B2(n_194), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_61), .A2(n_69), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_61), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_63), .A2(n_77), .B1(n_154), .B2(n_193), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_64), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_65), .A2(n_79), .B1(n_155), .B2(n_176), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_66), .A2(n_100), .B1(n_145), .B2(n_207), .Y(n_253) );
AND2x4_ASAP7_75t_L g141 ( .A(n_67), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g164 ( .A(n_68), .Y(n_164) );
INVx1_ASAP7_75t_L g127 ( .A(n_69), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_70), .A2(n_92), .B1(n_193), .B2(n_194), .Y(n_522) );
AO22x1_ASAP7_75t_L g584 ( .A1(n_71), .A2(n_78), .B1(n_219), .B2(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g142 ( .A(n_72), .Y(n_142) );
AND2x2_ASAP7_75t_L g542 ( .A(n_73), .B(n_186), .Y(n_542) );
INVx1_ASAP7_75t_L g831 ( .A(n_74), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_75), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_76), .B(n_235), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_80), .B(n_191), .Y(n_568) );
INVx2_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_82), .B(n_186), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_83), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_84), .A2(n_99), .B1(n_194), .B2(n_235), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_85), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_86), .B(n_162), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_87), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_90), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_91), .B(n_186), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_93), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_94), .B(n_186), .Y(n_564) );
INVx1_ASAP7_75t_L g114 ( .A(n_95), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_95), .B(n_472), .Y(n_471) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_96), .B(n_146), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_97), .A2(n_210), .B(n_235), .C(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g597 ( .A(n_98), .B(n_598), .Y(n_597) );
NAND2xp33_ASAP7_75t_L g572 ( .A(n_102), .B(n_181), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_122), .B(n_843), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx4_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx8_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_117), .Y(n_107) );
OR2x6_ASAP7_75t_L g846 ( .A(n_108), .B(n_117), .Y(n_846) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g472 ( .A(n_111), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g502 ( .A(n_114), .Y(n_502) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_483), .B(n_488), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_468), .Y(n_124) );
INVx1_ASAP7_75t_L g478 ( .A(n_125), .Y(n_478) );
XOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
INVx2_ASAP7_75t_L g503 ( .A(n_129), .Y(n_503) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_371), .Y(n_129) );
NAND4xp25_ASAP7_75t_L g130 ( .A(n_131), .B(n_295), .C(n_326), .D(n_355), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_262), .Y(n_131) );
OAI322xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_198), .A3(n_227), .B1(n_240), .B2(n_248), .C1(n_257), .C2(n_259), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_134), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
AND2x2_ASAP7_75t_L g292 ( .A(n_135), .B(n_293), .Y(n_292) );
INVx4_ASAP7_75t_L g328 ( .A(n_135), .Y(n_328) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g303 ( .A(n_136), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g306 ( .A(n_136), .B(n_200), .Y(n_306) );
AND2x2_ASAP7_75t_L g323 ( .A(n_136), .B(n_216), .Y(n_323) );
AND2x2_ASAP7_75t_L g421 ( .A(n_136), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g244 ( .A(n_137), .Y(n_244) );
AND2x4_ASAP7_75t_L g427 ( .A(n_137), .B(n_422), .Y(n_427) );
AO31x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_143), .A3(n_159), .B(n_165), .Y(n_137) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_138), .A2(n_211), .A3(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_139), .A2(n_590), .B(n_593), .Y(n_589) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AO31x2_ASAP7_75t_L g188 ( .A1(n_140), .A2(n_189), .A3(n_195), .B(n_196), .Y(n_188) );
AO31x2_ASAP7_75t_L g201 ( .A1(n_140), .A2(n_202), .A3(n_211), .B(n_213), .Y(n_201) );
AO31x2_ASAP7_75t_L g216 ( .A1(n_140), .A2(n_217), .A3(n_224), .B(n_225), .Y(n_216) );
AO31x2_ASAP7_75t_L g625 ( .A1(n_140), .A2(n_167), .A3(n_626), .B(n_629), .Y(n_625) );
BUFx10_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
BUFx10_ASAP7_75t_L g517 ( .A(n_141), .Y(n_517) );
INVx1_ASAP7_75t_L g541 ( .A(n_141), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_150), .B1(n_153), .B2(n_156), .Y(n_143) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_146), .Y(n_585) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g149 ( .A(n_147), .Y(n_149) );
INVx3_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
INVx1_ASAP7_75t_L g206 ( .A(n_147), .Y(n_206) );
INVx1_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
INVx2_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
INVx1_ASAP7_75t_L g235 ( .A(n_147), .Y(n_235) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_149), .B(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_179), .B(n_182), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_150), .A2(n_156), .B1(n_190), .B2(n_192), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_150), .A2(n_203), .B1(n_208), .B2(n_209), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_150), .A2(n_156), .B1(n_218), .B2(n_221), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_150), .A2(n_231), .B1(n_234), .B2(n_236), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_150), .A2(n_209), .B1(n_253), .B2(n_254), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_150), .A2(n_156), .B1(n_272), .B2(n_273), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_150), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_150), .A2(n_236), .B1(n_522), .B2(n_523), .Y(n_521) );
OAI22x1_ASAP7_75t_L g626 ( .A1(n_150), .A2(n_236), .B1(n_627), .B2(n_628), .Y(n_626) );
INVx6_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
O2A1O1Ixp5_ASAP7_75t_L g174 ( .A1(n_151), .A2(n_175), .B(n_176), .C(n_177), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_151), .A2(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_151), .B(n_584), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_151), .A2(n_580), .B(n_584), .C(n_587), .Y(n_641) );
BUFx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx1_ASAP7_75t_L g210 ( .A(n_152), .Y(n_210) );
INVx1_ASAP7_75t_L g537 ( .A(n_152), .Y(n_537) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx1_ASAP7_75t_L g207 ( .A(n_155), .Y(n_207) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g516 ( .A(n_157), .Y(n_516) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g570 ( .A(n_158), .Y(n_570) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_159), .A2(n_237), .A3(n_271), .B(n_274), .Y(n_270) );
AO21x2_ASAP7_75t_L g588 ( .A1(n_159), .A2(n_589), .B(n_597), .Y(n_588) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_161), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_161), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g167 ( .A(n_162), .Y(n_167) );
INVx2_ASAP7_75t_L g212 ( .A(n_162), .Y(n_212) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_162), .A2(n_541), .B(n_582), .Y(n_587) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_167), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g432 ( .A(n_168), .B(n_333), .Y(n_432) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g261 ( .A(n_169), .Y(n_261) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_169), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_187), .Y(n_169) );
AND2x2_ASAP7_75t_L g249 ( .A(n_170), .B(n_188), .Y(n_249) );
INVx1_ASAP7_75t_L g290 ( .A(n_170), .Y(n_290) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_185), .Y(n_170) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_171), .A2(n_173), .B(n_185), .Y(n_285) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_172), .B(n_197), .Y(n_196) );
BUFx3_ASAP7_75t_L g224 ( .A(n_172), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_172), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_172), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g554 ( .A(n_172), .B(n_517), .Y(n_554) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_178), .B(n_183), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_176), .A2(n_567), .B(n_568), .C(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g193 ( .A(n_181), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_181), .A2(n_223), .B1(n_595), .B2(n_596), .Y(n_594) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_SL g237 ( .A(n_184), .Y(n_237) );
INVx2_ASAP7_75t_L g195 ( .A(n_186), .Y(n_195) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_186), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
AND2x2_ASAP7_75t_L g345 ( .A(n_187), .B(n_284), .Y(n_345) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g299 ( .A(n_188), .Y(n_299) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_188), .Y(n_352) );
OR2x2_ASAP7_75t_L g423 ( .A(n_188), .B(n_229), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_191), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g524 ( .A(n_194), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_194), .B(n_549), .Y(n_548) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_195), .A2(n_513), .A3(n_517), .B(n_518), .Y(n_512) );
NAND4xp25_ASAP7_75t_L g301 ( .A(n_198), .B(n_302), .C(n_305), .D(n_307), .Y(n_301) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g439 ( .A(n_199), .B(n_427), .Y(n_439) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_215), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_200), .B(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g293 ( .A(n_200), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g313 ( .A(n_200), .Y(n_313) );
INVx1_ASAP7_75t_L g330 ( .A(n_200), .Y(n_330) );
INVx1_ASAP7_75t_L g338 ( .A(n_200), .Y(n_338) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_200), .Y(n_452) );
INVx4_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_201), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g370 ( .A(n_201), .B(n_270), .Y(n_370) );
AND2x2_ASAP7_75t_L g378 ( .A(n_201), .B(n_216), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_201), .B(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g443 ( .A(n_201), .Y(n_443) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_206), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g236 ( .A(n_210), .Y(n_236) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_211), .A2(n_237), .A3(n_521), .B(n_525), .Y(n_520) );
AOI21x1_ASAP7_75t_L g529 ( .A1(n_211), .A2(n_530), .B(n_542), .Y(n_529) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_212), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_212), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g598 ( .A(n_212), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_212), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g247 ( .A(n_216), .Y(n_247) );
OR2x2_ASAP7_75t_L g308 ( .A(n_216), .B(n_270), .Y(n_308) );
INVx2_ASAP7_75t_L g315 ( .A(n_216), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_216), .B(n_268), .Y(n_339) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_216), .Y(n_426) );
OAI21xp33_ASAP7_75t_SL g546 ( .A1(n_219), .A2(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AO31x2_ASAP7_75t_L g229 ( .A1(n_224), .A2(n_230), .A3(n_237), .B(n_238), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_227), .B(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g250 ( .A(n_229), .B(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g260 ( .A(n_229), .Y(n_260) );
INVx2_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
AND2x4_ASAP7_75t_L g310 ( .A(n_229), .B(n_282), .Y(n_310) );
OR2x2_ASAP7_75t_L g390 ( .A(n_229), .B(n_290), .Y(n_390) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_233), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_236), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_245), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_242), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g307 ( .A(n_242), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_242), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_243), .B(n_313), .Y(n_321) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
OR2x2_ASAP7_75t_L g359 ( .A(n_244), .B(n_269), .Y(n_359) );
INVx1_ASAP7_75t_L g286 ( .A(n_245), .Y(n_286) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g258 ( .A(n_246), .Y(n_258) );
INVx1_ASAP7_75t_L g294 ( .A(n_247), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
OAI322xp33_ASAP7_75t_L g262 ( .A1(n_249), .A2(n_263), .A3(n_276), .B1(n_279), .B2(n_286), .C1(n_287), .C2(n_291), .Y(n_262) );
AND2x4_ASAP7_75t_L g309 ( .A(n_249), .B(n_310), .Y(n_309) );
AOI211xp5_ASAP7_75t_SL g340 ( .A1(n_249), .A2(n_341), .B(n_342), .C(n_346), .Y(n_340) );
AND2x2_ASAP7_75t_L g360 ( .A(n_249), .B(n_250), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_249), .B(n_277), .Y(n_366) );
AND2x4_ASAP7_75t_SL g288 ( .A(n_250), .B(n_289), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_250), .B(n_306), .C(n_334), .Y(n_379) );
AND2x2_ASAP7_75t_L g410 ( .A(n_250), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g277 ( .A(n_251), .B(n_278), .Y(n_277) );
INVx3_ASAP7_75t_L g282 ( .A(n_251), .Y(n_282) );
BUFx2_ASAP7_75t_L g350 ( .A(n_251), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_260), .B(n_284), .Y(n_283) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_260), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_261), .B(n_277), .Y(n_408) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g351 ( .A(n_266), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_270), .Y(n_304) );
AND2x4_ASAP7_75t_L g314 ( .A(n_270), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g401 ( .A(n_270), .Y(n_401) );
INVx2_ASAP7_75t_L g422 ( .A(n_270), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_276), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g346 ( .A(n_277), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g300 ( .A(n_278), .B(n_284), .Y(n_300) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x4_ASAP7_75t_L g289 ( .A(n_281), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g411 ( .A(n_281), .Y(n_411) );
INVx2_ASAP7_75t_L g297 ( .A(n_282), .Y(n_297) );
AND2x2_ASAP7_75t_L g325 ( .A(n_282), .B(n_284), .Y(n_325) );
INVx3_ASAP7_75t_L g333 ( .A(n_282), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_282), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g318 ( .A(n_283), .Y(n_318) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
OAI222xp33_ASAP7_75t_L g457 ( .A1(n_287), .A2(n_447), .B1(n_458), .B2(n_461), .C1(n_463), .C2(n_465), .Y(n_457) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g398 ( .A(n_289), .Y(n_398) );
AND2x2_ASAP7_75t_L g462 ( .A(n_289), .B(n_332), .Y(n_462) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_292), .B(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_301), .B1(n_309), .B2(n_311), .C(n_316), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g384 ( .A(n_297), .Y(n_384) );
INVx2_ASAP7_75t_L g446 ( .A(n_298), .Y(n_446) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g347 ( .A(n_299), .Y(n_347) );
AND2x2_ASAP7_75t_L g383 ( .A(n_299), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g349 ( .A(n_300), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g375 ( .A(n_300), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g464 ( .A(n_300), .Y(n_464) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g413 ( .A(n_304), .Y(n_413) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g436 ( .A(n_306), .B(n_314), .Y(n_436) );
AND2x2_ASAP7_75t_L g459 ( .A(n_306), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g320 ( .A(n_308), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g455 ( .A(n_308), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_309), .A2(n_363), .B1(n_397), .B2(n_399), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_309), .A2(n_425), .B(n_428), .Y(n_424) );
INVxp67_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
INVx2_ASAP7_75t_SL g445 ( .A(n_310), .Y(n_445) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
OR2x2_ASAP7_75t_L g358 ( .A(n_312), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g456 ( .A(n_312), .B(n_455), .Y(n_456) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g329 ( .A(n_314), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_314), .B(n_338), .Y(n_354) );
INVx2_ASAP7_75t_L g381 ( .A(n_314), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B1(n_322), .B2(n_324), .Y(n_316) );
NOR2xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_318), .A2(n_392), .B1(n_405), .B2(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g414 ( .A(n_323), .B(n_415), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_331), .B(n_335), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g395 ( .A(n_328), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_328), .B(n_378), .Y(n_406) );
INVx1_ASAP7_75t_L g364 ( .A(n_330), .Y(n_364) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_332), .B(n_345), .Y(n_437) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g450 ( .A1(n_333), .A2(n_451), .B(n_453), .Y(n_450) );
OAI21xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_340), .B(n_348), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
INVx1_ASAP7_75t_L g460 ( .A(n_339), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g433 ( .A(n_343), .Y(n_433) );
OR2x2_ASAP7_75t_L g444 ( .A(n_344), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .C(n_353), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_349), .A2(n_410), .B1(n_412), .B2(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g376 ( .A(n_350), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_351), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_354), .B(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_354), .A2(n_417), .B1(n_420), .B2(n_423), .C(n_424), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B(n_361), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g365 ( .A(n_359), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B1(n_367), .B2(n_848), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g448 ( .A(n_370), .B(n_426), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g371 ( .A(n_372), .B(n_402), .C(n_429), .D(n_449), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_385), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_379), .B2(n_380), .C(n_382), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_375), .A2(n_432), .B1(n_454), .B2(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g412 ( .A(n_378), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_378), .B(n_421), .Y(n_420) );
NAND2x1_ASAP7_75t_L g465 ( .A(n_378), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_380), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g387 ( .A(n_384), .B(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_391), .B(n_396), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g429 ( .A1(n_401), .A2(n_430), .B(n_434), .C(n_440), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_416), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_404), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g463 ( .A(n_411), .B(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx3_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp33_ASAP7_75t_R g440 ( .A1(n_441), .A2(n_444), .B1(n_446), .B2(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g454 ( .A(n_443), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_457), .Y(n_449) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx5_ASAP7_75t_L g477 ( .A(n_470), .Y(n_477) );
INVx5_ASAP7_75t_L g482 ( .A(n_470), .Y(n_482) );
AND2x6_ASAP7_75t_SL g470 ( .A(n_471), .B(n_473), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_473), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2x1_ASAP7_75t_L g842 ( .A(n_474), .B(n_496), .Y(n_842) );
BUFx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx8_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g493 ( .A(n_487), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_487), .B(n_840), .Y(n_839) );
OAI321xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_497), .A3(n_828), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_490), .B(n_828), .Y(n_834) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx6_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x6_ASAP7_75t_SL g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g833 ( .A(n_497), .Y(n_833) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_501), .Y(n_504) );
BUFx8_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g841 ( .A(n_502), .B(n_842), .Y(n_841) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_720), .Y(n_505) );
NOR2xp67_ASAP7_75t_L g506 ( .A(n_507), .B(n_662), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g507 ( .A(n_508), .B(n_599), .C(n_644), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_555), .B(n_576), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_509), .A2(n_600), .B1(n_619), .B2(n_631), .Y(n_599) );
AOI22x1_ASAP7_75t_L g724 ( .A1(n_509), .A2(n_725), .B1(n_729), .B2(n_730), .Y(n_724) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_527), .Y(n_510) );
OR2x2_ASAP7_75t_L g685 ( .A(n_511), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .Y(n_511) );
OR2x2_ASAP7_75t_L g560 ( .A(n_512), .B(n_520), .Y(n_560) );
AND2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g611 ( .A(n_512), .Y(n_611) );
BUFx2_ASAP7_75t_L g661 ( .A(n_512), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_516), .A2(n_552), .B(n_553), .Y(n_551) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_516), .A2(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
AND2x2_ASAP7_75t_L g606 ( .A(n_520), .B(n_543), .Y(n_606) );
INVx1_ASAP7_75t_L g613 ( .A(n_520), .Y(n_613) );
INVx1_ASAP7_75t_L g618 ( .A(n_520), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_520), .B(n_611), .Y(n_680) );
INVx1_ASAP7_75t_L g701 ( .A(n_520), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_520), .B(n_604), .Y(n_771) );
INVx1_ASAP7_75t_L g664 ( .A(n_527), .Y(n_664) );
OR2x2_ASAP7_75t_L g716 ( .A(n_527), .B(n_680), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_543), .Y(n_527) );
AND2x2_ASAP7_75t_L g561 ( .A(n_528), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g609 ( .A(n_528), .B(n_610), .Y(n_609) );
INVxp67_ASAP7_75t_L g615 ( .A(n_528), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_528), .B(n_558), .Y(n_692) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g604 ( .A(n_529), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_538), .B(n_541), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_534), .B(n_536), .Y(n_531) );
BUFx4f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_537), .B(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g558 ( .A(n_543), .Y(n_558) );
INVx1_ASAP7_75t_L g658 ( .A(n_543), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_543), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g678 ( .A(n_543), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g700 ( .A(n_543), .B(n_701), .Y(n_700) );
NAND2x1p5_ASAP7_75t_SL g711 ( .A(n_543), .B(n_687), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_543), .B(n_618), .Y(n_801) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_551), .B(n_554), .Y(n_545) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_561), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_556), .A2(n_740), .B1(n_741), .B2(n_743), .Y(n_739) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_557), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_557), .B(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g818 ( .A(n_557), .B(n_676), .Y(n_818) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g617 ( .A(n_558), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_558), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g706 ( .A(n_558), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g657 ( .A(n_559), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g747 ( .A(n_560), .Y(n_747) );
OR2x2_ASAP7_75t_L g821 ( .A(n_560), .B(n_748), .Y(n_821) );
INVx1_ASAP7_75t_L g652 ( .A(n_561), .Y(n_652) );
INVx3_ASAP7_75t_L g656 ( .A(n_562), .Y(n_656) );
BUFx2_ASAP7_75t_L g667 ( .A(n_562), .Y(n_667) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g637 ( .A(n_563), .B(n_588), .Y(n_637) );
INVx2_ASAP7_75t_L g683 ( .A(n_563), .Y(n_683) );
INVx1_ASAP7_75t_L g715 ( .A(n_563), .Y(n_715) );
AND2x2_ASAP7_75t_L g728 ( .A(n_563), .B(n_625), .Y(n_728) );
AND2x2_ASAP7_75t_L g750 ( .A(n_563), .B(n_649), .Y(n_750) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
OAI21x1_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_571), .B(n_574), .Y(n_565) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g741 ( .A(n_577), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_577), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g766 ( .A(n_577), .B(n_634), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_577), .B(n_768), .Y(n_767) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_588), .Y(n_577) );
INVx2_ASAP7_75t_L g623 ( .A(n_578), .Y(n_623) );
AND2x2_ASAP7_75t_L g650 ( .A(n_578), .B(n_651), .Y(n_650) );
AOI21x1_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_586), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g643 ( .A(n_588), .Y(n_643) );
INVx2_ASAP7_75t_L g651 ( .A(n_588), .Y(n_651) );
OR2x2_ASAP7_75t_L g671 ( .A(n_588), .B(n_625), .Y(n_671) );
AND2x2_ASAP7_75t_L g682 ( .A(n_588), .B(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B1(n_607), .B2(n_612), .C(n_614), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI32xp33_ASAP7_75t_L g712 ( .A1(n_602), .A2(n_616), .A3(n_713), .B1(n_716), .B2(n_717), .Y(n_712) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g702 ( .A(n_603), .Y(n_702) );
AND2x2_ASAP7_75t_L g738 ( .A(n_603), .B(n_617), .Y(n_738) );
INVx1_ASAP7_75t_L g802 ( .A(n_603), .Y(n_802) );
OR2x2_ASAP7_75t_L g676 ( .A(n_604), .B(n_611), .Y(n_676) );
INVx2_ASAP7_75t_L g687 ( .A(n_604), .Y(n_687) );
BUFx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g826 ( .A(n_606), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g813 ( .A(n_609), .Y(n_813) );
INVx1_ASAP7_75t_L g827 ( .A(n_609), .Y(n_827) );
OR2x2_ASAP7_75t_L g707 ( .A(n_610), .B(n_687), .Y(n_707) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_612), .B(n_707), .Y(n_729) );
INVx1_ASAP7_75t_L g760 ( .A(n_612), .Y(n_760) );
BUFx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g794 ( .A(n_613), .Y(n_794) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2x1_ASAP7_75t_L g763 ( .A(n_615), .B(n_764), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g785 ( .A1(n_616), .A2(n_786), .B(n_791), .Y(n_785) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
AND2x2_ASAP7_75t_L g695 ( .A(n_621), .B(n_637), .Y(n_695) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_621), .Y(n_825) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g727 ( .A(n_622), .Y(n_727) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g709 ( .A(n_623), .B(n_683), .Y(n_709) );
AND2x2_ASAP7_75t_L g780 ( .A(n_623), .B(n_651), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_624), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g708 ( .A(n_624), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g787 ( .A(n_624), .B(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g636 ( .A(n_625), .Y(n_636) );
INVx2_ASAP7_75t_L g649 ( .A(n_625), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_625), .B(n_640), .Y(n_697) );
AND2x2_ASAP7_75t_L g757 ( .A(n_625), .B(n_651), .Y(n_757) );
NAND2xp33_ASAP7_75t_SL g631 ( .A(n_632), .B(n_638), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g732 ( .A(n_635), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_635), .B(n_715), .Y(n_807) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g639 ( .A(n_636), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g768 ( .A(n_636), .B(n_683), .Y(n_768) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
OR2x2_ASAP7_75t_L g713 ( .A(n_639), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g670 ( .A(n_640), .Y(n_670) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g696 ( .A(n_643), .B(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_652), .B(n_653), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g659 ( .A(n_647), .B(n_656), .Y(n_659) );
BUFx2_ASAP7_75t_L g677 ( .A(n_647), .Y(n_677) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g688 ( .A(n_648), .Y(n_688) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g703 ( .A(n_650), .B(n_667), .Y(n_703) );
INVx2_ASAP7_75t_L g719 ( .A(n_650), .Y(n_719) );
AND2x2_ASAP7_75t_L g761 ( .A(n_650), .B(n_683), .Y(n_761) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g736 ( .A(n_656), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g783 ( .A(n_657), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g814 ( .A(n_658), .Y(n_814) );
INVx2_ASAP7_75t_L g753 ( .A(n_661), .Y(n_753) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_672), .C(n_689), .D(n_704), .Y(n_662) );
NAND2xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_665), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_665), .A2(n_743), .B1(n_759), .B2(n_761), .C(n_762), .Y(n_758) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g740 ( .A(n_669), .Y(n_740) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_L g733 ( .A(n_670), .Y(n_733) );
INVx2_ASAP7_75t_L g805 ( .A(n_671), .Y(n_805) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_677), .B1(n_678), .B2(n_681), .C1(n_684), .C2(n_688), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g759 ( .A(n_675), .B(n_760), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_675), .A2(n_787), .B(n_789), .Y(n_786) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g798 ( .A(n_676), .B(n_742), .Y(n_798) );
OAI21xp33_ASAP7_75t_SL g772 ( .A1(n_677), .A2(n_698), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g691 ( .A(n_680), .B(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_680), .Y(n_743) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g742 ( .A(n_683), .Y(n_742) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g748 ( .A(n_687), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_693), .B1(n_698), .B2(n_703), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_695), .A2(n_705), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_704) );
INVx3_ASAP7_75t_R g819 ( .A(n_696), .Y(n_819) );
INVx1_ASAP7_75t_L g737 ( .A(n_697), .Y(n_737) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_700), .Y(n_754) );
INVx1_ASAP7_75t_L g764 ( .A(n_700), .Y(n_764) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_709), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g782 ( .A(n_709), .Y(n_782) );
AND2x2_ASAP7_75t_L g810 ( .A(n_709), .B(n_757), .Y(n_810) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g804 ( .A(n_714), .B(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_776), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_758), .C(n_772), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_734), .C(n_744), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI21xp33_ASAP7_75t_L g735 ( .A1(n_725), .A2(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g775 ( .A(n_727), .Y(n_775) );
AND2x2_ASAP7_75t_L g816 ( .A(n_727), .B(n_805), .Y(n_816) );
NAND2x1_ASAP7_75t_L g774 ( .A(n_728), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g796 ( .A(n_733), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_739), .Y(n_734) );
INVx1_ASAP7_75t_L g788 ( .A(n_742), .Y(n_788) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_749), .B1(n_751), .B2(n_755), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g784 ( .A(n_748), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_750), .B(n_780), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g823 ( .A(n_756), .Y(n_823) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI22xp33_ASAP7_75t_SL g762 ( .A1(n_763), .A2(n_765), .B1(n_767), .B2(n_769), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_803), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_781), .B(n_783), .C(n_785), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI21xp33_ASAP7_75t_L g792 ( .A1(n_779), .A2(n_793), .B(n_795), .Y(n_792) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
O2A1O1Ixp5_ASAP7_75t_SL g803 ( .A1(n_783), .A2(n_804), .B(n_806), .C(n_808), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_787), .A2(n_792), .B1(n_797), .B2(n_799), .Y(n_791) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_811), .B(n_815), .C(n_822), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OAI21xp5_ASAP7_75t_SL g822 ( .A1(n_823), .A2(n_824), .B(n_826), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
BUFx10_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_R g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx5_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
endmodule