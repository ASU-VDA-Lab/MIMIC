module fake_aes_2492_n_19 (n_1, n_2, n_4, n_3, n_5, n_0, n_19);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_19;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g6 ( .A(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_1), .B(n_0), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
BUFx3_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
CKINVDCx11_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
OAI21x1_ASAP7_75t_L g13 ( .A1(n_8), .A2(n_0), .B(n_1), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_11), .B(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
AOI22xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_12), .B1(n_15), .B2(n_9), .Y(n_17) );
NAND4xp25_ASAP7_75t_L g18 ( .A(n_17), .B(n_14), .C(n_9), .D(n_11), .Y(n_18) );
AOI222xp33_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_2), .B1(n_6), .B2(n_13), .C1(n_14), .C2(n_10), .Y(n_19) );
endmodule