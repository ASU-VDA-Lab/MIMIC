module real_aes_7663_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g413 ( .A(n_0), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_1), .A2(n_121), .B(n_126), .C(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g233 ( .A(n_2), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_3), .A2(n_116), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_4), .B(n_193), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_5), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g194 ( .A1(n_6), .A2(n_116), .B(n_195), .Y(n_194) );
AND2x6_ASAP7_75t_L g121 ( .A(n_7), .B(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_8), .A2(n_115), .B(n_123), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_9), .B(n_40), .Y(n_414) );
INVx1_ASAP7_75t_L g531 ( .A(n_10), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_11), .B(n_165), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_12), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g200 ( .A(n_13), .Y(n_200) );
INVx1_ASAP7_75t_L g113 ( .A(n_14), .Y(n_113) );
INVx1_ASAP7_75t_L g133 ( .A(n_15), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_16), .A2(n_134), .B(n_148), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_17), .B(n_193), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_18), .B(n_150), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_19), .B(n_116), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_20), .B(n_455), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_21), .A2(n_181), .B(n_207), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_22), .B(n_193), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_23), .B(n_165), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_24), .A2(n_130), .B(n_132), .C(n_134), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_25), .B(n_165), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_26), .Y(n_459) );
INVx1_ASAP7_75t_L g427 ( .A(n_27), .Y(n_427) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_28), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_29), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_30), .B(n_165), .Y(n_234) );
INVx1_ASAP7_75t_L g452 ( .A(n_31), .Y(n_452) );
INVx1_ASAP7_75t_L g212 ( .A(n_32), .Y(n_212) );
INVx2_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_34), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_35), .A2(n_181), .B(n_201), .C(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g453 ( .A(n_36), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_37), .A2(n_121), .B(n_126), .C(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_38), .A2(n_126), .B(n_426), .C(n_431), .Y(n_425) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_39), .Y(n_438) );
INVx1_ASAP7_75t_L g210 ( .A(n_41), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_42), .A2(n_152), .B(n_198), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_43), .B(n_165), .Y(n_164) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_44), .A2(n_99), .B1(n_691), .B2(n_700), .C1(n_710), .C2(n_716), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_44), .A2(n_415), .B1(n_684), .B2(n_703), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_44), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_45), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_46), .Y(n_449) );
INVx1_ASAP7_75t_L g497 ( .A(n_47), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_48), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_49), .B(n_116), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_50), .A2(n_126), .B1(n_207), .B2(n_209), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_51), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_52), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_53), .A2(n_198), .B(n_199), .C(n_201), .Y(n_197) );
CKINVDCx14_ASAP7_75t_R g528 ( .A(n_54), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_55), .Y(n_169) );
INVx1_ASAP7_75t_L g196 ( .A(n_56), .Y(n_196) );
INVx1_ASAP7_75t_L g122 ( .A(n_57), .Y(n_122) );
INVx1_ASAP7_75t_L g112 ( .A(n_58), .Y(n_112) );
INVx1_ASAP7_75t_SL g441 ( .A(n_59), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_60), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_61), .B(n_193), .Y(n_501) );
INVx1_ASAP7_75t_L g462 ( .A(n_62), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_SL g220 ( .A1(n_63), .A2(n_150), .B(n_201), .C(n_221), .Y(n_220) );
INVxp67_ASAP7_75t_L g222 ( .A(n_64), .Y(n_222) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_65), .A2(n_66), .B1(n_101), .B2(n_679), .C1(n_680), .C2(n_687), .Y(n_100) );
INVx1_ASAP7_75t_L g679 ( .A(n_66), .Y(n_679) );
INVx1_ASAP7_75t_L g695 ( .A(n_67), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_68), .A2(n_116), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_69), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_70), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_71), .A2(n_116), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g160 ( .A(n_72), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_73), .A2(n_115), .B(n_448), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_74), .Y(n_424) );
INVx1_ASAP7_75t_L g489 ( .A(n_75), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_76), .A2(n_121), .B(n_126), .C(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_77), .A2(n_116), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g492 ( .A(n_78), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_79), .B(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g110 ( .A(n_80), .Y(n_110) );
INVx1_ASAP7_75t_L g481 ( .A(n_81), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_82), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_83), .A2(n_121), .B(n_126), .C(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g411 ( .A(n_84), .Y(n_411) );
OR2x2_ASAP7_75t_L g678 ( .A(n_84), .B(n_412), .Y(n_678) );
OR2x2_ASAP7_75t_L g699 ( .A(n_84), .B(n_690), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_85), .A2(n_126), .B(n_461), .C(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_86), .B(n_109), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_87), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_88), .A2(n_121), .B(n_126), .C(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_89), .Y(n_186) );
INVx1_ASAP7_75t_L g219 ( .A(n_90), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_91), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_92), .B(n_147), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_93), .B(n_138), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_94), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_95), .A2(n_116), .B(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g500 ( .A(n_96), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_97), .B(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_410), .B1(n_415), .B2(n_678), .Y(n_101) );
INVx2_ASAP7_75t_SL g681 ( .A(n_102), .Y(n_681) );
OR4x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_306), .C(n_365), .D(n_392), .Y(n_102) );
NAND3xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_248), .C(n_273), .Y(n_103) );
O2A1O1Ixp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_171), .B(n_191), .C(n_224), .Y(n_104) );
AOI211xp5_ASAP7_75t_SL g396 ( .A1(n_105), .A2(n_397), .B(n_399), .C(n_402), .Y(n_396) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_140), .Y(n_105) );
INVx1_ASAP7_75t_L g271 ( .A(n_106), .Y(n_271) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g246 ( .A(n_107), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g278 ( .A(n_107), .Y(n_278) );
AND2x2_ASAP7_75t_L g333 ( .A(n_107), .B(n_302), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_107), .B(n_189), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_107), .B(n_190), .Y(n_391) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g252 ( .A(n_108), .Y(n_252) );
AND2x2_ASAP7_75t_L g295 ( .A(n_108), .B(n_158), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_108), .B(n_190), .Y(n_313) );
OA21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_114), .B(n_137), .Y(n_108) );
INVx1_ASAP7_75t_L g170 ( .A(n_109), .Y(n_170) );
INVx2_ASAP7_75t_L g175 ( .A(n_109), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g423 ( .A1(n_109), .A2(n_161), .B(n_424), .C(n_425), .Y(n_423) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_109), .A2(n_526), .B(n_532), .Y(n_525) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x2_ASAP7_75t_L g139 ( .A(n_110), .B(n_111), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_117), .B(n_121), .Y(n_161) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
INVx1_ASAP7_75t_L g430 ( .A(n_118), .Y(n_430) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g127 ( .A(n_119), .Y(n_127) );
INVx1_ASAP7_75t_L g208 ( .A(n_119), .Y(n_208) );
INVx1_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_120), .Y(n_131) );
INVx3_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
INVx1_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_120), .Y(n_165) );
INVx4_ASAP7_75t_SL g136 ( .A(n_121), .Y(n_136) );
BUFx3_ASAP7_75t_L g431 ( .A(n_121), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B(n_129), .C(n_136), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_125), .A2(n_136), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_125), .A2(n_136), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_125), .A2(n_136), .B(n_438), .C(n_439), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_SL g448 ( .A1(n_125), .A2(n_136), .B(n_449), .C(n_450), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_125), .A2(n_136), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_125), .A2(n_136), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_125), .A2(n_136), .B(n_528), .C(n_529), .Y(n_527) );
INVx5_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
BUFx3_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_127), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_130), .B(n_133), .Y(n_132) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_130), .A2(n_147), .B1(n_452), .B2(n_453), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_130), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_130), .B(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g209 ( .A1(n_131), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_209) );
INVx2_ASAP7_75t_L g211 ( .A(n_131), .Y(n_211) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g152 ( .A(n_135), .Y(n_152) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_136), .A2(n_161), .B1(n_206), .B2(n_213), .Y(n_205) );
INVx1_ASAP7_75t_L g465 ( .A(n_136), .Y(n_465) );
INVx4_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_138), .A2(n_217), .B(n_223), .Y(n_216) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_138), .Y(n_435) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx4_ASAP7_75t_L g245 ( .A(n_140), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_140), .A2(n_301), .B(n_303), .Y(n_300) );
AND2x2_ASAP7_75t_L g381 ( .A(n_140), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_158), .Y(n_140) );
INVx1_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
AND2x2_ASAP7_75t_L g250 ( .A(n_141), .B(n_190), .Y(n_250) );
OR2x2_ASAP7_75t_L g279 ( .A(n_141), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g293 ( .A(n_141), .Y(n_293) );
INVx3_ASAP7_75t_L g302 ( .A(n_141), .Y(n_302) );
AND2x2_ASAP7_75t_L g312 ( .A(n_141), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g345 ( .A(n_141), .B(n_251), .Y(n_345) );
AND2x2_ASAP7_75t_L g369 ( .A(n_141), .B(n_325), .Y(n_369) );
OR2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_155), .Y(n_141) );
AOI21xp5_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_144), .B(n_153), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_151), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_147), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_147), .A2(n_427), .B(n_428), .C(n_429), .Y(n_426) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_148), .B(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_148), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_148), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_151), .A2(n_164), .B(n_166), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_151), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
O2A1O1Ixp5_ASAP7_75t_L g480 ( .A1(n_151), .A2(n_463), .B(n_481), .C(n_482), .Y(n_480) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g167 ( .A(n_153), .Y(n_167) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_154), .A2(n_205), .B(n_214), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_154), .B(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_154), .A2(n_229), .B(n_236), .Y(n_228) );
NOR2xp33_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx3_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_157), .B(n_433), .Y(n_432) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_157), .A2(n_458), .B(n_466), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_157), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
AND2x2_ASAP7_75t_L g405 ( .A(n_158), .B(n_247), .Y(n_405) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_167), .B(n_168), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_162), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_161), .A2(n_230), .B(n_231), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_161), .A2(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_161), .A2(n_478), .B(n_479), .Y(n_477) );
INVx4_ASAP7_75t_L g181 ( .A(n_165), .Y(n_181) );
INVx2_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx1_ASAP7_75t_L g446 ( .A(n_167), .Y(n_446) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_167), .A2(n_471), .B(n_472), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_170), .B(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_170), .B(n_237), .Y(n_236) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_170), .A2(n_477), .B(n_483), .Y(n_476) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_173), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g325 ( .A(n_173), .B(n_313), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_173), .B(n_302), .Y(n_387) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g247 ( .A(n_174), .Y(n_247) );
AND2x2_ASAP7_75t_L g251 ( .A(n_174), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g292 ( .A(n_174), .B(n_293), .Y(n_292) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_185), .Y(n_174) );
INVx1_ASAP7_75t_L g455 ( .A(n_175), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_175), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_184), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_182), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_181), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g201 ( .A(n_183), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_187), .B(n_288), .Y(n_310) );
INVx1_ASAP7_75t_L g349 ( .A(n_187), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_187), .B(n_276), .Y(n_393) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
AND2x2_ASAP7_75t_L g256 ( .A(n_188), .B(n_251), .Y(n_256) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_190), .B(n_247), .Y(n_280) );
INVx1_ASAP7_75t_L g359 ( .A(n_190), .Y(n_359) );
AOI322xp5_ASAP7_75t_L g383 ( .A1(n_191), .A2(n_298), .A3(n_358), .B1(n_384), .B2(n_386), .C1(n_388), .C2(n_390), .Y(n_383) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_192), .B(n_203), .Y(n_191) );
AND2x2_ASAP7_75t_L g238 ( .A(n_192), .B(n_216), .Y(n_238) );
INVx1_ASAP7_75t_SL g241 ( .A(n_192), .Y(n_241) );
AND2x2_ASAP7_75t_L g243 ( .A(n_192), .B(n_204), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_192), .B(n_260), .Y(n_266) );
INVx2_ASAP7_75t_L g285 ( .A(n_192), .Y(n_285) );
AND2x2_ASAP7_75t_L g298 ( .A(n_192), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g336 ( .A(n_192), .B(n_260), .Y(n_336) );
BUFx2_ASAP7_75t_L g353 ( .A(n_192), .Y(n_353) );
AND2x2_ASAP7_75t_L g367 ( .A(n_192), .B(n_227), .Y(n_367) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_202), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_203), .B(n_255), .Y(n_282) );
AND2x2_ASAP7_75t_L g409 ( .A(n_203), .B(n_285), .Y(n_409) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_216), .Y(n_203) );
OR2x2_ASAP7_75t_L g254 ( .A(n_204), .B(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g260 ( .A(n_204), .Y(n_260) );
AND2x2_ASAP7_75t_L g305 ( .A(n_204), .B(n_228), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_204), .B(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_204), .Y(n_389) );
INVx2_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g463 ( .A(n_211), .Y(n_463) );
AND2x2_ASAP7_75t_L g240 ( .A(n_216), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g262 ( .A(n_216), .Y(n_262) );
BUFx2_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
AND2x2_ASAP7_75t_L g287 ( .A(n_216), .B(n_260), .Y(n_287) );
INVx3_ASAP7_75t_L g299 ( .A(n_216), .Y(n_299) );
OR2x2_ASAP7_75t_L g309 ( .A(n_216), .B(n_260), .Y(n_309) );
AOI31xp33_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_239), .A3(n_242), .B(n_244), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_238), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_226), .B(n_261), .Y(n_272) );
OR2x2_ASAP7_75t_L g296 ( .A(n_226), .B(n_266), .Y(n_296) );
INVx1_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_227), .B(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g317 ( .A(n_227), .B(n_309), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_227), .B(n_299), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_227), .B(n_335), .Y(n_334) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_227), .B(n_298), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_227), .B(n_353), .Y(n_363) );
AND2x2_ASAP7_75t_L g375 ( .A(n_227), .B(n_260), .Y(n_375) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g255 ( .A(n_228), .Y(n_255) );
INVx1_ASAP7_75t_L g321 ( .A(n_238), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_238), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_240), .B(n_316), .Y(n_350) );
AND2x4_ASAP7_75t_L g261 ( .A(n_241), .B(n_262), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g340 ( .A(n_246), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_246), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g288 ( .A(n_247), .B(n_278), .Y(n_288) );
AND2x2_ASAP7_75t_L g382 ( .A(n_247), .B(n_252), .Y(n_382) );
INVx1_ASAP7_75t_L g407 ( .A(n_247), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_253), .B1(n_256), .B2(n_257), .C(n_263), .Y(n_248) );
CKINVDCx14_ASAP7_75t_R g269 ( .A(n_249), .Y(n_269) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_250), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_253), .B(n_304), .Y(n_323) );
INVx3_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g372 ( .A(n_254), .B(n_268), .Y(n_372) );
AND2x2_ASAP7_75t_L g286 ( .A(n_255), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g316 ( .A(n_255), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_255), .B(n_299), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g386 ( .A(n_255), .B(n_356), .C(n_387), .Y(n_386) );
AOI211xp5_ASAP7_75t_SL g319 ( .A1(n_256), .A2(n_320), .B(n_322), .C(n_330), .Y(n_319) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_258), .A2(n_309), .B1(n_310), .B2(n_311), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_259), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_259), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g401 ( .A(n_261), .B(n_375), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_269), .B1(n_270), .B2(n_272), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_267), .B(n_316), .Y(n_347) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_270), .A2(n_362), .B1(n_393), .B2(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_281), .B1(n_283), .B2(n_288), .C(n_289), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_279), .A2(n_290), .B1(n_296), .B2(n_297), .C(n_300), .Y(n_289) );
INVx1_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_SL g304 ( .A(n_285), .Y(n_304) );
OR2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_309), .Y(n_377) );
AND2x2_ASAP7_75t_L g379 ( .A(n_285), .B(n_287), .Y(n_379) );
INVx1_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
AOI21xp33_ASAP7_75t_SL g348 ( .A1(n_291), .A2(n_349), .B(n_350), .Y(n_348) );
OR2x2_ASAP7_75t_L g355 ( .A(n_291), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_292), .B(n_313), .Y(n_329) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp33_ASAP7_75t_SL g346 ( .A(n_297), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_298), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_299), .B(n_335), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_302), .A2(n_315), .B(n_317), .C(n_318), .Y(n_314) );
NAND2x1_ASAP7_75t_SL g339 ( .A(n_302), .B(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_303), .A2(n_352), .B1(n_354), .B2(n_357), .Y(n_351) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_305), .B(n_395), .Y(n_394) );
NAND5xp2_ASAP7_75t_L g306 ( .A(n_307), .B(n_319), .C(n_337), .D(n_351), .E(n_360), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_314), .Y(n_307) );
INVx1_ASAP7_75t_L g364 ( .A(n_310), .Y(n_364) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_312), .A2(n_331), .B1(n_371), .B2(n_373), .C(n_376), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_313), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_316), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_316), .B(n_382), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_326), .B2(n_328), .Y(n_322) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g404 ( .A(n_333), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B1(n_345), .B2(n_346), .C(n_348), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g388 ( .A(n_343), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g395 ( .A(n_353), .Y(n_395) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_363), .B(n_364), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_368), .B(n_370), .C(n_383), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_368), .A2(n_393), .B(n_394), .C(n_396), .Y(n_392) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_372), .B(n_374), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_380), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .B(n_408), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g683 ( .A(n_410), .Y(n_683) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
NOR2x2_ASAP7_75t_L g689 ( .A(n_411), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_412), .Y(n_690) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g684 ( .A(n_415), .Y(n_684) );
OR3x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_589), .C(n_636), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_535), .C(n_560), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_475), .B1(n_502), .B2(n_505), .C(n_513), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_443), .B(n_468), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_420), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_420), .B(n_518), .Y(n_633) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_434), .Y(n_420) );
AND2x2_ASAP7_75t_L g504 ( .A(n_421), .B(n_474), .Y(n_504) );
AND2x2_ASAP7_75t_L g553 ( .A(n_421), .B(n_473), .Y(n_553) );
AND2x2_ASAP7_75t_L g574 ( .A(n_421), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g579 ( .A(n_421), .B(n_546), .Y(n_579) );
OR2x2_ASAP7_75t_L g587 ( .A(n_421), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g659 ( .A(n_421), .B(n_456), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_421), .B(n_608), .Y(n_673) );
INVx3_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g519 ( .A(n_422), .B(n_434), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_422), .B(n_456), .Y(n_520) );
AND2x4_ASAP7_75t_L g541 ( .A(n_422), .B(n_474), .Y(n_541) );
AND2x2_ASAP7_75t_L g571 ( .A(n_422), .B(n_445), .Y(n_571) );
AND2x2_ASAP7_75t_L g580 ( .A(n_422), .B(n_570), .Y(n_580) );
AND2x2_ASAP7_75t_L g596 ( .A(n_422), .B(n_457), .Y(n_596) );
OR2x2_ASAP7_75t_L g605 ( .A(n_422), .B(n_588), .Y(n_605) );
AND2x2_ASAP7_75t_L g611 ( .A(n_422), .B(n_546), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_422), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g625 ( .A(n_422), .B(n_470), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_422), .B(n_515), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_422), .B(n_575), .Y(n_664) );
OR2x6_ASAP7_75t_L g422 ( .A(n_423), .B(n_432), .Y(n_422) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_430), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
AND2x2_ASAP7_75t_L g570 ( .A(n_434), .B(n_456), .Y(n_570) );
AND2x2_ASAP7_75t_L g575 ( .A(n_434), .B(n_457), .Y(n_575) );
INVx1_ASAP7_75t_L g631 ( .A(n_434), .Y(n_631) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_442), .Y(n_434) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_435), .A2(n_487), .B(n_493), .Y(n_486) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_435), .A2(n_495), .B(n_501), .Y(n_494) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g540 ( .A(n_444), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_456), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_445), .B(n_504), .Y(n_503) );
BUFx3_ASAP7_75t_L g518 ( .A(n_445), .Y(n_518) );
OR2x2_ASAP7_75t_L g588 ( .A(n_445), .B(n_456), .Y(n_588) );
OR2x2_ASAP7_75t_L g649 ( .A(n_445), .B(n_556), .Y(n_649) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_454), .Y(n_445) );
INVx1_ASAP7_75t_L g471 ( .A(n_447), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_454), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_456), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g608 ( .A(n_456), .B(n_470), .Y(n_608) );
INVx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g547 ( .A(n_457), .Y(n_547) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_469), .A2(n_653), .B1(n_657), .B2(n_660), .C(n_661), .Y(n_652) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
INVx1_ASAP7_75t_SL g516 ( .A(n_470), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_470), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g647 ( .A(n_470), .B(n_504), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_473), .B(n_518), .Y(n_639) );
AND2x2_ASAP7_75t_L g546 ( .A(n_474), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g550 ( .A(n_475), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_475), .B(n_556), .Y(n_586) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
AND2x2_ASAP7_75t_L g512 ( .A(n_476), .B(n_486), .Y(n_512) );
INVx4_ASAP7_75t_L g524 ( .A(n_476), .Y(n_524) );
BUFx3_ASAP7_75t_L g566 ( .A(n_476), .Y(n_566) );
AND3x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_582), .C(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_L g663 ( .A(n_485), .B(n_577), .Y(n_663) );
AND2x2_ASAP7_75t_L g671 ( .A(n_485), .B(n_556), .Y(n_671) );
INVx1_ASAP7_75t_SL g676 ( .A(n_485), .Y(n_676) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
INVx1_ASAP7_75t_SL g534 ( .A(n_486), .Y(n_534) );
AND2x2_ASAP7_75t_L g557 ( .A(n_486), .B(n_524), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_486), .B(n_508), .Y(n_559) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_486), .Y(n_599) );
OR2x2_ASAP7_75t_L g604 ( .A(n_486), .B(n_524), .Y(n_604) );
INVx2_ASAP7_75t_L g510 ( .A(n_494), .Y(n_510) );
AND2x2_ASAP7_75t_L g544 ( .A(n_494), .B(n_525), .Y(n_544) );
OR2x2_ASAP7_75t_L g564 ( .A(n_494), .B(n_525), .Y(n_564) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_494), .Y(n_584) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g634 ( .A1(n_503), .A2(n_543), .B(n_635), .Y(n_634) );
AOI322xp5_ASAP7_75t_L g670 ( .A1(n_505), .A2(n_515), .A3(n_541), .B1(n_671), .B2(n_672), .C1(n_674), .C2(n_677), .Y(n_670) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_507), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_508), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g533 ( .A(n_509), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g601 ( .A(n_510), .B(n_524), .Y(n_601) );
AND2x2_ASAP7_75t_L g668 ( .A(n_510), .B(n_525), .Y(n_668) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g609 ( .A(n_512), .B(n_563), .Y(n_609) );
AOI31xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_517), .A3(n_520), .B(n_521), .Y(n_513) );
AND2x2_ASAP7_75t_L g568 ( .A(n_515), .B(n_546), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_515), .B(n_538), .Y(n_650) );
AND2x2_ASAP7_75t_L g669 ( .A(n_515), .B(n_574), .Y(n_669) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_518), .B(n_546), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g592 ( .A(n_518), .B(n_575), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_518), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_518), .B(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_519), .B(n_575), .Y(n_607) );
INVx1_ASAP7_75t_L g651 ( .A(n_519), .Y(n_651) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_533), .Y(n_522) );
INVxp67_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_524), .B(n_534), .Y(n_539) );
INVx1_ASAP7_75t_L g645 ( .A(n_524), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_524), .B(n_622), .Y(n_656) );
BUFx3_ASAP7_75t_L g556 ( .A(n_525), .Y(n_556) );
AND2x2_ASAP7_75t_L g582 ( .A(n_525), .B(n_534), .Y(n_582) );
INVx2_ASAP7_75t_L g622 ( .A(n_525), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_533), .B(n_655), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_540), .B(n_542), .C(n_551), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_537), .A2(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_538), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_538), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g618 ( .A(n_539), .B(n_564), .Y(n_618) );
INVx3_ASAP7_75t_L g549 ( .A(n_541), .Y(n_549) );
OAI22xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_545), .B1(n_548), .B2(n_550), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_544), .A2(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_544), .B(n_557), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_544), .B(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g548 ( .A(n_547), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g617 ( .A(n_547), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g561 ( .A1(n_548), .A2(n_562), .B(n_567), .Y(n_561) );
OAI22xp33_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_554), .B1(n_558), .B2(n_559), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_553), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g577 ( .A(n_556), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_556), .B(n_599), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_572), .C(n_585), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g627 ( .A1(n_562), .A2(n_628), .B1(n_632), .B2(n_633), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g632 ( .A(n_564), .B(n_565), .Y(n_632) );
AND2x2_ASAP7_75t_L g640 ( .A(n_565), .B(n_621), .Y(n_640) );
CKINVDCx16_ASAP7_75t_R g565 ( .A(n_566), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_SL g648 ( .A1(n_566), .A2(n_649), .B(n_650), .C(n_651), .Y(n_648) );
OR2x2_ASAP7_75t_L g675 ( .A(n_566), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_576), .B(n_578), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_574), .A2(n_611), .B(n_612), .C(n_615), .Y(n_610) );
OAI21xp33_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_580), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g643 ( .A(n_582), .B(n_601), .Y(n_643) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g621 ( .A(n_584), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_586), .Y(n_626) );
NAND3xp33_ASAP7_75t_SL g589 ( .A(n_590), .B(n_610), .C(n_623), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B(n_594), .C(n_602), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g660 ( .A(n_597), .Y(n_660) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g620 ( .A(n_599), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_599), .B(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_605), .C(n_606), .Y(n_602) );
INVx2_ASAP7_75t_SL g614 ( .A(n_604), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_605), .A2(n_616), .B1(n_618), .B2(n_619), .Y(n_615) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_627), .C(n_634), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVxp33_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g677 ( .A(n_631), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_637), .B(n_652), .C(n_665), .D(n_670), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_641), .C(n_648), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B(n_646), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_642), .A2(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_649), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g686 ( .A(n_678), .Y(n_686) );
OAI22xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B1(n_684), .B2(n_685), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx3_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NAND2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_697), .Y(n_692) );
NOR2xp33_ASAP7_75t_SL g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_SL g715 ( .A(n_694), .Y(n_715) );
INVx1_ASAP7_75t_L g714 ( .A(n_696), .Y(n_714) );
OA21x2_ASAP7_75t_L g717 ( .A1(n_696), .A2(n_715), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g705 ( .A(n_699), .Y(n_705) );
INVx1_ASAP7_75t_SL g708 ( .A(n_699), .Y(n_708) );
BUFx2_ASAP7_75t_L g718 ( .A(n_699), .Y(n_718) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
endmodule