module fake_jpeg_18077_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_41),
.Y(n_43)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_27),
.Y(n_58)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_18),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_23),
.B1(n_24),
.B2(n_0),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_19),
.B1(n_13),
.B2(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_58),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_27),
.B1(n_21),
.B2(n_17),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_32),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_68),
.B(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_15),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_11),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_24),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_87),
.B1(n_77),
.B2(n_63),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_60),
.B(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_57),
.B1(n_60),
.B2(n_35),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_41),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_93),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_73),
.C(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_95),
.B1(n_33),
.B2(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_100),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_69),
.B1(n_78),
.B2(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_104),
.B1(n_105),
.B2(n_92),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_88),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_65),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_81),
.B1(n_93),
.B2(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_86),
.C(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_111),
.C(n_39),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_83),
.B(n_87),
.C(n_92),
.D(n_89),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_99),
.B(n_100),
.C(n_96),
.D(n_39),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_100),
.C(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_32),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_114),
.A2(n_95),
.B(n_33),
.C(n_46),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_32),
.C(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_120),
.B(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_4),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_123),
.C(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_37),
.Y(n_131)
);

OAI221xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_112),
.B1(n_37),
.B2(n_10),
.C(n_11),
.Y(n_128)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.C(n_47),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_130),
.B(n_47),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_1),
.B1(n_9),
.B2(n_46),
.C(n_128),
.Y(n_134)
);


endmodule