module fake_jpeg_2411_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_0),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_59),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_55),
.B1(n_46),
.B2(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_56),
.B1(n_39),
.B2(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_56),
.B1(n_52),
.B2(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_55),
.B1(n_46),
.B2(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_43),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_53),
.B(n_41),
.C(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_51),
.B1(n_49),
.B2(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_41),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_43),
.B1(n_47),
.B2(n_45),
.Y(n_74)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_63),
.B1(n_61),
.B2(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_83),
.B1(n_85),
.B2(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_81),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_59),
.B1(n_57),
.B2(n_2),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_89),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_74),
.C(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_92),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_74),
.C(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_74),
.B1(n_62),
.B2(n_63),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_99),
.B1(n_24),
.B2(n_7),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_63),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_89),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_57),
.B(n_1),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_0),
.B(n_3),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_57),
.B1(n_31),
.B2(n_30),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_29),
.C(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_80),
.B1(n_1),
.B2(n_2),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_123),
.B1(n_9),
.B2(n_11),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_117),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_80),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_120),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_106),
.C(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_130),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_105),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_136),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_6),
.B(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_22),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_12),
.B(n_13),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_141),
.B1(n_119),
.B2(n_112),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_14),
.B(n_15),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_114),
.B1(n_115),
.B2(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_150),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_129),
.B1(n_127),
.B2(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_130),
.C(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_161),
.A2(n_160),
.B(n_152),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_143),
.B1(n_161),
.B2(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_143),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_162),
.C(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_147),
.C(n_144),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_136),
.C(n_150),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_137),
.Y(n_169)
);


endmodule