module real_jpeg_26119_n_16 (n_5, n_4, n_8, n_0, n_12, n_353, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_353;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g88 ( 
.A(n_3),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_92),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_31),
.C(n_47),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_82),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_75),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_28),
.B1(n_168),
.B2(n_171),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_52),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_5),
.A2(n_52),
.B1(n_66),
.B2(n_69),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_5),
.A2(n_52),
.B1(n_81),
.B2(n_91),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_6),
.A2(n_39),
.B1(n_49),
.B2(n_50),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_6),
.A2(n_39),
.B1(n_66),
.B2(n_69),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_6),
.A2(n_39),
.B1(n_84),
.B2(n_286),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_68),
.B1(n_81),
.B2(n_91),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_68),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_9),
.A2(n_36),
.B1(n_66),
.B2(n_69),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_9),
.A2(n_36),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_10),
.A2(n_62),
.B1(n_90),
.B2(n_91),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_11),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_77),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_77),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_11),
.A2(n_77),
.B1(n_90),
.B2(n_91),
.Y(n_233)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_12),
.B(n_69),
.C(n_88),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_81),
.B1(n_84),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_66),
.B1(n_69),
.B2(n_95),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_95),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_95),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_346),
.C(n_351),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_344),
.B(n_349),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_331),
.B(n_343),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_294),
.A3(n_324),
.B1(n_329),
.B2(n_330),
.C(n_353),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_267),
.B(n_293),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_239),
.B(n_266),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_130),
.B(n_218),
.C(n_238),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_116),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_24),
.B(n_116),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_96),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_59),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_26),
.B(n_59),
.C(n_96),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_27),
.B(n_44),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_28),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_28),
.A2(n_41),
.B1(n_161),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_37),
.B(n_150),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_28),
.A2(n_150),
.B(n_175),
.Y(n_245)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_29),
.A2(n_35),
.B1(n_40),
.B2(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_29),
.B(n_38),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_29),
.A2(n_40),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_30),
.B(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_33),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_43),
.A2(n_112),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_43),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_53),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_45),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_45),
.A2(n_55),
.B1(n_143),
.B2(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_45),
.B(n_82),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_45),
.A2(n_55),
.B(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_46),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_48),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_50),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_49),
.A2(n_73),
.B(n_184),
.C(n_186),
.Y(n_183)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_50),
.B(n_138),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g186 ( 
.A(n_50),
.B(n_69),
.C(n_72),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_53),
.B(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_61),
.B(n_63),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_54),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_54),
.A2(n_141),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_54),
.A2(n_141),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_55),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_55),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.C(n_78),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_64),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_61),
.B(n_141),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_61),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_63),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_69),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_83),
.B(n_87),
.C(n_114),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_66),
.B(n_82),
.CON(n_185),
.SN(n_185)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_70),
.A2(n_75),
.B1(n_128),
.B2(n_185),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_70),
.A2(n_107),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_70),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_70),
.A2(n_75),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_70),
.A2(n_235),
.B(n_274),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_70),
.A2(n_75),
.B(n_107),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_105),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_74),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_74),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_80),
.Y(n_286)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_81),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_82),
.B(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_85),
.A2(n_92),
.B1(n_102),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_85),
.B(n_285),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_85),
.A2(n_92),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_85),
.A2(n_319),
.B(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_85),
.A2(n_92),
.B(n_256),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_94),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_86),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_92),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_92),
.B(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_108),
.B2(n_115),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_99),
.B(n_103),
.C(n_115),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_100),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_100),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_106),
.B(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_117),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_121),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_126),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_123),
.B(n_147),
.Y(n_224)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_217),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_212),
.B(n_216),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_196),
.B(n_211),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_179),
.B(n_195),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_157),
.B(n_178),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_144),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_139),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_151),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_152),
.C(n_155),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_164),
.B(n_177),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_163),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_169),
.B(n_176),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_194),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_194),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_190),
.C(n_191),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_206),
.C(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_229),
.C(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_265),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_250),
.B1(n_263),
.B2(n_264),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_264),
.C(n_265),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_249),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_245),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_244),
.A2(n_278),
.B(n_282),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_257),
.C(n_262),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_255),
.B(n_300),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_277),
.B1(n_288),
.B2(n_289),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_275),
.B(n_276),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_276),
.A2(n_296),
.B1(n_308),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_288),
.C(n_292),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_287),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_284),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_290),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_310),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_310),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_308),
.C(n_309),
.Y(n_295)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_298),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_303),
.C(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_313),
.C(n_323),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_304),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_315),
.C(n_317),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_323),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_333),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_341),
.B2(n_342),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_337),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_339),
.C(n_341),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_346),
.Y(n_350)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_348),
.B(n_350),
.Y(n_349)
);


endmodule