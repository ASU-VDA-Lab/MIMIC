module real_jpeg_32726_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g156 ( 
.A(n_0),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_0),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g447 ( 
.A(n_0),
.Y(n_447)
);

NAND2x1p5_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_R g357 ( 
.A(n_1),
.B(n_358),
.Y(n_357)
);

NAND2x1_ASAP7_75t_L g363 ( 
.A(n_1),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_1),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_1),
.B(n_456),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_1),
.B(n_268),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_1),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_1),
.B(n_355),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

NAND2x1p5_ASAP7_75t_L g62 ( 
.A(n_2),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_2),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_2),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_121),
.Y(n_190)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_2),
.B(n_204),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_3),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_3),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_3),
.B(n_396),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_3),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_3),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_3),
.B(n_489),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_556),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_4),
.B(n_557),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_5),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_6),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_6),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_6),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_6),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_6),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_6),
.B(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_6),
.B(n_503),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_9),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_9),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_9),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_10),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_10),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_193),
.Y(n_197)
);

NAND2x1_ASAP7_75t_L g207 ( 
.A(n_10),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_10),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_10),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_10),
.B(n_355),
.Y(n_362)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_11),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_13),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_155),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_14),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

NAND2x1_ASAP7_75t_SL g56 ( 
.A(n_15),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_15),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_15),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_15),
.B(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

AND2x4_ASAP7_75t_SL g158 ( 
.A(n_17),
.B(n_59),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_17),
.B(n_213),
.Y(n_212)
);

NAND2x1_ASAP7_75t_L g233 ( 
.A(n_17),
.B(n_63),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_17),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_17),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_17),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_17),
.B(n_430),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_17),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_179),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_178),
.Y(n_20)
);

INVxp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_108),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_23),
.B(n_108),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_85),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.C(n_48),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_27),
.B(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.C(n_37),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_61),
.C(n_65),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_28),
.A2(n_29),
.B1(n_65),
.B2(n_79),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_28),
.A2(n_29),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_29),
.B(n_250),
.C(n_253),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_29),
.B(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_31),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_32),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_33),
.A2(n_112),
.B1(n_113),
.B2(n_124),
.Y(n_111)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_33),
.A2(n_37),
.B1(n_124),
.B2(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_33),
.A2(n_124),
.B1(n_306),
.B2(n_387),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_34),
.Y(n_426)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_35),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_37),
.Y(n_174)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_42),
.A2(n_48),
.B1(n_49),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_47),
.Y(n_161)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_47),
.Y(n_214)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_52),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_70),
.B2(n_71),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_120),
.C(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_61),
.A2(n_62),
.B1(n_138),
.B2(n_139),
.Y(n_290)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_64),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_65),
.Y(n_296)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_66),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_68),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_81),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_74),
.B(n_218),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g286 ( 
.A1(n_74),
.A2(n_222),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_79),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_82),
.B(n_127),
.C(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_130),
.B1(n_131),
.B2(n_135),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_R g85 ( 
.A(n_86),
.B(n_102),
.C(n_105),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_86),
.B(n_103),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.C(n_97),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_91),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_92),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_94),
.B(n_154),
.C(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_94),
.A2(n_144),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_96),
.Y(n_308)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_96),
.Y(n_467)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_167),
.C(n_170),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_109),
.B(n_542),
.Y(n_541)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_141),
.C(n_145),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_110),
.B(n_535),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_125),
.C(n_136),
.Y(n_110)
);

XOR2x2_ASAP7_75t_L g325 ( 
.A(n_111),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_123),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_120),
.C(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_120),
.B(n_203),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_120),
.Y(n_435)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_123),
.B(n_290),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_123),
.A2(n_203),
.B(n_434),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_124),
.B(n_306),
.C(n_309),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_126),
.A2(n_136),
.B1(n_137),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_126),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_131),
.A2(n_132),
.B1(n_233),
.B2(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_141),
.B(n_146),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_159),
.C(n_162),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_147),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.C(n_157),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_152),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_153),
.A2(n_154),
.B1(n_190),
.B2(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_284)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_154),
.B(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_154),
.B(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_156),
.Y(n_278)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_160),
.B1(n_192),
.B2(n_197),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_159),
.B(n_192),
.Y(n_335)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_160),
.A2(n_189),
.B(n_334),
.C(n_335),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_163),
.Y(n_332)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_168),
.B(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_170),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_171),
.B(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_175),
.B(n_177),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_227),
.C(n_233),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_529),
.B(n_552),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_408),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_345),
.B(n_404),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_183),
.B(n_409),
.C(n_411),
.Y(n_408)
);

AOI22x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_291),
.B1(n_322),
.B2(n_341),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_185),
.B(n_292),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_238),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_186),
.B(n_343),
.C(n_344),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_215),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_198),
.Y(n_187)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_188),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_190),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_190),
.A2(n_236),
.B1(n_302),
.B2(n_390),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_192),
.Y(n_334)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_196),
.Y(n_402)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_198),
.B(n_215),
.C(n_340),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.C(n_210),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_202),
.B(n_203),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_203),
.B(n_435),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_207),
.A2(n_212),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_209),
.Y(n_458)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_214),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_225),
.C(n_234),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_216),
.A2(n_217),
.B1(n_225),
.B2(n_226),
.Y(n_318)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_219),
.B(n_222),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_221),
.Y(n_463)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_229),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_230),
.Y(n_505)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_281),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_258),
.C(n_263),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_240),
.B(n_258),
.C(n_263),
.Y(n_343)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_241),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.C(n_255),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_242),
.B(n_255),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.C(n_246),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_243),
.B(n_283),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_246),
.B(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_250),
.B(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_259),
.B(n_264),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.C(n_276),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_276),
.A2(n_354),
.B(n_357),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_286),
.C(n_289),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_315),
.C(n_319),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_293),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.C(n_312),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_313),
.Y(n_349)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

XOR2x2_ASAP7_75t_SL g348 ( 
.A(n_298),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_301),
.B(n_305),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_306),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_386),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_316),
.B(n_320),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_342),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_323),
.B(n_342),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_339),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_325),
.Y(n_549)
);

INVxp33_ASAP7_75t_SL g550 ( 
.A(n_328),
.Y(n_550)
);

OAI22x1_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_328)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g539 ( 
.A(n_330),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_333),
.Y(n_540)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_337),
.B(n_539),
.C(n_540),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_339),
.A2(n_548),
.B(n_551),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_372),
.B(n_403),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_346),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_370),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_370),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.C(n_367),
.Y(n_347)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_367),
.Y(n_374)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.C(n_359),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_359),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.C(n_363),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_361),
.B(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_362),
.B(n_363),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2x2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_375),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.C(n_383),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_384),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.C(n_391),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_385),
.B(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_389),
.B1(n_391),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.C(n_398),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_392),
.A2(n_393),
.B1(n_398),
.B2(n_399),
.Y(n_519)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_395),
.B(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B(n_407),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_436),
.B(n_527),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_416),
.B(n_528),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_423),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_417),
.B(n_523),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_420),
.A2(n_421),
.B1(n_423),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_427),
.C(n_433),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_424),
.A2(n_425),
.B1(n_433),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_427),
.B(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_433),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_521),
.B(n_526),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_510),
.B(n_520),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_480),
.B(n_509),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_472),
.Y(n_439)
);

OAI22xp33_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_454),
.B1(n_470),
.B2(n_471),
.Y(n_440)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

AOI221xp5_ASAP7_75t_L g509 ( 
.A1(n_441),
.A2(n_454),
.B1(n_470),
.B2(n_471),
.C(n_472),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_452),
.B2(n_453),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_442),
.B(n_453),
.C(n_471),
.Y(n_511)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_448),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_448),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

INVx8_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_451),
.Y(n_487)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_454),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_459),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_455),
.B(n_460),
.C(n_464),
.Y(n_517)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_464),
.B1(n_468),
.B2(n_469),
.Y(n_459)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_460),
.Y(n_468)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_464),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.C(n_476),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_473),
.A2(n_474),
.B1(n_492),
.B2(n_493),
.Y(n_491)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_475),
.A2(n_476),
.B1(n_477),
.B2(n_494),
.Y(n_493)
);

CKINVDCx12_ASAP7_75t_R g494 ( 
.A(n_475),
.Y(n_494)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_495),
.B(n_508),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_491),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_491),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_488),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_488),
.Y(n_497)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_501),
.B(n_507),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_498),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_506),
.Y(n_501)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_512),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_517),
.C(n_518),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_SL g526 ( 
.A(n_522),
.B(n_525),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_544),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_554),
.B(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_541),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_541),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_536),
.C(n_538),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_546),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_538),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_547),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_550),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_550),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);


endmodule