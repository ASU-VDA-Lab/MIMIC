module fake_jpeg_21259_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_28),
.B1(n_32),
.B2(n_16),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_40),
.C(n_33),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_65),
.C(n_80),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_71),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_40),
.C(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_84),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_78),
.B1(n_56),
.B2(n_42),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_82),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_39),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_39),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_39),
.B(n_40),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_39),
.B(n_47),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_40),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_34),
.B1(n_32),
.B2(n_56),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_94),
.B1(n_97),
.B2(n_102),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_31),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_103),
.C(n_101),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_83),
.B(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_19),
.B1(n_29),
.B2(n_21),
.Y(n_97)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_76),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_19),
.B1(n_29),
.B2(n_22),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_17),
.C(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_30),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_27),
.B1(n_24),
.B2(n_18),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_26),
.B1(n_23),
.B2(n_30),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_77),
.B1(n_65),
.B2(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_125),
.B2(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_77),
.B1(n_63),
.B2(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_117),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_24),
.C(n_26),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_121),
.B(n_133),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_72),
.B(n_70),
.Y(n_121)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_63),
.B1(n_76),
.B2(n_81),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_91),
.B(n_108),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_109),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_20),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_113),
.B1(n_118),
.B2(n_127),
.Y(n_151)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_94),
.B1(n_92),
.B2(n_95),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_147),
.B1(n_137),
.B2(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_92),
.B1(n_90),
.B2(n_102),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_135),
.C(n_132),
.Y(n_172)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_95),
.B1(n_99),
.B2(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_90),
.B(n_1),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_160),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_30),
.B(n_23),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_9),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_165),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_9),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_170),
.B1(n_189),
.B2(n_158),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_150),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_126),
.B1(n_128),
.B2(n_119),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_124),
.C(n_119),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_186),
.C(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_123),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_20),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_20),
.B1(n_1),
.B2(n_0),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_185),
.B1(n_169),
.B2(n_171),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_2),
.C(n_4),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_142),
.B(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_4),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_6),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_145),
.B1(n_157),
.B2(n_161),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_212),
.B(n_173),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_146),
.C(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_8),
.C(n_9),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_150),
.B1(n_151),
.B2(n_139),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_156),
.B1(n_154),
.B2(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_143),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_143),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_207),
.C(n_184),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_150),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_169),
.B1(n_190),
.B2(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_221),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_226),
.B1(n_200),
.B2(n_207),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_190),
.C(n_187),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_227),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_181),
.B1(n_186),
.B2(n_138),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_181),
.C(n_163),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_180),
.B(n_163),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_198),
.Y(n_237)
);

AO221x1_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.C(n_211),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_223),
.B1(n_226),
.B2(n_202),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_230),
.B1(n_221),
.B2(n_214),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_223),
.C(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_220),
.B(n_218),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_8),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_198),
.C(n_217),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_217),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_10),
.Y(n_261)
);

XOR2x1_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_235),
.Y(n_256)
);

OAI21x1_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_10),
.B(n_11),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_259),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_8),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_10),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_252),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_262),
.B(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_268),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_266),
.A2(n_269),
.B(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_255),
.C(n_258),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_272),
.Y(n_275)
);

OAI211xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_259),
.B(n_13),
.C(n_14),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_271),
.B(n_14),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_278),
.A2(n_275),
.B(n_273),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_12),
.B(n_15),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_12),
.B(n_15),
.Y(n_281)
);


endmodule