module real_aes_1463_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_0), .A2(n_42), .B1(n_130), .B2(n_131), .Y(n_129) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_1), .A2(n_53), .B1(n_91), .B2(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g163 ( .A(n_2), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_3), .B(n_190), .Y(n_213) );
INVx1_ASAP7_75t_L g235 ( .A(n_4), .Y(n_235) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_5), .A2(n_16), .B1(n_91), .B2(n_99), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_6), .Y(n_251) );
INVx2_ASAP7_75t_L g189 ( .A(n_7), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_8), .A2(n_68), .B1(n_118), .B2(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g223 ( .A(n_9), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_10), .A2(n_37), .B1(n_134), .B2(n_135), .Y(n_133) );
INVx1_ASAP7_75t_L g220 ( .A(n_11), .Y(n_220) );
INVx1_ASAP7_75t_SL g295 ( .A(n_12), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_13), .B(n_200), .Y(n_199) );
AOI33xp33_ASAP7_75t_L g272 ( .A1(n_14), .A2(n_38), .A3(n_180), .B1(n_195), .B2(n_273), .B3(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g244 ( .A(n_15), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_15), .A2(n_80), .B1(n_81), .B2(n_244), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g155 ( .A1(n_16), .A2(n_53), .B1(n_56), .B2(n_156), .C(n_158), .Y(n_155) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_17), .A2(n_69), .B(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_L g191 ( .A(n_17), .B(n_69), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_18), .B(n_233), .Y(n_292) );
INVx3_ASAP7_75t_L g91 ( .A(n_19), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_20), .A2(n_80), .B1(n_81), .B2(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_20), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_21), .A2(n_71), .B1(n_104), .B2(n_108), .Y(n_103) );
INVx1_ASAP7_75t_SL g92 ( .A(n_22), .Y(n_92) );
INVx1_ASAP7_75t_L g165 ( .A(n_23), .Y(n_165) );
AND2x2_ASAP7_75t_L g184 ( .A(n_23), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g209 ( .A(n_23), .B(n_163), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_24), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_25), .B(n_85), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_26), .B(n_233), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_27), .A2(n_177), .B1(n_187), .B2(n_190), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_28), .B(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_29), .A2(n_80), .B1(n_81), .B2(n_142), .Y(n_79) );
INVx1_ASAP7_75t_L g142 ( .A(n_29), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_30), .B(n_200), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_31), .A2(n_54), .B1(n_126), .B2(n_127), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_32), .B(n_211), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_33), .B(n_200), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_34), .A2(n_38), .B1(n_148), .B2(n_149), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_34), .Y(n_149) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_35), .A2(n_56), .B1(n_91), .B2(n_95), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_36), .Y(n_186) );
INVx1_ASAP7_75t_L g148 ( .A(n_38), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_39), .B(n_200), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_40), .A2(n_47), .B1(n_112), .B2(n_115), .Y(n_111) );
INVx1_ASAP7_75t_L g181 ( .A(n_41), .Y(n_181) );
INVx1_ASAP7_75t_L g202 ( .A(n_41), .Y(n_202) );
AND2x2_ASAP7_75t_L g264 ( .A(n_43), .B(n_265), .Y(n_264) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_44), .A2(n_58), .B1(n_193), .B2(n_233), .C(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_45), .B(n_233), .Y(n_287) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_48), .B(n_187), .Y(n_253) );
INVx1_ASAP7_75t_L g556 ( .A(n_48), .Y(n_556) );
AOI21xp5_ASAP7_75t_SL g283 ( .A1(n_49), .A2(n_193), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g216 ( .A(n_50), .Y(n_216) );
INVx1_ASAP7_75t_L g262 ( .A(n_51), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_52), .A2(n_193), .B(n_261), .Y(n_260) );
INVxp33_ASAP7_75t_L g160 ( .A(n_53), .Y(n_160) );
INVx1_ASAP7_75t_L g185 ( .A(n_55), .Y(n_185) );
INVx1_ASAP7_75t_L g204 ( .A(n_55), .Y(n_204) );
INVxp67_ASAP7_75t_L g159 ( .A(n_56), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_57), .B(n_233), .Y(n_275) );
AND2x2_ASAP7_75t_L g297 ( .A(n_59), .B(n_240), .Y(n_297) );
INVx1_ASAP7_75t_L g217 ( .A(n_60), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_61), .A2(n_193), .B(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_62), .A2(n_65), .B1(n_137), .B2(n_140), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_63), .A2(n_193), .B(n_198), .C(n_210), .Y(n_192) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_64), .B(n_240), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_66), .A2(n_193), .B1(n_270), .B2(n_271), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_67), .A2(n_146), .B1(n_147), .B2(n_150), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_67), .Y(n_146) );
INVx1_ASAP7_75t_L g285 ( .A(n_70), .Y(n_285) );
AND2x2_ASAP7_75t_L g276 ( .A(n_72), .B(n_240), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_73), .A2(n_242), .B(n_243), .C(n_245), .Y(n_241) );
BUFx2_ASAP7_75t_SL g157 ( .A(n_74), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g143 ( .A1(n_75), .A2(n_144), .B1(n_145), .B2(n_151), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_75), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_76), .B(n_200), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_152), .B1(n_166), .B2(n_537), .C(n_539), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_143), .Y(n_78) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_81), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_82), .Y(n_81) );
NOR2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_124), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_103), .C(n_111), .D(n_117), .Y(n_83) );
INVx4_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
INVx6_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_96), .Y(n_87) );
AND2x2_ASAP7_75t_L g115 ( .A(n_88), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g121 ( .A(n_88), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g106 ( .A(n_89), .B(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_89), .Y(n_109) );
INVx2_ASAP7_75t_L g114 ( .A(n_89), .Y(n_114) );
OAI22x1_ASAP7_75t_L g89 ( .A1(n_90), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
INVx2_ASAP7_75t_L g99 ( .A(n_91), .Y(n_99) );
INVx1_ASAP7_75t_L g102 ( .A(n_91), .Y(n_102) );
INVx2_ASAP7_75t_L g107 ( .A(n_94), .Y(n_107) );
AND2x2_ASAP7_75t_L g113 ( .A(n_94), .B(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
AND2x6_ASAP7_75t_L g126 ( .A(n_96), .B(n_113), .Y(n_126) );
AND2x2_ASAP7_75t_L g134 ( .A(n_96), .B(n_106), .Y(n_134) );
AND2x4_ASAP7_75t_L g139 ( .A(n_96), .B(n_128), .Y(n_139) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_100), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x4_ASAP7_75t_L g105 ( .A(n_98), .B(n_100), .Y(n_105) );
AND2x2_ASAP7_75t_L g110 ( .A(n_98), .B(n_101), .Y(n_110) );
INVx1_ASAP7_75t_L g120 ( .A(n_98), .Y(n_120) );
INVxp67_ASAP7_75t_L g116 ( .A(n_100), .Y(n_116) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g119 ( .A(n_101), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g112 ( .A(n_105), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g141 ( .A(n_105), .B(n_128), .Y(n_141) );
AND2x4_ASAP7_75t_L g118 ( .A(n_106), .B(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g128 ( .A(n_107), .B(n_114), .Y(n_128) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g131 ( .A(n_110), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g135 ( .A(n_110), .B(n_128), .Y(n_135) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_113), .B(n_119), .Y(n_130) );
AND2x6_ASAP7_75t_L g127 ( .A(n_119), .B(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_120), .Y(n_123) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .C(n_133), .D(n_136), .Y(n_124) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx8_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx1_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_154), .Y(n_153) );
AND3x1_ASAP7_75t_SL g154 ( .A(n_155), .B(n_161), .C(n_164), .Y(n_154) );
INVxp67_ASAP7_75t_L g546 ( .A(n_155), .Y(n_546) );
CKINVDCx8_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_161), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_161), .A2(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g179 ( .A(n_162), .B(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_SL g551 ( .A(n_162), .B(n_164), .Y(n_551) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g197 ( .A(n_163), .B(n_181), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_164), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2x1p5_ASAP7_75t_L g194 ( .A(n_165), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_471), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_394), .Y(n_169) );
NAND3xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_341), .C(n_374), .Y(n_170) );
AOI211xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_298), .B(n_307), .C(n_331), .Y(n_171) );
OAI21xp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_227), .B(n_277), .Y(n_172) );
OR2x2_ASAP7_75t_L g351 ( .A(n_173), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g506 ( .A(n_173), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_174), .A2(n_397), .B1(n_401), .B2(n_403), .Y(n_396) );
AND2x2_ASAP7_75t_L g433 ( .A(n_174), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_212), .Y(n_174) );
INVx1_ASAP7_75t_L g330 ( .A(n_175), .Y(n_330) );
AND2x4_ASAP7_75t_L g347 ( .A(n_175), .B(n_328), .Y(n_347) );
INVx2_ASAP7_75t_L g369 ( .A(n_175), .Y(n_369) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_175), .Y(n_452) );
AND2x2_ASAP7_75t_L g523 ( .A(n_175), .B(n_280), .Y(n_523) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_192), .Y(n_175) );
NOR3xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_182), .C(n_186), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g233 ( .A(n_179), .B(n_183), .Y(n_233) );
OR2x6_ASAP7_75t_L g207 ( .A(n_180), .B(n_196), .Y(n_207) );
INVxp33_ASAP7_75t_L g273 ( .A(n_180), .Y(n_273) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_180), .Y(n_554) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x4_ASAP7_75t_L g225 ( .A(n_181), .B(n_203), .Y(n_225) );
INVxp67_ASAP7_75t_L g555 ( .A(n_182), .Y(n_555) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g196 ( .A(n_185), .Y(n_196) );
AND2x6_ASAP7_75t_L g222 ( .A(n_185), .B(n_201), .Y(n_222) );
INVx4_ASAP7_75t_L g240 ( .A(n_187), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_187), .B(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_188), .Y(n_211) );
AND2x4_ASAP7_75t_L g190 ( .A(n_189), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_189), .B(n_191), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_190), .B(n_208), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_190), .A2(n_283), .B(n_287), .Y(n_282) );
INVxp67_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_197), .Y(n_193) );
INVx1_ASAP7_75t_L g274 ( .A(n_195), .Y(n_274) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_205), .B(n_208), .Y(n_198) );
INVx1_ASAP7_75t_L g218 ( .A(n_200), .Y(n_218) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_203), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_207), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_207), .A2(n_208), .B(n_235), .C(n_236), .Y(n_234) );
INVxp67_ASAP7_75t_L g242 ( .A(n_207), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_207), .A2(n_208), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g284 ( .A1(n_207), .A2(n_208), .B(n_285), .C(n_286), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_SL g294 ( .A1(n_207), .A2(n_208), .B(n_295), .C(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g270 ( .A(n_208), .Y(n_270) );
INVx5_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_210), .A2(n_268), .B(n_276), .Y(n_267) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_210), .A2(n_268), .B(n_276), .Y(n_312) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_211), .A2(n_232), .B(n_237), .Y(n_231) );
AND2x2_ASAP7_75t_L g288 ( .A(n_212), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g317 ( .A(n_212), .Y(n_317) );
INVx3_ASAP7_75t_L g328 ( .A(n_212), .Y(n_328) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_219), .B(n_226), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_218), .B(n_244), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B1(n_223), .B2(n_224), .Y(n_219) );
INVxp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVxp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_227), .A2(n_518), .B1(n_520), .B2(n_522), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_227), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_255), .Y(n_228) );
INVx3_ASAP7_75t_L g301 ( .A(n_229), .Y(n_301) );
AND2x2_ASAP7_75t_L g309 ( .A(n_229), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_229), .Y(n_339) );
NAND2x1_ASAP7_75t_SL g533 ( .A(n_229), .B(n_300), .Y(n_533) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_238), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g306 ( .A(n_231), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_231), .B(n_312), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_231), .B(n_238), .Y(n_337) );
AND2x4_ASAP7_75t_L g344 ( .A(n_231), .B(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_231), .Y(n_393) );
INVxp67_ASAP7_75t_L g400 ( .A(n_231), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_231), .Y(n_405) );
INVx1_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
INVx1_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_238), .B(n_314), .Y(n_323) );
INVx2_ASAP7_75t_L g391 ( .A(n_238), .Y(n_391) );
INVx1_ASAP7_75t_L g430 ( .A(n_238), .Y(n_430) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B1(n_246), .B2(n_247), .Y(n_239) );
INVx3_ASAP7_75t_L g247 ( .A(n_240), .Y(n_247) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_247), .A2(n_258), .B(n_264), .Y(n_257) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_247), .A2(n_258), .B(n_264), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_252), .B1(n_253), .B2(n_254), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_254), .Y(n_538) );
AND2x2_ASAP7_75t_L g360 ( .A(n_255), .B(n_337), .Y(n_360) );
AND2x2_ASAP7_75t_L g428 ( .A(n_255), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g442 ( .A(n_255), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_255), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_267), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2x1_ASAP7_75t_L g305 ( .A(n_257), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g398 ( .A(n_257), .B(n_391), .Y(n_398) );
AND2x2_ASAP7_75t_L g489 ( .A(n_257), .B(n_311), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_265), .Y(n_290) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
INVx2_ASAP7_75t_L g345 ( .A(n_267), .Y(n_345) );
AND2x2_ASAP7_75t_L g390 ( .A(n_267), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_269), .B(n_275), .Y(n_268) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_288), .Y(n_278) );
AND2x2_ASAP7_75t_L g432 ( .A(n_279), .B(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g491 ( .A(n_279), .B(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx4_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
AND2x4_ASAP7_75t_L g329 ( .A(n_280), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g364 ( .A(n_280), .B(n_289), .Y(n_364) );
INVx2_ASAP7_75t_L g413 ( .A(n_280), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_280), .B(n_387), .Y(n_462) );
AND2x2_ASAP7_75t_L g499 ( .A(n_280), .B(n_317), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_280), .B(n_382), .Y(n_507) );
OR2x6_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g340 ( .A(n_288), .B(n_329), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_288), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_288), .B(n_367), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_288), .B(n_380), .Y(n_501) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
AND2x2_ASAP7_75t_L g327 ( .A(n_289), .B(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_289), .Y(n_350) );
INVx2_ASAP7_75t_L g353 ( .A(n_289), .Y(n_353) );
INVx1_ASAP7_75t_L g386 ( .A(n_289), .Y(n_386) );
INVx1_ASAP7_75t_L g434 ( .A(n_289), .Y(n_434) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_297), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_300), .B(n_303), .Y(n_376) );
OR2x2_ASAP7_75t_L g448 ( .A(n_300), .B(n_449), .Y(n_448) );
AND4x1_ASAP7_75t_SL g494 ( .A(n_300), .B(n_476), .C(n_495), .D(n_496), .Y(n_494) );
OR2x2_ASAP7_75t_L g518 ( .A(n_301), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g355 ( .A(n_304), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_304), .B(n_313), .Y(n_505) );
AND2x2_ASAP7_75t_L g530 ( .A(n_305), .B(n_390), .Y(n_530) );
OAI32xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_315), .A3(n_320), .B1(n_322), .B2(n_325), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_310), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g503 ( .A(n_310), .B(n_457), .Y(n_503) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x2_ASAP7_75t_L g399 ( .A(n_311), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g485 ( .A(n_311), .Y(n_485) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_312), .B(n_314), .Y(n_519) );
INVx3_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_313), .B(n_441), .Y(n_514) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_314), .Y(n_373) );
AND2x2_ASAP7_75t_L g392 ( .A(n_314), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g526 ( .A(n_316), .Y(n_526) );
NAND2x1_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_317), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_320), .B(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_326), .Y(n_358) );
AND2x4_ASAP7_75t_L g380 ( .A(n_321), .B(n_330), .Y(n_380) );
AND2x4_ASAP7_75t_SL g451 ( .A(n_321), .B(n_452), .Y(n_451) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_321), .B(n_402), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_322), .A2(n_445), .B1(n_448), .B2(n_450), .Y(n_444) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_SL g464 ( .A(n_323), .Y(n_464) );
INVx2_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_327), .B(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_327), .A2(n_463), .B1(n_466), .B2(n_469), .Y(n_465) );
INVx1_ASAP7_75t_L g387 ( .A(n_328), .Y(n_387) );
AND2x2_ASAP7_75t_L g410 ( .A(n_328), .B(n_369), .Y(n_410) );
INVx2_ASAP7_75t_L g333 ( .A(n_329), .Y(n_333) );
OAI21xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_334), .B(n_338), .Y(n_331) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_335), .A2(n_407), .B1(n_411), .B2(n_412), .Y(n_406) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_336), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_336), .B(n_404), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_336), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_357), .C(n_361), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B1(n_351), .B2(n_354), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g411 ( .A(n_344), .B(n_398), .Y(n_411) );
AND2x2_ASAP7_75t_L g463 ( .A(n_344), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g480 ( .A(n_344), .B(n_430), .Y(n_480) );
AND2x2_ASAP7_75t_L g535 ( .A(n_344), .B(n_429), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx4_ASAP7_75t_L g402 ( .A(n_347), .Y(n_402) );
AND2x2_ASAP7_75t_L g412 ( .A(n_347), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
AND2x2_ASAP7_75t_L g426 ( .A(n_350), .B(n_410), .Y(n_426) );
INVx1_ASAP7_75t_L g461 ( .A(n_352), .Y(n_461) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_355), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_356), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_370), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_363), .B(n_402), .Y(n_511) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AOI21xp33_ASAP7_75t_SL g374 ( .A1(n_366), .A2(n_375), .B(n_377), .Y(n_374) );
AND2x2_ASAP7_75t_L g521 ( .A(n_366), .B(n_380), .Y(n_521) );
AND2x4_ASAP7_75t_L g384 ( .A(n_367), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_SL g418 ( .A(n_367), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_367), .B(n_434), .Y(n_500) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_383), .B(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_380), .B(n_385), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_381), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g443 ( .A(n_381), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_381), .Y(n_447) );
AND2x2_ASAP7_75t_L g531 ( .A(n_381), .B(n_499), .Y(n_531) );
AND2x2_ASAP7_75t_L g534 ( .A(n_381), .B(n_451), .Y(n_534) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_386), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g513 ( .A(n_390), .Y(n_513) );
AND2x2_ASAP7_75t_L g404 ( .A(n_391), .B(n_405), .Y(n_404) );
NAND4xp75_ASAP7_75t_L g394 ( .A(n_395), .B(n_414), .C(n_435), .D(n_453), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_406), .Y(n_395) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_398), .B(n_485), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_399), .B(n_464), .Y(n_470) );
NAND2xp5_ASAP7_75t_R g486 ( .A(n_402), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g536 ( .A(n_402), .Y(n_536) );
INVx2_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
BUFx3_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g492 ( .A(n_410), .Y(n_492) );
AND2x2_ASAP7_75t_L g446 ( .A(n_412), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g468 ( .A(n_413), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_419), .B(n_421), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_417), .B(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_418), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_420), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B1(n_427), .B2(n_431), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
OA21x2_ASAP7_75t_L g436 ( .A1(n_429), .A2(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g457 ( .A(n_429), .Y(n_457) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g488 ( .A(n_430), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g496 ( .A(n_430), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_431), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g466 ( .A(n_434), .B(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_442), .B(n_444), .Y(n_435) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g483 ( .A(n_440), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_447), .Y(n_495) );
INVx2_ASAP7_75t_SL g487 ( .A(n_451), .Y(n_487) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_465), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B1(n_460), .B2(n_463), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_508), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .C(n_493), .Y(n_472) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_486), .B1(n_488), .B2(n_490), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .C(n_504), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_501), .B(n_502), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_527), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .C(n_524), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_515), .B2(n_516), .Y(n_510) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_518), .B(n_523), .C(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI222xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_531), .B1(n_532), .B2(n_534), .C1(n_535), .C2(n_536), .Y(n_527) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
OAI222xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_547), .B2(n_549), .C1(n_552), .C2(n_556), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
endmodule