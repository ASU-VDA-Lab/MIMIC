module real_jpeg_12707_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx4_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_55),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_4),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_121),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_47),
.B1(n_49),
.B2(n_121),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_4),
.A2(n_65),
.B1(n_67),
.B2(n_121),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_7),
.A2(n_51),
.B1(n_65),
.B2(n_67),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_36),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_8),
.B(n_63),
.C(n_65),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_8),
.A2(n_47),
.B1(n_49),
.B2(n_145),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_103),
.B1(n_106),
.B2(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_8),
.B(n_43),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_12),
.A2(n_47),
.B1(n_49),
.B2(n_123),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_12),
.A2(n_65),
.B1(n_67),
.B2(n_123),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_13),
.A2(n_47),
.B1(n_49),
.B2(n_152),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_13),
.A2(n_65),
.B1(n_67),
.B2(n_152),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_14),
.A2(n_38),
.B1(n_65),
.B2(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_14),
.A2(n_38),
.B1(n_47),
.B2(n_49),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_15),
.A2(n_24),
.B1(n_47),
.B2(n_49),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_15),
.A2(n_24),
.B1(n_65),
.B2(n_67),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_15),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_75),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_72),
.Y(n_321)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_41),
.C(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_23),
.A2(n_36),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_25),
.B(n_145),
.CON(n_144),
.SN(n_144)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_25),
.B(n_32),
.C(n_34),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_28),
.A2(n_37),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_28),
.A2(n_36),
.B1(n_144),
.B2(n_151),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_28),
.A2(n_87),
.B(n_165),
.Y(n_302)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_29),
.A2(n_33),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_29),
.A2(n_33),
.B1(n_120),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_29),
.A2(n_122),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_31),
.A2(n_35),
.B(n_144),
.C(n_146),
.Y(n_143)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g215 ( 
.A(n_35),
.B(n_145),
.CON(n_215),
.SN(n_215)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_35),
.B(n_45),
.C(n_49),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_36),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_58),
.B2(n_70),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_42),
.A2(n_78),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_50),
.B(n_56),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_43),
.A2(n_56),
.B1(n_192),
.B2(n_215),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_43),
.A2(n_56),
.B1(n_80),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x4_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_54),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_44),
.A2(n_52),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_44),
.A2(n_78),
.B1(n_148),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_44),
.A2(n_78),
.B1(n_183),
.B2(n_191),
.Y(n_190)
);

OA22x2_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_46),
.A2(n_47),
.B(n_215),
.C(n_216),
.Y(n_214)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_49),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_47),
.B(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_50),
.A2(n_56),
.B(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_72),
.C(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_58),
.A2(n_70),
.B1(n_77),
.B2(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_68),
.B(n_69),
.Y(n_58)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_59),
.A2(n_68),
.B1(n_113),
.B2(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_59),
.A2(n_135),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_59),
.A2(n_69),
.B(n_172),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_59),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_59),
.A2(n_68),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_59),
.A2(n_68),
.B1(n_220),
.B2(n_245),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_SL g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_64),
.B(n_115),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_64),
.A2(n_116),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_64),
.B(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_67),
.B(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_68),
.B(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_69),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_71),
.A2(n_72),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_75),
.A2(n_76),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_77),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_81),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_311),
.B(n_328),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_291),
.B(n_310),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_175),
.B(n_290),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_153),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_99),
.B(n_153),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_126),
.C(n_136),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_100),
.B(n_126),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_117),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_118),
.C(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_102),
.B(n_112),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B(n_109),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_103),
.A2(n_106),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_103),
.A2(n_106),
.B1(n_248),
.B2(n_256),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_103),
.A2(n_131),
.B(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_104),
.A2(n_110),
.B(n_132),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_104),
.A2(n_105),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_106),
.A2(n_129),
.B(n_142),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_106),
.B(n_145),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_114),
.B(n_230),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_133),
.B2(n_134),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_134),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_136),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.C(n_149),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_138),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_149),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_174),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_166),
.B2(n_167),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_155),
.B(n_167),
.C(n_174),
.Y(n_309)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_157),
.B(n_161),
.C(n_163),
.Y(n_294)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_162),
.Y(n_307)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_168),
.A2(n_169),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_169),
.B(n_171),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_169),
.A2(n_299),
.B(n_302),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_203),
.B(n_285),
.C(n_289),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_196),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.C(n_189),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_178),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_181),
.C(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_190),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_197),
.B(n_201),
.C(n_202),
.Y(n_286)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_279),
.B(n_284),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_234),
.B(n_278),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_222),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_222),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_217),
.C(n_218),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_209),
.A2(n_210),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_218),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_223),
.B(n_228),
.C(n_232),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_272),
.B(n_277),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_262),
.B(n_271),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_251),
.B(n_261),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_246),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_257),
.B(n_260),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_276),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_309),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_309),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_297),
.C(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_303),
.B2(n_304),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B(n_308),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_314),
.C(n_319),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_308),
.A2(n_314),
.B1(n_315),
.B2(n_327),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_323),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_320),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);


endmodule