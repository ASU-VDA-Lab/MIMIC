module real_jpeg_30652_n_32 (n_17, n_232, n_8, n_0, n_233, n_21, n_2, n_229, n_226, n_29, n_10, n_31, n_9, n_12, n_235, n_24, n_6, n_230, n_231, n_28, n_236, n_234, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_228, n_30, n_227, n_16, n_15, n_13, n_225, n_32);

input n_17;
input n_232;
input n_8;
input n_0;
input n_233;
input n_21;
input n_2;
input n_229;
input n_226;
input n_29;
input n_10;
input n_31;
input n_9;
input n_12;
input n_235;
input n_24;
input n_6;
input n_230;
input n_231;
input n_28;
input n_236;
input n_234;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_228;
input n_30;
input n_227;
input n_16;
input n_15;
input n_13;
input n_225;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_150;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_60),
.B1(n_62),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_3),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_5),
.B(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_6),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_103),
.Y(n_200)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_7),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_8),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_9),
.A2(n_112),
.B(n_116),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_10),
.Y(n_223)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_156),
.A3(n_158),
.B1(n_161),
.B2(n_183),
.C1(n_185),
.C2(n_236),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_58),
.C(n_211),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_13),
.B(n_87),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_40),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_16),
.A2(n_112),
.B(n_116),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_16),
.B(n_126),
.C(n_129),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_19),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_21),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_21),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_49),
.C(n_215),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_23),
.B(n_51),
.Y(n_214)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_24),
.B(n_93),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_26),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_27),
.Y(n_192)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_29),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_29),
.B(n_163),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_30),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_30),
.B(n_167),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_47),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g216 ( 
.A(n_37),
.Y(n_216)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_42),
.Y(n_170)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_44),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.C(n_218),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_50),
.B(n_57),
.C(n_214),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_52),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_55),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_107),
.B(n_188),
.Y(n_58)
);

NAND4xp25_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.C(n_91),
.D(n_101),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_82),
.C(n_84),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_73),
.B(n_199),
.C(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_81),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_74),
.B(n_81),
.Y(n_203)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_83),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_85),
.A2(n_191),
.B(n_194),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_85),
.B(n_91),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_88),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_88),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_91),
.A2(n_205),
.B(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI221xp5_ASAP7_75t_L g189 ( 
.A1(n_92),
.A2(n_190),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_232),
.Y(n_158)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI31xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_148),
.A3(n_171),
.B(n_178),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_140),
.C(n_141),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_130),
.B(n_139),
.Y(n_109)
);

OAI221xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_118),
.B1(n_124),
.B2(n_125),
.C(n_225),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_227),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_160),
.C(n_166),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_179),
.B(n_182),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_166),
.C(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_226),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_228),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_229),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_230),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_231),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_233),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_234),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_235),
.Y(n_174)
);


endmodule