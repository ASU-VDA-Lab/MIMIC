module fake_netlist_5_720_n_1871 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1871);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1871;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_50),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_0),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_56),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_78),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_15),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_83),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_20),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_56),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_89),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_150),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_18),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_58),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_103),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_62),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_6),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_151),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_19),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_10),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_92),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_126),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_140),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_1),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_13),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_21),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_115),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_121),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_17),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_119),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_111),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_46),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_105),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_81),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_138),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_180),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_136),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_36),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_110),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_77),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_186),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_184),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_99),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_95),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_82),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_46),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_164),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_175),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_189),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_96),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_84),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_90),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_13),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_135),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_1),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_16),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_36),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_154),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_33),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_53),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_50),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_191),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_30),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_40),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_159),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_192),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_104),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_100),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_26),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_2),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_118),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_144),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_40),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_41),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_75),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_183),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_86),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_107),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_169),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_12),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_98),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_6),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_72),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_29),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_3),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_109),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_9),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_122),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_25),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_88),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_4),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_176),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_12),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_28),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_69),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_71),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_20),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_163),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_114),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_97),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_73),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_18),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_22),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_162),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_23),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_65),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_67),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_74),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_139),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_52),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_42),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_23),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_87),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_174),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_131),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_51),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_79),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_91),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_85),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_30),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_123),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_55),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_168),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_54),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_173),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_22),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_143),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_141),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_31),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_16),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_172),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_31),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_48),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_44),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_120),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_153),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_63),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_94),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_44),
.Y(n_373)
);

CKINVDCx12_ASAP7_75t_R g374 ( 
.A(n_65),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_61),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_35),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_158),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_34),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_7),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_157),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_165),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_39),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_62),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_3),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_142),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_80),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_52),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_55),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_28),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_246),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_234),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_246),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_197),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_276),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_4),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_258),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_213),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_238),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_254),
.B(n_5),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_214),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_225),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_260),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_300),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_197),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_338),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_218),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_242),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_277),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_235),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_249),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_228),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_247),
.Y(n_414)
);

BUFx8_ASAP7_75t_SL g415 ( 
.A(n_357),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_216),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_195),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_279),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_363),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_280),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_374),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_252),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_285),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_194),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_253),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_194),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_255),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_270),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_198),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_304),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_198),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_201),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_201),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_222),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_274),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_275),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_206),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_326),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_297),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_339),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_203),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_203),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_206),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_228),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_233),
.Y(n_451)
);

BUFx6f_ASAP7_75t_SL g452 ( 
.A(n_277),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_210),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_302),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_311),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_228),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_313),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_210),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_373),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_226),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_195),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_228),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_268),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_388),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_226),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_321),
.B(n_5),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_233),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_292),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_229),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_292),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_229),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_337),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_315),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_230),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_230),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_337),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_353),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_320),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_353),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_254),
.B(n_7),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_204),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_207),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_211),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_322),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_366),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_391),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_451),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_398),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_418),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_409),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_396),
.B(n_366),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_462),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_414),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_R g504 ( 
.A(n_410),
.B(n_257),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_416),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_462),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_417),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_396),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_423),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_397),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_426),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_R g515 ( 
.A(n_428),
.B(n_265),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_429),
.B(n_259),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_437),
.B(n_259),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_438),
.B(n_282),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_450),
.Y(n_519)
);

INVxp33_ASAP7_75t_SL g520 ( 
.A(n_441),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g521 ( 
.A(n_455),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_470),
.B(n_272),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_487),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_471),
.B(n_473),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_400),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_456),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_404),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_404),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_411),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_406),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_452),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_458),
.B(n_307),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_393),
.B(n_307),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_476),
.B(n_196),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_272),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_481),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_419),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_488),
.Y(n_547)
);

AND3x2_ASAP7_75t_L g548 ( 
.A(n_395),
.B(n_382),
.C(n_349),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_406),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_405),
.B(n_196),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_405),
.B(n_244),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_464),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_415),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_424),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_435),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_446),
.B(n_236),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_464),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_466),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_394),
.B(n_243),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_446),
.B(n_244),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_401),
.B(n_273),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_420),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_479),
.B(n_205),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_390),
.B(n_392),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_436),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_403),
.B(n_277),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_531),
.Y(n_569)
);

INVx6_ASAP7_75t_L g570 ( 
.A(n_538),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_534),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_500),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_515),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_557),
.B(n_483),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_493),
.B(n_248),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_518),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_510),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_536),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_563),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_493),
.B(n_399),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_493),
.B(n_440),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_510),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_557),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_519),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_500),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_512),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_542),
.B(n_484),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_560),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_522),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_519),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_516),
.B(n_278),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_541),
.B(n_248),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_565),
.A2(n_355),
.B1(n_267),
.B2(n_221),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_554),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_565),
.A2(n_355),
.B1(n_267),
.B2(n_221),
.Y(n_597)
);

HAxp5_ASAP7_75t_SL g598 ( 
.A(n_498),
.B(n_420),
.CON(n_598),
.SN(n_598)
);

NOR2x1p5_ASAP7_75t_L g599 ( 
.A(n_491),
.B(n_368),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_517),
.B(n_341),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_525),
.B(n_541),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_528),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_539),
.B(n_452),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_520),
.A2(n_281),
.B1(n_309),
.B2(n_352),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_519),
.B(n_195),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_541),
.B(n_303),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_552),
.B(n_341),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_519),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_523),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_492),
.B(n_463),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_568),
.A2(n_367),
.B1(n_305),
.B2(n_323),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_500),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_523),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_492),
.B(n_550),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_504),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_552),
.B(n_351),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_511),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_552),
.B(n_351),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_529),
.B(n_442),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_530),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_490),
.B(n_325),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_490),
.B(n_329),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_530),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_523),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_562),
.B(n_354),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_500),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_521),
.A2(n_489),
.B1(n_482),
.B2(n_480),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_523),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_562),
.A2(n_205),
.B1(n_345),
.B2(n_354),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_540),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_540),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_529),
.B(n_452),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_491),
.A2(n_469),
.B1(n_289),
.B2(n_314),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_566),
.B(n_562),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_500),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_553),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_508),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_527),
.B(n_444),
.C(n_443),
.Y(n_642)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_498),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_490),
.B(n_332),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_546),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_499),
.B(n_334),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_533),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_543),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_514),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_499),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_494),
.A2(n_283),
.B1(n_287),
.B2(n_291),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_494),
.A2(n_489),
.B1(n_482),
.B2(n_480),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_527),
.B(n_544),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_556),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_543),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_558),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_546),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_558),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_551),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_535),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_544),
.B(n_327),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_537),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_551),
.A2(n_345),
.B1(n_467),
.B2(n_465),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_558),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_549),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_495),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_495),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_497),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_497),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_496),
.B(n_195),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_555),
.B(n_445),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_501),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_502),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_502),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_506),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_506),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_555),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_567),
.B(n_346),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_567),
.B(n_347),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_538),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_538),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_448),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_496),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_503),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_503),
.B(n_195),
.Y(n_687)
);

BUFx4f_ASAP7_75t_L g688 ( 
.A(n_505),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_559),
.B(n_454),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_505),
.Y(n_690)
);

AND2x2_ASAP7_75t_SL g691 ( 
.A(n_509),
.B(n_294),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_509),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_513),
.B(n_427),
.Y(n_693)
);

INVxp33_ASAP7_75t_L g694 ( 
.A(n_564),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_513),
.A2(n_460),
.B1(n_294),
.B2(n_299),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_532),
.B(n_294),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_532),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_559),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_545),
.Y(n_699)
);

INVx6_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_547),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_547),
.B(n_212),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_507),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_500),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_542),
.B(n_199),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_531),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_557),
.Y(n_707)
);

INVx4_ASAP7_75t_SL g708 ( 
.A(n_519),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_531),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_508),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_531),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_557),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_519),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_678),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_619),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_587),
.B(n_215),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_583),
.B(n_427),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_691),
.B(n_294),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_659),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_707),
.B(n_478),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_587),
.B(n_220),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_678),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_581),
.B(n_223),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_712),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_654),
.B(n_574),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_629),
.B(n_239),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_629),
.B(n_241),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_611),
.Y(n_729)
);

O2A1O1Ixp5_ASAP7_75t_L g730 ( 
.A1(n_575),
.A2(n_263),
.B(n_245),
.C(n_251),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_610),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_575),
.A2(n_298),
.B1(n_256),
.B2(n_261),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_580),
.A2(n_262),
.B1(n_271),
.B2(n_288),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_638),
.B(n_296),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_670),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_621),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_624),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_601),
.B(n_478),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_627),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_654),
.B(n_430),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_638),
.B(n_308),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_634),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_705),
.B(n_592),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_670),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_691),
.A2(n_310),
.B1(n_318),
.B2(n_328),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_684),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_632),
.A2(n_340),
.B(n_342),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_697),
.B(n_199),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_641),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_675),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_577),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_614),
.B(n_237),
.C(n_240),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_582),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_626),
.A2(n_331),
.B(n_333),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_582),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_581),
.B(n_294),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_705),
.A2(n_477),
.B1(n_474),
.B2(n_472),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_581),
.B(n_228),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_669),
.B(n_200),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_695),
.B(n_228),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_594),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_695),
.B(n_228),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_606),
.A2(n_477),
.B1(n_474),
.B2(n_472),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_635),
.B(n_200),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_645),
.B(n_202),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_594),
.A2(n_228),
.B1(n_269),
.B2(n_358),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_702),
.A2(n_468),
.B1(n_461),
.B2(n_459),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_658),
.B(n_202),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_586),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_660),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_594),
.A2(n_358),
.B1(n_269),
.B2(n_459),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_586),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_569),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_594),
.A2(n_468),
.B1(n_461),
.B2(n_453),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_600),
.B(n_319),
.C(n_264),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_675),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_618),
.B(n_453),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_665),
.B(n_208),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_579),
.B(n_430),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_665),
.B(n_209),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_671),
.B(n_432),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_697),
.B(n_269),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_594),
.A2(n_358),
.B1(n_269),
.B2(n_434),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_571),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_651),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_600),
.B(n_209),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_603),
.A2(n_449),
.B1(n_439),
.B2(n_434),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_671),
.B(n_432),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_651),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_697),
.B(n_269),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_603),
.A2(n_449),
.B1(n_439),
.B2(n_433),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_687),
.B(n_433),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_623),
.A2(n_356),
.B(n_224),
.C(n_227),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_623),
.A2(n_358),
.B1(n_269),
.B2(n_385),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_578),
.B(n_219),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_612),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_588),
.B(n_227),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_589),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_623),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_590),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_700),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_687),
.B(n_231),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_679),
.B(n_269),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_579),
.B(n_422),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_602),
.A2(n_360),
.B1(n_348),
.B2(n_350),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_706),
.B(n_232),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_572),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_697),
.B(n_269),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_572),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_709),
.B(n_232),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_711),
.B(n_348),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_667),
.B(n_350),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_607),
.A2(n_358),
.B1(n_385),
.B2(n_306),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_667),
.B(n_356),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_650),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_607),
.A2(n_620),
.B1(n_622),
.B2(n_633),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_579),
.B(n_422),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_667),
.B(n_358),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_674),
.B(n_360),
.Y(n_820)
);

AND2x6_ASAP7_75t_SL g821 ( 
.A(n_703),
.B(n_368),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_674),
.B(n_361),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_696),
.B(n_361),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_681),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_668),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_633),
.B(n_358),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_677),
.B(n_362),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_640),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_640),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_651),
.Y(n_830)
);

NOR2x1p5_ASAP7_75t_L g831 ( 
.A(n_619),
.B(n_371),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_362),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_620),
.B(n_70),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_673),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_644),
.A2(n_365),
.B(n_369),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_696),
.B(n_365),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_680),
.B(n_358),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_625),
.B(n_369),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_676),
.B(n_370),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_681),
.B(n_372),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_676),
.B(n_372),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_652),
.A2(n_389),
.B1(n_387),
.B2(n_371),
.C(n_376),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_672),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_573),
.B(n_377),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_637),
.B(n_380),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_672),
.A2(n_380),
.B(n_386),
.C(n_266),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_646),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_700),
.B(n_306),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_688),
.B(n_386),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_701),
.B(n_284),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_576),
.B(n_286),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_572),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_576),
.B(n_290),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_576),
.B(n_343),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_649),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_686),
.B(n_306),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_701),
.B(n_344),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_SL g858 ( 
.A(n_688),
.B(n_655),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_656),
.B(n_657),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_686),
.B(n_385),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_657),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_584),
.B(n_316),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_584),
.B(n_293),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_651),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_585),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_585),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_699),
.B(n_295),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_701),
.B(n_312),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_744),
.B(n_604),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_803),
.A2(n_636),
.B(n_685),
.C(n_690),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_747),
.Y(n_871)
);

AND2x2_ASAP7_75t_SL g872 ( 
.A(n_858),
.B(n_693),
.Y(n_872)
);

OA21x2_ASAP7_75t_L g873 ( 
.A1(n_837),
.A2(n_622),
.B(n_647),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_721),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_726),
.B(n_692),
.Y(n_875)
);

OR2x6_ASAP7_75t_SL g876 ( 
.A(n_715),
.B(n_655),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_843),
.B(n_595),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_740),
.B(n_692),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_718),
.A2(n_642),
.B(n_597),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_716),
.B(n_595),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_722),
.B(n_597),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_741),
.B(n_700),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_817),
.A2(n_631),
.B1(n_653),
.B2(n_664),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_859),
.A2(n_713),
.B(n_584),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_761),
.A2(n_599),
.B1(n_689),
.B2(n_613),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_734),
.B(n_591),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_816),
.Y(n_887)
);

BUFx4f_ASAP7_75t_L g888 ( 
.A(n_848),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_800),
.B(n_682),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_750),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_803),
.A2(n_683),
.B(n_682),
.C(n_698),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_808),
.A2(n_628),
.B(n_613),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_721),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_777),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_717),
.B(n_689),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_727),
.A2(n_628),
.B(n_613),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_717),
.B(n_598),
.C(n_689),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_825),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_728),
.A2(n_628),
.B(n_609),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_746),
.A2(n_605),
.B(n_683),
.C(n_664),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_848),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_735),
.B(n_609),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_778),
.B(n_661),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_782),
.A2(n_609),
.B1(n_710),
.B2(n_663),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_735),
.A2(n_608),
.B(n_616),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_802),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_823),
.A2(n_694),
.B(n_643),
.C(n_666),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_777),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_802),
.B(n_641),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_745),
.A2(n_608),
.B(n_616),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_751),
.B(n_708),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_729),
.B(n_596),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_834),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_782),
.A2(n_570),
.B1(n_704),
.B2(n_630),
.Y(n_914)
);

AO21x2_ASAP7_75t_L g915 ( 
.A1(n_742),
.A2(n_704),
.B(n_585),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_759),
.A2(n_616),
.B(n_593),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_725),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_731),
.B(n_585),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_719),
.Y(n_919)
);

O2A1O1Ixp5_ASAP7_75t_L g920 ( 
.A1(n_757),
.A2(n_694),
.B(n_643),
.C(n_570),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_810),
.A2(n_593),
.B(n_608),
.Y(n_921)
);

INVx11_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_810),
.A2(n_593),
.B(n_608),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_848),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_810),
.A2(n_593),
.B(n_616),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_852),
.A2(n_615),
.B(n_630),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_777),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_852),
.A2(n_615),
.B(n_630),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_774),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_850),
.Y(n_930)
);

AND2x2_ASAP7_75t_SL g931 ( 
.A(n_789),
.B(n_598),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_736),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_737),
.B(n_704),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_852),
.A2(n_704),
.B(n_615),
.Y(n_934)
);

OA22x2_ASAP7_75t_L g935 ( 
.A1(n_758),
.A2(n_376),
.B1(n_378),
.B2(n_379),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_862),
.A2(n_630),
.B(n_615),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_833),
.B(n_570),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_761),
.A2(n_648),
.B(n_387),
.C(n_383),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_777),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_833),
.B(n_639),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_833),
.B(n_639),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_863),
.A2(n_639),
.B(n_301),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_719),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_763),
.A2(n_648),
.B(n_383),
.C(n_379),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_778),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_789),
.B(n_617),
.Y(n_946)
);

NOR2x1_ASAP7_75t_L g947 ( 
.A(n_831),
.B(n_617),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_857),
.B(n_617),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_739),
.B(n_639),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_752),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_823),
.A2(n_11),
.B(n_14),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_836),
.A2(n_378),
.B(n_596),
.C(n_24),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_837),
.A2(n_188),
.B(n_185),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_757),
.A2(n_182),
.B(n_170),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_826),
.A2(n_160),
.B(n_156),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_793),
.B(n_596),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_865),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_819),
.A2(n_147),
.B(n_137),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_786),
.A2(n_133),
.B(n_132),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_793),
.A2(n_11),
.B1(n_14),
.B2(n_24),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_743),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_771),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_836),
.B(n_25),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_786),
.A2(n_790),
.B(n_865),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_738),
.B(n_26),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_790),
.A2(n_129),
.B(n_108),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_763),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_866),
.A2(n_106),
.B(n_102),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_738),
.B(n_27),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_752),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_838),
.B(n_32),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_780),
.B(n_34),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_733),
.A2(n_35),
.B(n_37),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_804),
.A2(n_779),
.B(n_781),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_840),
.A2(n_37),
.B(n_38),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_714),
.B(n_38),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_724),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_754),
.B(n_39),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_754),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_830),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_723),
.B(n_41),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_820),
.A2(n_43),
.B(n_45),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_826),
.A2(n_43),
.B(n_45),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_851),
.B(n_47),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_851),
.B(n_47),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_756),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_855),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_785),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_853),
.B(n_66),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_724),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_822),
.A2(n_49),
.B(n_57),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_830),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_853),
.B(n_57),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_L g994 ( 
.A(n_776),
.B(n_58),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_783),
.A2(n_59),
.B(n_60),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_827),
.A2(n_60),
.B(n_61),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_845),
.A2(n_66),
.B(n_63),
.C(n_64),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_854),
.B(n_840),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_799),
.A2(n_64),
.B1(n_801),
.B2(n_724),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_732),
.A2(n_772),
.B1(n_784),
.B2(n_845),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_756),
.B(n_770),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_832),
.A2(n_864),
.B(n_815),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_760),
.B(n_867),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_775),
.B(n_749),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_867),
.B(n_813),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_868),
.A2(n_860),
.B1(n_856),
.B2(n_854),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_770),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_783),
.A2(n_791),
.B(n_809),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_868),
.A2(n_856),
.B1(n_860),
.B2(n_787),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_847),
.B(n_861),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_773),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_773),
.A2(n_828),
.B(n_797),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_768),
.B(n_764),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_797),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_795),
.A2(n_814),
.B1(n_788),
.B2(n_792),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_762),
.B(n_769),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_765),
.A2(n_766),
.B1(n_839),
.B2(n_841),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_828),
.B(n_829),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_796),
.B(n_807),
.Y(n_1019)
);

AO32x1_ASAP7_75t_L g1020 ( 
.A1(n_730),
.A2(n_846),
.A3(n_794),
.B1(n_805),
.B2(n_818),
.Y(n_1020)
);

BUFx12f_ASAP7_75t_L g1021 ( 
.A(n_821),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_798),
.B(n_811),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_842),
.A2(n_753),
.B(n_806),
.Y(n_1023)
);

O2A1O1Ixp5_ASAP7_75t_L g1024 ( 
.A1(n_812),
.A2(n_849),
.B(n_748),
.C(n_755),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_844),
.B(n_767),
.C(n_835),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_762),
.B(n_744),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_762),
.A2(n_587),
.B(n_744),
.C(n_803),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_762),
.A2(n_718),
.B(n_716),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_762),
.A2(n_632),
.B(n_859),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_SL g1030 ( 
.A(n_762),
.B(n_758),
.C(n_604),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_762),
.A2(n_587),
.B(n_744),
.C(n_803),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_777),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_744),
.B(n_697),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_859),
.A2(n_632),
.B(n_720),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_777),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_747),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_744),
.B(n_520),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_777),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1007),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_998),
.B(n_1003),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_906),
.B(n_1030),
.Y(n_1042)
);

AO31x2_ASAP7_75t_L g1043 ( 
.A1(n_1027),
.A2(n_1031),
.A3(n_951),
.B(n_1026),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1037),
.B(n_1005),
.Y(n_1044)
);

AOI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_869),
.A2(n_1013),
.B(n_1023),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_1015),
.A2(n_931),
.B(n_883),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_984),
.A2(n_985),
.B(n_1000),
.C(n_1006),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_1032),
.B(n_1035),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_882),
.B(n_977),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1015),
.A2(n_883),
.B(n_946),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_880),
.A2(n_881),
.B(n_1000),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_880),
.A2(n_881),
.B(n_1008),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_887),
.B(n_1036),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1002),
.A2(n_899),
.B(n_896),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1016),
.A2(n_974),
.B(n_1019),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_L g1056 ( 
.A1(n_1033),
.A2(n_902),
.B(n_884),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_890),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1022),
.B(n_930),
.Y(n_1058)
);

NOR2xp67_ASAP7_75t_SL g1059 ( 
.A(n_977),
.B(n_990),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_875),
.B(n_877),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1034),
.A2(n_941),
.B(n_940),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_956),
.A2(n_903),
.B(n_963),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_940),
.A2(n_941),
.B(n_1025),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1001),
.A2(n_892),
.B(n_900),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_SL g1065 ( 
.A1(n_1032),
.A2(n_1035),
.B(n_1038),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1001),
.A2(n_873),
.B(n_1018),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_877),
.B(n_1017),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_964),
.A2(n_934),
.B(n_926),
.Y(n_1068)
);

OA22x2_ASAP7_75t_L g1069 ( 
.A1(n_945),
.A2(n_893),
.B1(n_874),
.B2(n_972),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_928),
.A2(n_905),
.B(n_910),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_916),
.A2(n_923),
.B(n_925),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1009),
.A2(n_948),
.B1(n_1004),
.B2(n_872),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_916),
.A2(n_921),
.B(n_953),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_932),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_878),
.B(n_895),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_SL g1076 ( 
.A1(n_983),
.A2(n_995),
.B(n_958),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_965),
.A2(n_969),
.B(n_993),
.C(n_989),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_873),
.A2(n_879),
.B(n_1024),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_939),
.B(n_1038),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_879),
.A2(n_933),
.B(n_918),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_971),
.A2(n_891),
.B(n_913),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_890),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_961),
.B(n_962),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_939),
.A2(n_1038),
.B(n_977),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_938),
.A2(n_944),
.B(n_920),
.C(n_870),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_911),
.A2(n_1010),
.B(n_1007),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_SL g1087 ( 
.A1(n_939),
.A2(n_990),
.B(n_914),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_876),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_915),
.A2(n_949),
.B(n_1020),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_990),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_917),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1010),
.A2(n_992),
.B(n_987),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_919),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_949),
.A2(n_1020),
.B(n_942),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_972),
.B(n_909),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_973),
.A2(n_978),
.A3(n_997),
.B(n_960),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_929),
.B(n_904),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_943),
.A2(n_986),
.B(n_970),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_SL g1099 ( 
.A1(n_975),
.A2(n_960),
.B1(n_952),
.B2(n_976),
.C(n_967),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_978),
.A2(n_898),
.B(n_950),
.Y(n_1100)
);

AND3x4_ASAP7_75t_L g1101 ( 
.A(n_947),
.B(n_981),
.C(n_889),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_999),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_889),
.B(n_894),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_992),
.A2(n_1014),
.B(n_979),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_888),
.B(n_924),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_871),
.B(n_907),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_894),
.A2(n_927),
.B(n_908),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_871),
.B(n_935),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_SL g1109 ( 
.A1(n_982),
.A2(n_996),
.B(n_991),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_888),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_994),
.A2(n_885),
.B(n_972),
.C(n_927),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_897),
.A2(n_988),
.B1(n_981),
.B2(n_901),
.C(n_924),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1011),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_SL g1114 ( 
.A1(n_935),
.A2(n_959),
.B(n_966),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_901),
.B(n_912),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_908),
.B(n_1021),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1011),
.A2(n_980),
.B(n_954),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_957),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_968),
.A2(n_1011),
.B(n_980),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_957),
.B(n_922),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_957),
.A2(n_1012),
.B(n_936),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_998),
.B(n_744),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_875),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_906),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_L g1133 ( 
.A(n_1006),
.B(n_697),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_932),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_875),
.B(n_583),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_887),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_886),
.A2(n_1033),
.B(n_1002),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1027),
.A2(n_1031),
.B(n_1026),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1037),
.B(n_945),
.Y(n_1139)
);

BUFx12f_ASAP7_75t_L g1140 ( 
.A(n_906),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_998),
.B(n_744),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_983),
.A2(n_955),
.B(n_937),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_906),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_871),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_998),
.B(n_1037),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_998),
.B(n_744),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_998),
.B(n_744),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_998),
.B(n_744),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_932),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1027),
.A2(n_1031),
.A3(n_951),
.B(n_1026),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_SL g1156 ( 
.A1(n_963),
.A2(n_971),
.B(n_1005),
.Y(n_1156)
);

AND3x4_ASAP7_75t_L g1157 ( 
.A(n_909),
.B(n_598),
.C(n_692),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_932),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1027),
.A2(n_1031),
.B(n_1026),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_875),
.B(n_583),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_869),
.B(n_661),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1027),
.A2(n_1031),
.B(n_1026),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_998),
.B(n_1037),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_886),
.A2(n_1033),
.B(n_1002),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_L g1167 ( 
.A1(n_886),
.A2(n_1033),
.B(n_1002),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_998),
.B(n_744),
.Y(n_1168)
);

AO21x1_ASAP7_75t_L g1169 ( 
.A1(n_984),
.A2(n_985),
.B(n_963),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_985),
.B(n_1023),
.C(n_1000),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1027),
.A2(n_1031),
.A3(n_951),
.B(n_1026),
.Y(n_1171)
);

AO21x1_ASAP7_75t_L g1172 ( 
.A1(n_984),
.A2(n_985),
.B(n_963),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_917),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1026),
.A2(n_886),
.B(n_1028),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_932),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_998),
.B(n_744),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1027),
.A2(n_1031),
.A3(n_951),
.B(n_1026),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_886),
.A2(n_1033),
.B(n_1002),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1012),
.A2(n_936),
.B(n_1029),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1027),
.A2(n_1031),
.B(n_1026),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_875),
.B(n_583),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1027),
.A2(n_1031),
.A3(n_951),
.B(n_1026),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1110),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1170),
.A2(n_1047),
.B1(n_1044),
.B2(n_1150),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1135),
.B(n_1161),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1049),
.B(n_1120),
.Y(n_1191)
);

BUFx2_ASAP7_75t_R g1192 ( 
.A(n_1088),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1173),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1046),
.A2(n_1050),
.B1(n_1045),
.B2(n_1062),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1074),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1136),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1102),
.A2(n_1172),
.B1(n_1169),
.B2(n_1075),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1051),
.A2(n_1063),
.B(n_1122),
.Y(n_1198)
);

HAxp5_ASAP7_75t_L g1199 ( 
.A(n_1157),
.B(n_1057),
.CON(n_1199),
.SN(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1077),
.A2(n_1072),
.B(n_1139),
.C(n_1041),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1134),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1130),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1151),
.B(n_1152),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1063),
.A2(n_1128),
.B(n_1122),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1059),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1185),
.B(n_1126),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1048),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1091),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1168),
.B(n_1180),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1084),
.B(n_1049),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1126),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1049),
.B(n_1090),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1149),
.B(n_1165),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1147),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1067),
.A2(n_1133),
.B(n_1052),
.Y(n_1215)
);

OR2x6_ASAP7_75t_SL g1216 ( 
.A(n_1162),
.B(n_1058),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1060),
.B(n_1102),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1097),
.B(n_1053),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1140),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1146),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1082),
.B(n_1106),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1118),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1090),
.B(n_1115),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1048),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1112),
.A2(n_1069),
.B1(n_1108),
.B2(n_1042),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1055),
.A2(n_1143),
.B(n_1178),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_SL g1227 ( 
.A(n_1105),
.B(n_1111),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1069),
.B(n_1083),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1154),
.B(n_1158),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_SL g1230 ( 
.A1(n_1111),
.A2(n_1138),
.B(n_1159),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1128),
.B(n_1132),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1179),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1095),
.Y(n_1233)
);

O2A1O1Ixp5_ASAP7_75t_SL g1234 ( 
.A1(n_1081),
.A2(n_1184),
.B(n_1163),
.C(n_1156),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1112),
.B(n_1095),
.Y(n_1235)
);

CKINVDCx16_ASAP7_75t_R g1236 ( 
.A(n_1095),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1103),
.B(n_1093),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1132),
.A2(n_1178),
.B(n_1177),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1101),
.B(n_1085),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1143),
.B(n_1148),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1040),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1148),
.A2(n_1177),
.B(n_1160),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1113),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1079),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1160),
.A2(n_1176),
.B(n_1164),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_R g1246 ( 
.A(n_1100),
.B(n_1137),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1087),
.B(n_1116),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1065),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1164),
.A2(n_1176),
.B(n_1174),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1098),
.B(n_1092),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1096),
.B(n_1171),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1107),
.B(n_1119),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1096),
.B(n_1099),
.Y(n_1253)
);

O2A1O1Ixp5_ASAP7_75t_L g1254 ( 
.A1(n_1094),
.A2(n_1054),
.B(n_1166),
.C(n_1167),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1109),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1080),
.A2(n_1175),
.B(n_1061),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1064),
.A2(n_1061),
.B(n_1054),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1182),
.B(n_1080),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1096),
.B(n_1043),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1104),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1096),
.B(n_1117),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1078),
.A2(n_1066),
.B(n_1117),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1086),
.B(n_1071),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1089),
.A2(n_1078),
.B(n_1094),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1121),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1114),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1056),
.B(n_1070),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1155),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1073),
.B(n_1068),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1043),
.B(n_1181),
.Y(n_1270)
);

INVx3_ASAP7_75t_SL g1271 ( 
.A(n_1144),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1155),
.Y(n_1272)
);

AND2x2_ASAP7_75t_SL g1273 ( 
.A(n_1076),
.B(n_1043),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1043),
.B(n_1181),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1039),
.A2(n_1123),
.B(n_1125),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1186),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1127),
.A2(n_1129),
.B(n_1131),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_SL g1278 ( 
.A1(n_1171),
.A2(n_1181),
.B(n_1145),
.C(n_1153),
.Y(n_1278)
);

AND2x6_ASAP7_75t_L g1279 ( 
.A(n_1141),
.B(n_1183),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1173),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1173),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1057),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1135),
.B(n_1161),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1049),
.B(n_1120),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1046),
.A2(n_1047),
.B(n_1170),
.C(n_1045),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1044),
.B(n_701),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1136),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1049),
.B(n_1120),
.Y(n_1289)
);

INVx3_ASAP7_75t_SL g1290 ( 
.A(n_1088),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1046),
.A2(n_1047),
.B(n_1170),
.C(n_1045),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1173),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1173),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1170),
.A2(n_1077),
.B(n_1047),
.C(n_1046),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1136),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1074),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1173),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1173),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1046),
.A2(n_931),
.B1(n_1050),
.B2(n_1045),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1304)
);

INVx5_ASAP7_75t_L g1305 ( 
.A(n_1090),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1135),
.B(n_1161),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1041),
.B(n_661),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1041),
.B(n_661),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1044),
.A2(n_931),
.B1(n_897),
.B2(n_1013),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1074),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1173),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1170),
.A2(n_1047),
.B1(n_1044),
.B2(n_1124),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1041),
.B(n_661),
.Y(n_1315)
);

AND2x2_ASAP7_75t_SL g1316 ( 
.A(n_1105),
.B(n_931),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1050),
.A2(n_985),
.B(n_984),
.C(n_965),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1135),
.B(n_1161),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1173),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1124),
.B(n_1142),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1044),
.B(n_701),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1170),
.A2(n_1077),
.B(n_1047),
.C(n_1046),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1057),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1074),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1173),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1170),
.A2(n_1047),
.B1(n_1044),
.B2(n_1124),
.Y(n_1326)
);

OR2x2_ASAP7_75t_SL g1327 ( 
.A(n_1044),
.B(n_897),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1046),
.A2(n_931),
.B1(n_1050),
.B2(n_1045),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1195),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1201),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1212),
.B(n_1210),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1282),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1311),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1310),
.A2(n_1328),
.B1(n_1302),
.B2(n_1227),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1227),
.A2(n_1239),
.B1(n_1316),
.B2(n_1235),
.Y(n_1335)
);

BUFx4f_ASAP7_75t_SL g1336 ( 
.A(n_1187),
.Y(n_1336)
);

BUFx2_ASAP7_75t_R g1337 ( 
.A(n_1290),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1324),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1261),
.B(n_1250),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1275),
.A2(n_1277),
.B(n_1257),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1232),
.Y(n_1341)
);

INVxp67_ASAP7_75t_SL g1342 ( 
.A(n_1288),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1188),
.B(n_1203),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1200),
.B(n_1194),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1297),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1250),
.Y(n_1346)
);

CKINVDCx16_ASAP7_75t_R g1347 ( 
.A(n_1280),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1197),
.B(n_1188),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1296),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1189),
.A2(n_1314),
.B1(n_1326),
.B2(n_1221),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1323),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1196),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1203),
.B(n_1209),
.Y(n_1353)
);

AO21x1_ASAP7_75t_SL g1354 ( 
.A1(n_1259),
.A2(n_1268),
.B(n_1272),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1190),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1283),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1251),
.B(n_1274),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_SL g1358 ( 
.A(n_1281),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1261),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1229),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1225),
.A2(n_1327),
.B1(n_1216),
.B2(n_1217),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1210),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1292),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1255),
.B(n_1260),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1211),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1229),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1211),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1260),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1241),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1265),
.B(n_1273),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1237),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1217),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1206),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1213),
.A2(n_1218),
.B1(n_1228),
.B2(n_1306),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1210),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1189),
.A2(n_1326),
.B1(n_1314),
.B2(n_1266),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1318),
.A2(n_1247),
.B1(n_1301),
.B2(n_1320),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1212),
.B(n_1223),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1209),
.A2(n_1293),
.B1(n_1307),
.B2(n_1303),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1287),
.A2(n_1321),
.B1(n_1315),
.B2(n_1309),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1295),
.A2(n_1322),
.B(n_1259),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1286),
.B(n_1293),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1244),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1254),
.A2(n_1252),
.B(n_1226),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1276),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1252),
.A2(n_1249),
.B(n_1238),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1191),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1308),
.A2(n_1271),
.B1(n_1253),
.B2(n_1286),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1242),
.A2(n_1245),
.B(n_1234),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1300),
.A2(n_1313),
.B1(n_1320),
.B2(n_1301),
.Y(n_1390)
);

INVx8_ASAP7_75t_L g1391 ( 
.A(n_1305),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1300),
.A2(n_1313),
.B1(n_1303),
.B2(n_1304),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1231),
.A2(n_1240),
.B(n_1267),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1265),
.Y(n_1394)
);

OAI21xp33_ASAP7_75t_L g1395 ( 
.A1(n_1285),
.A2(n_1291),
.B(n_1230),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1222),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1298),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1208),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1304),
.A2(n_1307),
.B1(n_1284),
.B2(n_1289),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1223),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1264),
.A2(n_1204),
.B(n_1256),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1284),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1289),
.A2(n_1233),
.B1(n_1198),
.B2(n_1270),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1243),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1193),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1193),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1312),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1205),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1248),
.B(n_1236),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1274),
.Y(n_1410)
);

AO21x1_ASAP7_75t_L g1411 ( 
.A1(n_1198),
.A2(n_1231),
.B(n_1240),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1317),
.A2(n_1219),
.B1(n_1204),
.B2(n_1199),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1202),
.A2(n_1214),
.B1(n_1193),
.B2(n_1299),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1207),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1220),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1258),
.A2(n_1224),
.B1(n_1269),
.B2(n_1246),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1263),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1215),
.B(n_1263),
.Y(n_1418)
);

INVx8_ASAP7_75t_L g1419 ( 
.A(n_1279),
.Y(n_1419)
);

BUFx2_ASAP7_75t_R g1420 ( 
.A(n_1319),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1294),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1279),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1325),
.A2(n_1192),
.B1(n_1278),
.B2(n_1279),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1279),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1302),
.B(n_1046),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1195),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1275),
.A2(n_1277),
.B(n_1262),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1188),
.B(n_1044),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1188),
.B(n_1044),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1210),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1280),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1302),
.B(n_1046),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1227),
.A2(n_931),
.B1(n_956),
.B2(n_946),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1302),
.A2(n_1328),
.B1(n_1170),
.B2(n_1044),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1250),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1212),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1282),
.Y(n_1441)
);

BUFx2_ASAP7_75t_R g1442 ( 
.A(n_1290),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1288),
.Y(n_1444)
);

BUFx2_ASAP7_75t_SL g1445 ( 
.A(n_1305),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1282),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1195),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1302),
.A2(n_1046),
.B1(n_931),
.B2(n_1328),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1220),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1362),
.B(n_1375),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1419),
.B(n_1424),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1410),
.Y(n_1454)
);

NAND2x1_ASAP7_75t_L g1455 ( 
.A(n_1362),
.B(n_1375),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1382),
.B(n_1344),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1365),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1411),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1363),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1357),
.B(n_1401),
.Y(n_1460)
);

AND2x4_ASAP7_75t_SL g1461 ( 
.A(n_1378),
.B(n_1400),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1367),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1411),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1382),
.B(n_1392),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1373),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1450),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1342),
.Y(n_1467)
);

BUFx4f_ASAP7_75t_SL g1468 ( 
.A(n_1450),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1373),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1339),
.B(n_1357),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1391),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1384),
.A2(n_1427),
.B(n_1386),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1393),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1393),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1364),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1417),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1343),
.B(n_1353),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1419),
.B(n_1424),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1385),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1346),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1430),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1346),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1396),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1359),
.B(n_1348),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1389),
.A2(n_1381),
.B(n_1340),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1401),
.B(n_1439),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1419),
.B(n_1418),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1350),
.B(n_1439),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1417),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1401),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1336),
.B(n_1374),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1441),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1390),
.B(n_1428),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1362),
.B(n_1375),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1370),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1430),
.B(n_1331),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1341),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1438),
.A2(n_1423),
.B(n_1386),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1430),
.B(n_1331),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1376),
.B(n_1425),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1370),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1345),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1381),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1363),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1425),
.B(n_1434),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1434),
.B(n_1372),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1397),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1422),
.A2(n_1394),
.B(n_1368),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1349),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1418),
.B(n_1430),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1444),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1331),
.B(n_1387),
.Y(n_1512)
);

BUFx12f_ASAP7_75t_L g1513 ( 
.A(n_1415),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1369),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1377),
.B(n_1361),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1340),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1397),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1329),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1330),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1395),
.B(n_1354),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1354),
.B(n_1366),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1391),
.B(n_1445),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1332),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1332),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1333),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1338),
.Y(n_1526)
);

OAI211xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1437),
.A2(n_1412),
.B(n_1380),
.C(n_1335),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1426),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1351),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1334),
.A2(n_1449),
.B(n_1446),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1366),
.B(n_1371),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1431),
.A2(n_1433),
.B1(n_1443),
.B2(n_1435),
.C1(n_1436),
.C2(n_1403),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1388),
.A2(n_1399),
.B1(n_1379),
.B2(n_1402),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1429),
.B(n_1409),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1470),
.B(n_1416),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1530),
.A2(n_1360),
.B1(n_1351),
.B2(n_1447),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1470),
.B(n_1394),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1476),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1493),
.B(n_1408),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1473),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1452),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1515),
.A2(n_1409),
.B1(n_1415),
.B2(n_1404),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1486),
.B(n_1448),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1490),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1458),
.B(n_1463),
.Y(n_1545)
);

INVx5_ASAP7_75t_L g1546 ( 
.A(n_1452),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1490),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1460),
.B(n_1474),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1485),
.B(n_1447),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1485),
.B(n_1484),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1523),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1505),
.B(n_1414),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1475),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1451),
.B(n_1378),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1465),
.B(n_1352),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1456),
.B(n_1383),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1479),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1451),
.B(n_1378),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1524),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1469),
.B(n_1398),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1485),
.B(n_1400),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1489),
.B(n_1503),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1506),
.B(n_1454),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1508),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1475),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1489),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1455),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1521),
.B(n_1440),
.Y(n_1569)
);

INVx8_ASAP7_75t_L g1570 ( 
.A(n_1478),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1503),
.B(n_1347),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1513),
.Y(n_1572)
);

BUFx2_ASAP7_75t_SL g1573 ( 
.A(n_1459),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1467),
.B(n_1406),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1521),
.B(n_1405),
.Y(n_1575)
);

INVx5_ASAP7_75t_L g1576 ( 
.A(n_1522),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1488),
.B(n_1405),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1488),
.B(n_1405),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_1551),
.Y(n_1579)
);

AND2x2_ASAP7_75t_SL g1580 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1539),
.B(n_1457),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1536),
.B(n_1527),
.C(n_1532),
.Y(n_1582)
);

AOI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1536),
.A2(n_1534),
.B1(n_1500),
.B2(n_1462),
.C(n_1511),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1559),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1549),
.A2(n_1498),
.B(n_1533),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1559),
.B(n_1483),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1542),
.A2(n_1500),
.B1(n_1491),
.B2(n_1520),
.Y(n_1587)
);

AOI221xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1542),
.A2(n_1464),
.B1(n_1413),
.B2(n_1477),
.C(n_1492),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1560),
.B(n_1509),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1571),
.A2(n_1453),
.B1(n_1510),
.B2(n_1487),
.C(n_1495),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1561),
.A2(n_1466),
.B1(n_1459),
.B2(n_1517),
.C(n_1504),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1535),
.A2(n_1498),
.B(n_1496),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1550),
.B(n_1480),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1549),
.B(n_1482),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1555),
.A2(n_1466),
.B1(n_1504),
.B2(n_1507),
.C(n_1517),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1549),
.B(n_1482),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1564),
.B(n_1552),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1555),
.B(n_1519),
.C(n_1525),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1537),
.B(n_1543),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_1574),
.B(n_1519),
.C(n_1525),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1577),
.A2(n_1499),
.B(n_1461),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1544),
.A2(n_1516),
.B(n_1472),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1554),
.B(n_1558),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1574),
.B(n_1526),
.C(n_1518),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1471),
.C(n_1501),
.Y(n_1605)
);

NAND3xp33_ASAP7_75t_L g1606 ( 
.A(n_1557),
.B(n_1528),
.C(n_1514),
.Y(n_1606)
);

OAI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1556),
.A2(n_1531),
.B(n_1420),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1553),
.B(n_1566),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1577),
.A2(n_1512),
.B1(n_1499),
.B2(n_1494),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1547),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1570),
.A2(n_1494),
.B1(n_1510),
.B2(n_1468),
.Y(n_1611)
);

AND2x2_ASAP7_75t_SL g1612 ( 
.A(n_1538),
.B(n_1481),
.Y(n_1612)
);

OAI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1556),
.A2(n_1497),
.B(n_1502),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1548),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1610),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1610),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1606),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1606),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1602),
.Y(n_1620)
);

AND3x1_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1578),
.C(n_1575),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1593),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1594),
.B(n_1563),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1594),
.B(n_1563),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1612),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1597),
.B(n_1545),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1588),
.B(n_1554),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1599),
.B(n_1565),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1596),
.B(n_1567),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1567),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1608),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1600),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1605),
.B(n_1576),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1581),
.B(n_1540),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1599),
.B(n_1565),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1580),
.B(n_1612),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1580),
.B(n_1569),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1604),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1598),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1617),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1637),
.B(n_1580),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1641),
.B(n_1582),
.C(n_1588),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1637),
.B(n_1583),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1634),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1572),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1614),
.B(n_1513),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1625),
.B(n_1612),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1616),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1616),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1623),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1627),
.A2(n_1582),
.B1(n_1585),
.B2(n_1592),
.C(n_1591),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1635),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1625),
.B(n_1603),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1635),
.Y(n_1659)
);

AND2x6_ASAP7_75t_SL g1660 ( 
.A(n_1634),
.B(n_1337),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1628),
.B(n_1608),
.Y(n_1661)
);

OR4x1_ASAP7_75t_L g1662 ( 
.A(n_1618),
.B(n_1619),
.C(n_1642),
.D(n_1641),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1642),
.B(n_1632),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1634),
.B(n_1568),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1623),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1620),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1624),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1640),
.B(n_1586),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1620),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1632),
.B(n_1613),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1640),
.B(n_1639),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1624),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1639),
.B(n_1589),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1629),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1613),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1629),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1630),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1630),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1442),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1636),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1644),
.B(n_1636),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1663),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1663),
.B(n_1671),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_SL g1685 ( 
.A(n_1645),
.B(n_1590),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1671),
.B(n_1670),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1651),
.B(n_1638),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1618),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1643),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1648),
.B(n_1664),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1651),
.B(n_1638),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1670),
.B(n_1675),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1675),
.B(n_1633),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_SL g1694 ( 
.A(n_1656),
.B(n_1573),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1648),
.B(n_1631),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1643),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1648),
.B(n_1631),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1653),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1648),
.B(n_1655),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1664),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1646),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1646),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1664),
.B(n_1634),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1674),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1655),
.B(n_1622),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1664),
.B(n_1546),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1622),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1619),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1659),
.B(n_1615),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1656),
.A2(n_1585),
.B1(n_1592),
.B2(n_1595),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1665),
.B(n_1667),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1668),
.B(n_1615),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1676),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1666),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1666),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1676),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1668),
.B(n_1626),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1669),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1677),
.Y(n_1721)
);

OAI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1647),
.A2(n_1621),
.B(n_1607),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1649),
.B(n_1621),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1689),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1689),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1697),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1697),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1690),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1680),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1722),
.B(n_1673),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1673),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1681),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1688),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1702),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1686),
.B(n_1667),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1722),
.A2(n_1611),
.B1(n_1609),
.B2(n_1658),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1702),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1703),
.Y(n_1739)
);

AND3x2_ASAP7_75t_L g1740 ( 
.A(n_1685),
.B(n_1662),
.C(n_1658),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1681),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1685),
.B(n_1672),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1690),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1703),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1687),
.B(n_1677),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1694),
.A2(n_1607),
.B1(n_1570),
.B2(n_1541),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1682),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1705),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1705),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1692),
.B(n_1678),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1714),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1692),
.B(n_1683),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1686),
.B(n_1678),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1714),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1690),
.B(n_1652),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1691),
.B(n_1661),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1684),
.B(n_1652),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1691),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1715),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1715),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1734),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1759),
.B(n_1690),
.Y(n_1763)
);

AOI21xp33_ASAP7_75t_L g1764 ( 
.A1(n_1731),
.A2(n_1694),
.B(n_1711),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1740),
.B(n_1693),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1724),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1732),
.B(n_1723),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1742),
.A2(n_1662),
.B1(n_1693),
.B2(n_1709),
.C(n_1684),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1744),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

OAI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1737),
.A2(n_1707),
.B1(n_1709),
.B2(n_1701),
.C(n_1718),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1744),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1725),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1757),
.B(n_1704),
.Y(n_1776)
);

NAND5xp2_ASAP7_75t_L g1777 ( 
.A(n_1747),
.B(n_1707),
.C(n_1679),
.D(n_1700),
.E(n_1696),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1757),
.A2(n_1698),
.B(n_1696),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1753),
.B(n_1700),
.Y(n_1779)
);

OAI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1751),
.A2(n_1707),
.B1(n_1721),
.B2(n_1718),
.C(n_1698),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1756),
.B(n_1704),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1704),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1746),
.A2(n_1719),
.B(n_1713),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1725),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1729),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1754),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1729),
.A2(n_1704),
.B(n_1601),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1756),
.B(n_1721),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1754),
.A2(n_1710),
.B(n_1719),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1764),
.A2(n_1741),
.B1(n_1730),
.B2(n_1733),
.C(n_1761),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1776),
.B(n_1746),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1785),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1769),
.B(n_1736),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1785),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1777),
.A2(n_1730),
.B1(n_1741),
.B2(n_1733),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1762),
.B(n_1743),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1772),
.B(n_1743),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1774),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1786),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1763),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1770),
.B(n_1736),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1772),
.B(n_1750),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1766),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1782),
.B(n_1712),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1771),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1775),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1772),
.B(n_1712),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1767),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1784),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1768),
.A2(n_1758),
.B1(n_1752),
.B2(n_1755),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1796),
.B(n_1779),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1793),
.A2(n_1768),
.B1(n_1765),
.B2(n_1773),
.C(n_1780),
.Y(n_1812)
);

AOI211xp5_ASAP7_75t_L g1813 ( 
.A1(n_1799),
.A2(n_1781),
.B(n_1787),
.C(n_1788),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1797),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1810),
.A2(n_1781),
.B1(n_1778),
.B2(n_1782),
.C(n_1783),
.Y(n_1815)
);

AOI322xp5_ASAP7_75t_L g1816 ( 
.A1(n_1795),
.A2(n_1788),
.A3(n_1774),
.B1(n_1767),
.B2(n_1752),
.C1(n_1749),
.C2(n_1760),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1800),
.A2(n_1782),
.B1(n_1767),
.B2(n_1789),
.Y(n_1817)
);

NOR3xp33_ASAP7_75t_L g1818 ( 
.A(n_1801),
.B(n_1755),
.C(n_1749),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1808),
.A2(n_1713),
.B1(n_1710),
.B2(n_1758),
.Y(n_1819)
);

NOR3x1_ASAP7_75t_L g1820 ( 
.A(n_1802),
.B(n_1761),
.C(n_1760),
.Y(n_1820)
);

NAND4xp25_ASAP7_75t_L g1821 ( 
.A(n_1790),
.B(n_1727),
.C(n_1735),
.D(n_1726),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1807),
.A2(n_1727),
.B1(n_1745),
.B2(n_1739),
.C(n_1738),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1808),
.B(n_1660),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1797),
.A2(n_1735),
.B(n_1726),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1814),
.B(n_1797),
.Y(n_1825)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1826 ( 
.A1(n_1815),
.A2(n_1809),
.B(n_1803),
.C(n_1805),
.D(n_1806),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1811),
.Y(n_1827)
);

NOR3xp33_ASAP7_75t_L g1828 ( 
.A(n_1812),
.B(n_1798),
.C(n_1794),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1816),
.B(n_1794),
.C(n_1792),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1813),
.B(n_1792),
.C(n_1803),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1823),
.B(n_1791),
.Y(n_1831)
);

NOR2x1p5_ASAP7_75t_L g1832 ( 
.A(n_1821),
.B(n_1805),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1824),
.Y(n_1833)
);

NOR3x1_ASAP7_75t_L g1834 ( 
.A(n_1822),
.B(n_1809),
.C(n_1739),
.Y(n_1834)
);

NAND2x1p5_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1407),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1819),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_R g1837 ( 
.A(n_1827),
.B(n_1421),
.Y(n_1837)
);

AOI32xp33_ASAP7_75t_L g1838 ( 
.A1(n_1828),
.A2(n_1836),
.A3(n_1818),
.B1(n_1831),
.B2(n_1833),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1829),
.A2(n_1817),
.B1(n_1804),
.B2(n_1791),
.Y(n_1839)
);

OAI21xp33_ASAP7_75t_L g1840 ( 
.A1(n_1825),
.A2(n_1804),
.B(n_1745),
.Y(n_1840)
);

NAND4xp25_ASAP7_75t_L g1841 ( 
.A(n_1830),
.B(n_1738),
.C(n_1748),
.D(n_1407),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1835),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1839),
.A2(n_1832),
.B1(n_1826),
.B2(n_1748),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1842),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1840),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1841),
.A2(n_1826),
.B1(n_1706),
.B2(n_1708),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1838),
.B(n_1834),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1837),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1842),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1844),
.B(n_1706),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1849),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_L g1852 ( 
.A(n_1847),
.B(n_1432),
.C(n_1406),
.Y(n_1852)
);

NOR3xp33_ASAP7_75t_L g1853 ( 
.A(n_1845),
.B(n_1432),
.C(n_1358),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1843),
.B(n_1708),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_L g1855 ( 
.A(n_1848),
.B(n_1358),
.C(n_1682),
.Y(n_1855)
);

NAND2x1_ASAP7_75t_L g1856 ( 
.A(n_1850),
.B(n_1846),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1854),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1851),
.B(n_1654),
.Y(n_1858)
);

XOR2x2_ASAP7_75t_L g1859 ( 
.A(n_1852),
.B(n_1358),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1857),
.Y(n_1860)
);

XOR2xp5_ASAP7_75t_L g1861 ( 
.A(n_1859),
.B(n_1853),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1860),
.A2(n_1856),
.B1(n_1858),
.B2(n_1421),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1862),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1862),
.A2(n_1861),
.B(n_1855),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1863),
.A2(n_1682),
.B1(n_1695),
.B2(n_1699),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1864),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1866),
.A2(n_1720),
.B1(n_1695),
.B2(n_1699),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1865),
.B(n_1699),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1868),
.Y(n_1869)
);

OAI221xp5_ASAP7_75t_R g1870 ( 
.A1(n_1869),
.A2(n_1660),
.B1(n_1720),
.B2(n_1695),
.C(n_1717),
.Y(n_1870)
);

AOI211xp5_ASAP7_75t_L g1871 ( 
.A1(n_1870),
.A2(n_1720),
.B(n_1717),
.C(n_1716),
.Y(n_1871)
);


endmodule