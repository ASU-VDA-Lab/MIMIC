module fake_jpeg_12263_n_589 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_589);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_67),
.Y(n_132)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_77),
.Y(n_134)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_16),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_85),
.Y(n_182)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_35),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_87),
.B(n_97),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_35),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_99),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_35),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_33),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_111),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_33),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_113),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_41),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_115),
.Y(n_148)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_41),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_22),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_121),
.B(n_18),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_72),
.A2(n_52),
.B1(n_48),
.B2(n_34),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_130),
.A2(n_139),
.B1(n_66),
.B2(n_117),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_58),
.A2(n_48),
.B1(n_53),
.B2(n_57),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_78),
.A2(n_79),
.B1(n_84),
.B2(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_143),
.A2(n_191),
.B1(n_24),
.B2(n_37),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_39),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_184),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_109),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_156),
.B(n_183),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_60),
.A2(n_57),
.B1(n_53),
.B2(n_46),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_42),
.B1(n_47),
.B2(n_43),
.Y(n_207)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g167 ( 
.A(n_103),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_167),
.Y(n_204)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_59),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

AND2x4_ASAP7_75t_SL g175 ( 
.A(n_94),
.B(n_42),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_175),
.B(n_73),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_187),
.Y(n_208)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_103),
.B(n_18),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_107),
.B(n_20),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_46),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_75),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_195),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_119),
.A2(n_47),
.B1(n_43),
.B2(n_39),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_69),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_75),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_118),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_110),
.Y(n_213)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_198),
.Y(n_300)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_200),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_62),
.B1(n_74),
.B2(n_108),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_201),
.A2(n_207),
.B1(n_212),
.B2(n_266),
.Y(n_293)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_205),
.Y(n_314)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_206),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_130),
.A2(n_86),
.B1(n_90),
.B2(n_105),
.Y(n_212)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

CKINVDCx12_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_217),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_160),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_218),
.B(n_245),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_20),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_219),
.B(n_222),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_137),
.B(n_37),
.Y(n_222)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_228),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_239),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_154),
.A2(n_116),
.B1(n_114),
.B2(n_70),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_136),
.Y(n_231)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_231),
.Y(n_287)
);

BUFx4f_ASAP7_75t_SL g232 ( 
.A(n_127),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_232),
.Y(n_279)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_154),
.Y(n_233)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_242),
.Y(n_278)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_235),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_120),
.B1(n_28),
.B2(n_29),
.Y(n_236)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_24),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_R g271 ( 
.A(n_238),
.B(n_246),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_179),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_175),
.B(n_65),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_123),
.Y(n_243)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_255),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_160),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_30),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_124),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_251),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_134),
.B(n_110),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_250),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_140),
.B(n_104),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_159),
.A2(n_15),
.B(n_16),
.Y(n_252)
);

AOI32xp33_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_0),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_162),
.A2(n_27),
.B1(n_28),
.B2(n_89),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_139),
.B1(n_190),
.B2(n_171),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_126),
.B(n_15),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_164),
.B(n_159),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_256),
.B(n_143),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_144),
.B(n_0),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_261),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_138),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_171),
.Y(n_276)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_259),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_148),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_260),
.Y(n_316)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_141),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_164),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_263),
.Y(n_292)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_152),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_132),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_158),
.A2(n_92),
.B1(n_85),
.B2(n_82),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_201),
.A2(n_168),
.B1(n_190),
.B2(n_169),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_270),
.A2(n_301),
.B1(n_311),
.B2(n_263),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_272),
.A2(n_304),
.B1(n_320),
.B2(n_231),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_276),
.Y(n_357)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_281),
.B(n_278),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_242),
.A2(n_133),
.B(n_153),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_283),
.A2(n_310),
.B(n_204),
.Y(n_349)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_234),
.A2(n_185),
.B1(n_125),
.B2(n_181),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_284),
.B(n_211),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_122),
.B(n_102),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_286),
.B(n_302),
.C(n_322),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_256),
.A2(n_169),
.B1(n_152),
.B2(n_128),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_215),
.B(n_122),
.C(n_76),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_229),
.A2(n_174),
.B1(n_157),
.B2(n_194),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_209),
.B(n_174),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_309),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_0),
.C(n_6),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_250),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_250),
.A2(n_186),
.B(n_128),
.C(n_194),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_208),
.A2(n_186),
.B1(n_166),
.B2(n_182),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_236),
.A2(n_182),
.B1(n_172),
.B2(n_166),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_235),
.A2(n_0),
.B(n_5),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_274),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_324),
.B(n_328),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_342),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_304),
.A2(n_172),
.B1(n_237),
.B2(n_220),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_329),
.B1(n_358),
.B2(n_362),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_258),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_333),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_232),
.Y(n_328)
);

BUFx4f_ASAP7_75t_SL g330 ( 
.A(n_314),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_271),
.B(n_312),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_239),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_278),
.A2(n_232),
.B(n_225),
.C(n_233),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_338),
.Y(n_369)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_210),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_336),
.B(n_341),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_267),
.B(n_251),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_268),
.Y(n_339)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_253),
.B1(n_230),
.B2(n_200),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_340),
.A2(n_364),
.B1(n_276),
.B2(n_310),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_271),
.B(n_204),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_343),
.Y(n_371)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_344),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_210),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_277),
.B(n_267),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_346),
.Y(n_395)
);

INVx13_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_278),
.B(n_308),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_353),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_284),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_248),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_359),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_241),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_356),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_308),
.A2(n_216),
.B1(n_203),
.B2(n_221),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_302),
.B(n_248),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_319),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_365),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_315),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_361),
.A2(n_363),
.B1(n_282),
.B2(n_303),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_308),
.A2(n_224),
.B1(n_254),
.B2(n_223),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_293),
.A2(n_240),
.B1(n_254),
.B2(n_223),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_281),
.B(n_261),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_359),
.C(n_323),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_375),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_373),
.A2(n_398),
.B(n_303),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_309),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_283),
.C(n_286),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_378),
.B(n_381),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_322),
.C(n_276),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_394),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_327),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_396),
.Y(n_406)
);

XNOR2x2_ASAP7_75t_SL g390 ( 
.A(n_341),
.B(n_284),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_331),
.B(n_360),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_293),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_307),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_325),
.B(n_276),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_401),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_364),
.A2(n_321),
.B1(n_279),
.B2(n_291),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_400),
.A2(n_403),
.B1(n_362),
.B2(n_287),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_313),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_342),
.A2(n_291),
.B1(n_280),
.B2(n_298),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_379),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_405),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_346),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_329),
.B1(n_334),
.B2(n_335),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_420),
.B1(n_427),
.B2(n_403),
.Y(n_440)
);

AND2x4_ASAP7_75t_SL g409 ( 
.A(n_396),
.B(n_357),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_425),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_371),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_398),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

CKINVDCx10_ASAP7_75t_R g413 ( 
.A(n_399),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_413),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_401),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_343),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_416),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_385),
.B(n_339),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_358),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_369),
.A2(n_287),
.B(n_344),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_419),
.A2(n_410),
.B(n_406),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_394),
.A2(n_361),
.B1(n_363),
.B2(n_348),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_368),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_429),
.Y(n_445)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_423),
.A2(n_384),
.B1(n_383),
.B2(n_371),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_367),
.A2(n_361),
.B1(n_290),
.B2(n_275),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_426),
.A2(n_373),
.B(n_397),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_377),
.A2(n_280),
.B1(n_355),
.B2(n_288),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_388),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_298),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_376),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_434),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_372),
.B(n_375),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_378),
.C(n_373),
.Y(n_444)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_376),
.B(n_294),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_369),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_436),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_368),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

AOI322xp5_ASAP7_75t_L g438 ( 
.A1(n_390),
.A2(n_288),
.A3(n_347),
.B1(n_290),
.B2(n_289),
.C1(n_314),
.C2(n_296),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_438),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_440),
.A2(n_453),
.B1(n_417),
.B2(n_428),
.Y(n_484)
);

MAJx2_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_433),
.C(n_409),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_454),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_408),
.B(n_382),
.Y(n_450)
);

XNOR2x1_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_458),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_452),
.A2(n_420),
.B1(n_426),
.B2(n_419),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_436),
.A2(n_383),
.B1(n_400),
.B2(n_384),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_412),
.A2(n_381),
.B(n_380),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_380),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_459),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_399),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_460),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_414),
.B(n_366),
.Y(n_461)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_432),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_468),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_406),
.B(n_366),
.Y(n_465)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_370),
.Y(n_467)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_431),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_471),
.Y(n_501)
);

XOR2x2_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_433),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_481),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_474),
.A2(n_453),
.B1(n_443),
.B2(n_442),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_461),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_445),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_447),
.A2(n_412),
.B1(n_418),
.B2(n_423),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_493),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_408),
.C(n_409),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_488),
.C(n_489),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_425),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_410),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_484),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_413),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_427),
.C(n_418),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_437),
.C(n_317),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_462),
.C(n_443),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_462),
.C(n_467),
.Y(n_500)
);

XOR2x1_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_354),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_491),
.B(n_451),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_462),
.A2(n_393),
.B1(n_300),
.B2(n_228),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_317),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_479),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_502),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_499),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_500),
.B(n_507),
.Y(n_531)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_503),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_486),
.B(n_465),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_512),
.Y(n_528)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_506),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_492),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_442),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_481),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_451),
.C(n_469),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_514),
.C(n_515),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_485),
.A2(n_468),
.B1(n_448),
.B2(n_449),
.Y(n_511)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_478),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_441),
.Y(n_513)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_513),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_439),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_473),
.C(n_471),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_466),
.Y(n_517)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_517),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_488),
.A2(n_469),
.B1(n_456),
.B2(n_393),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_518),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_523),
.A2(n_525),
.B(n_498),
.Y(n_542)
);

A2O1A1Ixp33_ASAP7_75t_SL g525 ( 
.A1(n_503),
.A2(n_491),
.B(n_508),
.C(n_498),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_494),
.Y(n_526)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_526),
.Y(n_537)
);

NOR4xp25_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_480),
.C(n_476),
.D(n_493),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_529),
.A2(n_518),
.B1(n_515),
.B2(n_505),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_456),
.C(n_482),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_532),
.B(n_535),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_463),
.Y(n_534)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_534),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_330),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_496),
.C(n_516),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_538),
.B(n_543),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_519),
.B(n_527),
.Y(n_540)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_540),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_523),
.B(n_509),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_548),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_542),
.B(n_520),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_501),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_544),
.A2(n_549),
.B(n_550),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_502),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_545),
.B(n_547),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_460),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_449),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_448),
.B(n_330),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_522),
.B(n_315),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_528),
.B(n_300),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_551),
.B(n_525),
.C(n_533),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_539),
.C(n_550),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_556),
.Y(n_569)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_555),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_533),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_542),
.Y(n_564)
);

BUFx24_ASAP7_75t_SL g558 ( 
.A(n_540),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_558),
.B(n_526),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_536),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_562),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_524),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_564),
.B(n_205),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_552),
.B(n_521),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_565),
.B(n_205),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_560),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_525),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_567),
.A2(n_555),
.B(n_559),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_563),
.B(n_289),
.Y(n_571)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_571),
.Y(n_573)
);

AOI31xp67_ASAP7_75t_L g572 ( 
.A1(n_554),
.A2(n_525),
.A3(n_206),
.B(n_198),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_572),
.B(n_569),
.Y(n_578)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_574),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_575),
.A2(n_577),
.B(n_578),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_576),
.B(n_567),
.C(n_570),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_579),
.A2(n_582),
.B(n_7),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_SL g582 ( 
.A(n_573),
.B(n_568),
.C(n_564),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_583),
.B(n_584),
.Y(n_585)
);

AOI322xp5_ASAP7_75t_L g584 ( 
.A1(n_581),
.A2(n_7),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_14),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_585),
.A2(n_580),
.B(n_10),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_586),
.B(n_7),
.C(n_11),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_12),
.C(n_14),
.Y(n_588)
);

OAI31xp33_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_12),
.A3(n_14),
.B(n_572),
.Y(n_589)
);


endmodule