module fake_netlist_6_2449_n_1815 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1815);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1815;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_95),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_10),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_154),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_12),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_8),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_69),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_64),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_48),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_58),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_47),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_54),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_21),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_72),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_24),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_87),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_31),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_70),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_92),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_121),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_111),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_125),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_2),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_62),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_133),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_47),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_88),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_53),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_4),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_68),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_66),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_120),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_21),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_131),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_50),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_122),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_37),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_19),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_135),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_91),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_114),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_20),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_112),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_51),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_97),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_33),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_113),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_48),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_75),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_79),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_8),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_157),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_49),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_59),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_90),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_4),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_130),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_14),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_129),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_35),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_141),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_132),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_35),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_145),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_152),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_105),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_56),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_17),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_89),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_73),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_36),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_123),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_77),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_49),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_9),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_37),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_19),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_74),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_10),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_29),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_150),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_29),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_34),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_119),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_83),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_57),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_86),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_158),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_98),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_38),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_46),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_99),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_94),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_156),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_3),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_103),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_140),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_109),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_128),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_24),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_39),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_115),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_1),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_20),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_55),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_7),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_110),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_93),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_188),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_282),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_203),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_163),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_218),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_190),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_191),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_180),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_169),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_205),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_159),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_192),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_242),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_229),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_229),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_230),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_193),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_170),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_172),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_213),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_290),
.Y(n_351)
);

BUFx2_ASAP7_75t_SL g352 ( 
.A(n_233),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_302),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_196),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_221),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_222),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_223),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_173),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_240),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_254),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_259),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_283),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_176),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_178),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_197),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_178),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_226),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_189),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_185),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_189),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_187),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g374 ( 
.A(n_195),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_198),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_209),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_209),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_225),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_225),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_239),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_239),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_226),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_208),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_249),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_249),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_186),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_264),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_264),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_281),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_281),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_231),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_324),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_320),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_317),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_161),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_351),
.A2(n_183),
.B1(n_314),
.B2(n_175),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_317),
.B(n_322),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_296),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_235),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_330),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_247),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_253),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_337),
.B(n_260),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_354),
.B(n_162),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_364),
.B(n_176),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_177),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_319),
.B(n_176),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_323),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_286),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_334),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_366),
.Y(n_425)
);

CKINVDCx6p67_ASAP7_75t_R g426 ( 
.A(n_364),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_375),
.B(n_287),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_352),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_321),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_331),
.B(n_347),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_337),
.B(n_294),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_371),
.B(n_315),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_358),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_376),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_328),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_377),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_316),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_378),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_379),
.B(n_177),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_335),
.B(n_177),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_325),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_358),
.B(n_177),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_358),
.B(n_177),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_395),
.Y(n_463)
);

BUFx4f_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_427),
.Y(n_465)
);

AO22x1_ASAP7_75t_L g466 ( 
.A1(n_408),
.A2(n_383),
.B1(n_183),
.B2(n_175),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_L g467 ( 
.A1(n_412),
.A2(n_374),
.B1(n_373),
.B2(n_327),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_402),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

AO22x1_ASAP7_75t_L g473 ( 
.A1(n_408),
.A2(n_171),
.B1(n_168),
.B2(n_164),
.Y(n_473)
);

AND3x2_ASAP7_75t_L g474 ( 
.A(n_410),
.B(n_316),
.C(n_448),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_406),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_441),
.A2(n_391),
.B1(n_364),
.B2(n_389),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_416),
.B(n_391),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_409),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_399),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_422),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_399),
.B(n_384),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_438),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_397),
.A2(n_303),
.B1(n_168),
.B2(n_309),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_356),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_415),
.B(n_385),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_403),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

AND2x4_ASAP7_75t_SL g495 ( 
.A(n_426),
.B(n_206),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_421),
.B(n_206),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_446),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_415),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_431),
.B(n_206),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_435),
.B(n_238),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_394),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_433),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_408),
.B(n_385),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_401),
.B(n_364),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_394),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_404),
.B(n_238),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_397),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_456),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_438),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_405),
.A2(n_199),
.B1(n_280),
.B2(n_277),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_419),
.B(n_238),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_338),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_423),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_394),
.B(n_387),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_408),
.A2(n_389),
.B1(n_388),
.B2(n_387),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_417),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_440),
.A2(n_461),
.B1(n_459),
.B2(n_456),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_394),
.B(n_388),
.Y(n_523)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_457),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_440),
.B(n_424),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_440),
.B(n_390),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_398),
.A2(n_440),
.B(n_411),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_459),
.A2(n_390),
.B1(n_365),
.B2(n_363),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_396),
.B(n_344),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_436),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_459),
.B(n_291),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_436),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_442),
.Y(n_537)
);

AO21x2_ASAP7_75t_L g538 ( 
.A1(n_398),
.A2(n_461),
.B(n_459),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_414),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_436),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_461),
.A2(n_171),
.B1(n_164),
.B2(n_161),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_456),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_413),
.B(n_160),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_442),
.B(n_174),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_456),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_461),
.B(n_291),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_393),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_393),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_418),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_393),
.Y(n_552)
);

AO21x2_ASAP7_75t_L g553 ( 
.A1(n_424),
.A2(n_350),
.B(n_349),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_427),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_425),
.B(n_349),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_418),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_442),
.B(n_353),
.Y(n_557)
);

AO22x2_ASAP7_75t_L g558 ( 
.A1(n_425),
.A2(n_202),
.B1(n_220),
.B2(n_228),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_418),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_393),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_426),
.B(n_251),
.Y(n_561)
);

AND3x1_ASAP7_75t_L g562 ( 
.A(n_428),
.B(n_355),
.C(n_350),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_428),
.A2(n_234),
.B1(n_217),
.B2(n_219),
.Y(n_563)
);

INVx4_ASAP7_75t_SL g564 ( 
.A(n_413),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_413),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_418),
.B(n_258),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_420),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_393),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_458),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_413),
.A2(n_365),
.B(n_363),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_437),
.B(n_160),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_393),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_420),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_420),
.B(n_200),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_439),
.B(n_336),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_413),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_427),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_429),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_400),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_420),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_420),
.B(n_291),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_444),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_400),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_400),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_400),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_400),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_432),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_444),
.B(n_355),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_450),
.B(n_336),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_432),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_450),
.B(n_357),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_432),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_400),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_432),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_451),
.A2(n_272),
.B1(n_194),
.B2(n_201),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_432),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_458),
.B(n_207),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_451),
.B(n_165),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_447),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_447),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_447),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_447),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_447),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_458),
.B(n_210),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_525),
.B(n_357),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_571),
.B(n_226),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_496),
.B(n_359),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_571),
.B(n_454),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_597),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_499),
.B(n_482),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_597),
.B(n_454),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_553),
.A2(n_226),
.B1(n_413),
.B2(n_453),
.Y(n_621)
);

AOI221xp5_ASAP7_75t_L g622 ( 
.A1(n_509),
.A2(n_301),
.B1(n_307),
.B2(n_309),
.C(n_310),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_499),
.B(n_226),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_482),
.B(n_587),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_526),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_525),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_533),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_522),
.B(n_547),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_468),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_463),
.B(n_471),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_578),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_579),
.B(n_165),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_547),
.B(n_226),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_606),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_567),
.B(n_226),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_498),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_463),
.B(n_226),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_498),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_491),
.B(n_359),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_606),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_580),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_497),
.B(n_301),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_490),
.B(n_360),
.Y(n_643)
);

AO22x2_ASAP7_75t_L g644 ( 
.A1(n_490),
.A2(n_362),
.B1(n_361),
.B2(n_360),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_471),
.B(n_454),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_472),
.B(n_211),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_580),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_472),
.B(n_454),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_480),
.B(n_212),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_478),
.B(n_166),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_533),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_480),
.B(n_454),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_526),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_515),
.B(n_166),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_594),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_505),
.B(n_361),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_534),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_481),
.B(n_214),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_594),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_504),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_502),
.B(n_167),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_491),
.B(n_362),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_481),
.B(n_215),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_553),
.A2(n_413),
.B1(n_310),
.B2(n_312),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_484),
.B(n_454),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_468),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_484),
.B(n_460),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_526),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_485),
.B(n_460),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_534),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_536),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_485),
.B(n_460),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_567),
.B(n_503),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_494),
.B(n_460),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_460),
.Y(n_675)
);

AOI221xp5_ASAP7_75t_L g676 ( 
.A1(n_558),
.A2(n_307),
.B1(n_312),
.B2(n_314),
.C(n_262),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_505),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_469),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_511),
.B(n_460),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_511),
.B(n_462),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_527),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_516),
.B(n_462),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_467),
.B(n_167),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_527),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_555),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_561),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_504),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_553),
.A2(n_292),
.B1(n_261),
.B2(n_265),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_524),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_555),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_486),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_516),
.B(n_462),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_493),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_558),
.A2(n_298),
.B1(n_227),
.B2(n_236),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_466),
.B(n_204),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_466),
.B(n_245),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_495),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_555),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_486),
.B(n_340),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_493),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_536),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_493),
.B(n_340),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_506),
.A2(n_279),
.B1(n_216),
.B2(n_232),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_SL g704 ( 
.A(n_501),
.B(n_248),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_555),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_565),
.B(n_241),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_513),
.B(n_179),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_493),
.B(n_342),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_528),
.B(n_462),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_528),
.B(n_462),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_510),
.A2(n_184),
.B1(n_181),
.B2(n_182),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_528),
.B(n_462),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_469),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_565),
.B(n_243),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_583),
.B(n_455),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_557),
.A2(n_288),
.B1(n_244),
.B2(n_246),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_593),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_583),
.B(n_429),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_503),
.B(n_455),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_565),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_507),
.B(n_434),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_531),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_593),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_507),
.B(n_434),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_537),
.B(n_443),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_510),
.A2(n_543),
.B1(n_541),
.B2(n_514),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_558),
.A2(n_250),
.B1(n_275),
.B2(n_299),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_537),
.B(n_443),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_565),
.B(n_581),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_604),
.B(n_445),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_540),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_612),
.B(n_546),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_541),
.A2(n_276),
.B1(n_255),
.B2(n_256),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_476),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_508),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_SL g736 ( 
.A(n_489),
.B(n_289),
.C(n_252),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_605),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_574),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_538),
.B(n_445),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_581),
.B(n_257),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_538),
.B(n_449),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_538),
.B(n_449),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_558),
.A2(n_274),
.B1(n_271),
.B2(n_269),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_539),
.B(n_263),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_593),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_593),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_596),
.B(n_342),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_539),
.B(n_295),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_489),
.B(n_268),
.C(n_237),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_473),
.B(n_348),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_596),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_544),
.B(n_297),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_540),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_596),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_543),
.A2(n_266),
.B1(n_267),
.B2(n_273),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_487),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_544),
.B(n_285),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_596),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_518),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_473),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_551),
.B(n_452),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_581),
.B(n_305),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_523),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_567),
.A2(n_348),
.B1(n_346),
.B2(n_343),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_551),
.B(n_452),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_556),
.B(n_452),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_477),
.A2(n_304),
.B1(n_181),
.B2(n_182),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_556),
.B(n_452),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_519),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_577),
.A2(n_305),
.B(n_184),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_487),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_559),
.B(n_452),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_559),
.B(n_452),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_563),
.B(n_313),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_568),
.B(n_452),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_581),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_474),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_567),
.B(n_308),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_573),
.B(n_549),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_568),
.B(n_308),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_562),
.B(n_346),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_476),
.B(n_179),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_562),
.B(n_343),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_549),
.B(n_311),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_470),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_572),
.B(n_313),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_616),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_690),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_624),
.B(n_495),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_624),
.B(n_495),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_738),
.B(n_519),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_SL g792 ( 
.A(n_654),
.B(n_542),
.C(n_548),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_654),
.B(n_572),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_698),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_660),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_723),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_745),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_618),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_746),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_628),
.A2(n_567),
.B1(n_535),
.B2(n_586),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_664),
.A2(n_567),
.B1(n_542),
.B2(n_483),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_660),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_650),
.B(n_576),
.Y(n_805)
);

NAND2x2_ASAP7_75t_L g806 ( 
.A(n_777),
.B(n_601),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_629),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_626),
.B(n_677),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_751),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_754),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_758),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_687),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_638),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_722),
.B(n_576),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_685),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_691),
.B(n_529),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_685),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_650),
.B(n_585),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_683),
.A2(n_707),
.B(n_774),
.C(n_717),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_643),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_717),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_629),
.Y(n_822)
);

AND2x6_ASAP7_75t_L g823 ( 
.A(n_720),
.B(n_603),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_666),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_660),
.B(n_608),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_681),
.B(n_564),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_666),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_631),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_668),
.Y(n_829)
);

AND2x4_ASAP7_75t_SL g830 ( 
.A(n_702),
.B(n_520),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_653),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_732),
.B(n_585),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_684),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_634),
.B(n_567),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_640),
.B(n_759),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_664),
.A2(n_483),
.B1(n_521),
.B2(n_530),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_736),
.A2(n_521),
.B1(n_530),
.B2(n_532),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_769),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_763),
.B(n_600),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_688),
.A2(n_532),
.B1(n_512),
.B2(n_488),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_653),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_628),
.A2(n_600),
.B1(n_590),
.B2(n_588),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_630),
.B(n_588),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_708),
.B(n_464),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_678),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_678),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_705),
.B(n_590),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_709),
.A2(n_464),
.B(n_500),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_688),
.A2(n_488),
.B1(n_512),
.B2(n_545),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_614),
.B(n_564),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_747),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_715),
.Y(n_854)
);

NOR2x2_ASAP7_75t_L g855 ( 
.A(n_694),
.B(n_550),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_676),
.A2(n_569),
.B1(n_550),
.B2(n_552),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_641),
.B(n_647),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_655),
.B(n_591),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_689),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_693),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_713),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_700),
.B(n_608),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_639),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_668),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_SL g865 ( 
.A(n_694),
.B(n_237),
.C(n_300),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_662),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

CKINVDCx8_ASAP7_75t_R g868 ( 
.A(n_781),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_686),
.B(n_699),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_718),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_683),
.A2(n_591),
.B(n_603),
.C(n_552),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_614),
.B(n_464),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_656),
.B(n_659),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_710),
.B(n_554),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_760),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_632),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_SL g877 ( 
.A(n_697),
.B(n_300),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_712),
.B(n_554),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_656),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_737),
.B(n_500),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_SL g881 ( 
.A(n_749),
.B(n_304),
.C(n_311),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_668),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_781),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_619),
.B(n_500),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_632),
.B(n_554),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_734),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_619),
.B(n_564),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_783),
.B(n_564),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_783),
.B(n_566),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_720),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_734),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_617),
.B(n_554),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_735),
.B(n_609),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_750),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_620),
.B(n_582),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_695),
.B(n_582),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_720),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_785),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_SL g899 ( 
.A(n_774),
.B(n_1),
.C(n_2),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_739),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_627),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_716),
.B(n_613),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_741),
.A2(n_599),
.B(n_589),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_644),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_651),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_742),
.B(n_582),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_657),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_SL g908 ( 
.A(n_696),
.B(n_560),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_727),
.A2(n_743),
.B1(n_707),
.B2(n_622),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_661),
.A2(n_584),
.B(n_560),
.C(n_569),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_726),
.B(n_566),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_670),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_661),
.A2(n_584),
.B(n_575),
.C(n_589),
.Y(n_913)
);

CKINVDCx8_ASAP7_75t_R g914 ( 
.A(n_644),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_730),
.B(n_625),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_671),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_701),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_756),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_633),
.B(n_566),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_633),
.B(n_582),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_731),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_644),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_719),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_623),
.B(n_613),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_727),
.A2(n_575),
.B1(n_599),
.B2(n_609),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_721),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_771),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_642),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_623),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_646),
.B(n_649),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_704),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_711),
.B(n_598),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_645),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_724),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_648),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_652),
.Y(n_937)
);

AO22x1_ASAP7_75t_L g938 ( 
.A1(n_767),
.A2(n_611),
.B1(n_610),
.B2(n_598),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_615),
.A2(n_465),
.B1(n_595),
.B2(n_598),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_725),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_776),
.B(n_570),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_646),
.B(n_649),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_728),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_658),
.B(n_595),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_761),
.A2(n_611),
.B(n_610),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_665),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_621),
.A2(n_602),
.B1(n_465),
.B2(n_598),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_782),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_785),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_743),
.B(n_607),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_784),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_658),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_776),
.B(n_570),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_663),
.B(n_595),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_776),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_776),
.B(n_595),
.Y(n_956)
);

BUFx4f_ASAP7_75t_L g957 ( 
.A(n_663),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_784),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_780),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_786),
.B(n_667),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_637),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_669),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_SL g963 ( 
.A1(n_635),
.A2(n_5),
.B1(n_11),
.B2(n_14),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_733),
.B(n_492),
.Y(n_964)
);

AND2x4_ASAP7_75t_SL g965 ( 
.A(n_755),
.B(n_475),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_673),
.A2(n_475),
.B(n_479),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_672),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_744),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_674),
.B(n_465),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_703),
.B(n_607),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_675),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_679),
.B(n_602),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_706),
.A2(n_602),
.B1(n_607),
.B2(n_517),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_680),
.B(n_592),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_682),
.B(n_592),
.Y(n_975)
);

BUFx8_ASAP7_75t_L g976 ( 
.A(n_778),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_692),
.B(n_592),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_637),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_762),
.B(n_517),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_909),
.A2(n_762),
.B1(n_706),
.B2(n_714),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_833),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_849),
.A2(n_779),
.B(n_714),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_961),
.A2(n_779),
.B(n_621),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_900),
.B(n_740),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_852),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_SL g986 ( 
.A(n_909),
.B(n_770),
.C(n_740),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_961),
.A2(n_729),
.B(n_773),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_819),
.A2(n_729),
.B1(n_764),
.B2(n_752),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_865),
.A2(n_748),
.B(n_757),
.C(n_768),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_876),
.B(n_764),
.Y(n_990)
);

NOR2x1_ASAP7_75t_SL g991 ( 
.A(n_804),
.B(n_775),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_900),
.B(n_772),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_833),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_865),
.A2(n_766),
.B1(n_765),
.B2(n_592),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_854),
.B(n_592),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_801),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_859),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_876),
.A2(n_570),
.B1(n_492),
.B2(n_470),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_SL g999 ( 
.A1(n_812),
.A2(n_5),
.B1(n_15),
.B2(n_17),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_960),
.A2(n_517),
.B(n_479),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_807),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_SL g1002 ( 
.A1(n_896),
.A2(n_517),
.B(n_479),
.C(n_475),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_822),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_870),
.B(n_570),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_869),
.B(n_570),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_832),
.B(n_492),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_792),
.A2(n_492),
.B(n_470),
.C(n_22),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_852),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_967),
.B(n_492),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_863),
.B(n_15),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_849),
.A2(n_479),
.B(n_475),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_SL g1012 ( 
.A(n_932),
.B(n_18),
.C(n_22),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_863),
.B(n_18),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_866),
.B(n_959),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_804),
.A2(n_470),
.B(n_147),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_915),
.A2(n_470),
.B(n_144),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_804),
.A2(n_142),
.B(n_117),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_838),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_792),
.A2(n_894),
.B(n_789),
.C(n_790),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_831),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_795),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_788),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_866),
.B(n_116),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_957),
.B(n_104),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_906),
.A2(n_71),
.B(n_84),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_957),
.B(n_85),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_820),
.B(n_23),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_894),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_804),
.A2(n_955),
.B(n_878),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_831),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_959),
.B(n_80),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_794),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_SL g1033 ( 
.A1(n_922),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_796),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_931),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_824),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_813),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_955),
.A2(n_76),
.B(n_67),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_827),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_813),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_846),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_930),
.A2(n_65),
.B1(n_60),
.B2(n_34),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_SL g1043 ( 
.A(n_803),
.B(n_30),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_942),
.A2(n_958),
.B(n_952),
.C(n_951),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_820),
.B(n_32),
.Y(n_1045)
);

OA22x2_ASAP7_75t_L g1046 ( 
.A1(n_922),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_955),
.A2(n_41),
.B(n_42),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_787),
.B(n_42),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_860),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_826),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_835),
.B(n_43),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_963),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_951),
.A2(n_44),
.B(n_45),
.C(n_50),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_955),
.A2(n_874),
.B(n_966),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_873),
.B(n_868),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_797),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_930),
.A2(n_830),
.B1(n_793),
.B2(n_883),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_875),
.B(n_883),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_873),
.B(n_879),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_949),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_808),
.B(n_889),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_934),
.B(n_936),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_937),
.B(n_946),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_828),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_L g1065 ( 
.A(n_890),
.B(n_949),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_966),
.A2(n_898),
.B(n_892),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_799),
.Y(n_1067)
);

AO21x1_ASAP7_75t_L g1068 ( 
.A1(n_908),
.A2(n_896),
.B(n_979),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_809),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_791),
.B(n_914),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_889),
.B(n_831),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_968),
.B(n_828),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_R g1073 ( 
.A(n_850),
.B(n_882),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_825),
.B(n_888),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_880),
.A2(n_948),
.B(n_814),
.C(n_899),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_810),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_938),
.A2(n_945),
.B(n_953),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_816),
.B(n_798),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_SL g1079 ( 
.A(n_877),
.B(n_976),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_903),
.A2(n_974),
.B(n_975),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_976),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_798),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_811),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_924),
.B(n_927),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_857),
.A2(n_808),
.B(n_853),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_979),
.A2(n_818),
.B1(n_805),
.B2(n_817),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_847),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_943),
.B(n_814),
.Y(n_1088)
);

BUFx4f_ASAP7_75t_L g1089 ( 
.A(n_842),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_898),
.A2(n_941),
.B(n_895),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_948),
.A2(n_899),
.B(n_845),
.C(n_935),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_904),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_842),
.B(n_911),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_844),
.A2(n_977),
.B(n_972),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_842),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_885),
.A2(n_964),
.B(n_969),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_800),
.A2(n_920),
.B(n_978),
.C(n_933),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_929),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_935),
.B(n_962),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_855),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_911),
.B(n_817),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_841),
.B(n_940),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_962),
.B(n_971),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_890),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_933),
.A2(n_920),
.B(n_851),
.C(n_856),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_893),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_806),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_888),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_890),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_962),
.B(n_971),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_861),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_950),
.A2(n_902),
.B(n_802),
.C(n_970),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_834),
.A2(n_903),
.B(n_944),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_881),
.B(n_919),
.Y(n_1114)
);

CKINVDCx14_ASAP7_75t_R g1115 ( 
.A(n_825),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_862),
.B(n_917),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_971),
.B(n_815),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_867),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_949),
.B(n_890),
.Y(n_1119)
);

AOI222xp33_ASAP7_75t_L g1120 ( 
.A1(n_802),
.A2(n_858),
.B1(n_919),
.B2(n_872),
.C1(n_821),
.C2(n_839),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_897),
.A2(n_947),
.B(n_884),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_886),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_825),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_901),
.B(n_905),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_925),
.A2(n_843),
.B1(n_897),
.B2(n_851),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_881),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_963),
.A2(n_856),
.B(n_926),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_887),
.B(n_826),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_829),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_907),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_918),
.B(n_928),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_954),
.A2(n_848),
.B(n_891),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_912),
.B(n_923),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_916),
.B(n_921),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_1105),
.A2(n_871),
.B(n_910),
.C(n_913),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1018),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_SL g1137 ( 
.A(n_997),
.B(n_829),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_SL g1138 ( 
.A1(n_1019),
.A2(n_926),
.B(n_973),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1075),
.A2(n_925),
.B(n_837),
.C(n_850),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1011),
.A2(n_836),
.B(n_837),
.Y(n_1140)
);

AOI221x1_ASAP7_75t_L g1141 ( 
.A1(n_1127),
.A2(n_1007),
.B1(n_986),
.B2(n_1112),
.C(n_1125),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1037),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_1068),
.A2(n_864),
.A3(n_836),
.B(n_925),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1086),
.A2(n_864),
.A3(n_840),
.B(n_823),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_1097),
.A2(n_840),
.A3(n_823),
.B(n_939),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_SL g1146 ( 
.A1(n_1091),
.A2(n_823),
.B(n_956),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1113),
.A2(n_823),
.A3(n_956),
.B(n_965),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_996),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1113),
.A2(n_887),
.B(n_823),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1001),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1088),
.A2(n_882),
.B1(n_956),
.B2(n_1084),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1080),
.A2(n_956),
.B(n_1096),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1066),
.A2(n_956),
.B(n_1054),
.Y(n_1153)
);

BUFx8_ASAP7_75t_L g1154 ( 
.A(n_1100),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_980),
.B(n_1044),
.C(n_1070),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1094),
.A2(n_984),
.B(n_988),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_1049),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1088),
.B(n_1084),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1014),
.B(n_1078),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_984),
.A2(n_992),
.B(n_1121),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1021),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1003),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1099),
.B(n_1014),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_992),
.A2(n_1000),
.B(n_989),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1000),
.A2(n_1065),
.B(n_1006),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1099),
.B(n_1062),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1052),
.A2(n_1046),
.B1(n_1063),
.B2(n_1062),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1040),
.B(n_1064),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1063),
.B(n_1072),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1058),
.B(n_1126),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_982),
.A2(n_1077),
.B(n_1090),
.Y(n_1171)
);

AO21x2_ASAP7_75t_L g1172 ( 
.A1(n_1132),
.A2(n_1016),
.B(n_1002),
.Y(n_1172)
);

BUFx4f_ASAP7_75t_SL g1173 ( 
.A(n_1129),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_981),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_987),
.A2(n_1029),
.B(n_983),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1016),
.A2(n_1057),
.A3(n_1006),
.B(n_991),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_1082),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1022),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1005),
.B(n_1103),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1009),
.A2(n_995),
.B(n_1004),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_1109),
.B(n_985),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_993),
.B(n_1061),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1046),
.A2(n_990),
.B1(n_1051),
.B2(n_1076),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1035),
.A2(n_1053),
.B(n_1028),
.C(n_1107),
.Y(n_1184)
);

NAND2x1p5_ASAP7_75t_L g1185 ( 
.A(n_1089),
.B(n_1060),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_R g1186 ( 
.A(n_1055),
.B(n_1061),
.Y(n_1186)
);

AND3x4_ASAP7_75t_L g1187 ( 
.A(n_1012),
.B(n_1059),
.C(n_1116),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1051),
.B(n_1102),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_998),
.A2(n_1025),
.A3(n_1009),
.B(n_995),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1089),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1004),
.A2(n_994),
.B(n_1025),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1042),
.A2(n_1031),
.A3(n_1124),
.B(n_1134),
.Y(n_1192)
);

O2A1O1Ixp5_ASAP7_75t_L g1193 ( 
.A1(n_1031),
.A2(n_1026),
.B(n_1024),
.C(n_1101),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1109),
.A2(n_1120),
.B(n_1085),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1074),
.B(n_1059),
.Y(n_1195)
);

NAND2x1_ASAP7_75t_L g1196 ( 
.A(n_1060),
.B(n_1074),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1098),
.A2(n_1045),
.B(n_1048),
.C(n_1093),
.Y(n_1197)
);

CKINVDCx6p67_ASAP7_75t_R g1198 ( 
.A(n_1081),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_R g1199 ( 
.A(n_1114),
.B(n_1073),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1023),
.A2(n_1117),
.A3(n_1122),
.B(n_1047),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1036),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1110),
.B(n_1130),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1039),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1109),
.A2(n_1128),
.B(n_1119),
.Y(n_1205)
);

NAND2x1_ASAP7_75t_L g1206 ( 
.A(n_1074),
.B(n_1050),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1032),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1015),
.A2(n_1133),
.B(n_1005),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_1023),
.B(n_1017),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1108),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1027),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1104),
.A2(n_1123),
.B(n_1071),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1033),
.A2(n_1041),
.B(n_1118),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1020),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1034),
.B(n_1083),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1056),
.B(n_1069),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1038),
.A2(n_1087),
.B(n_1111),
.Y(n_1217)
);

AO32x2_ASAP7_75t_L g1218 ( 
.A1(n_999),
.A2(n_1115),
.A3(n_1092),
.B1(n_1067),
.B2(n_1123),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1131),
.A2(n_1050),
.B(n_1008),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1020),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1109),
.A2(n_1106),
.B(n_1008),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1020),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1123),
.A2(n_985),
.B1(n_1108),
.B2(n_1095),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1030),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1108),
.A2(n_1043),
.B(n_1030),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1030),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1095),
.B(n_1079),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1095),
.Y(n_1228)
);

OAI22x1_ASAP7_75t_L g1229 ( 
.A1(n_1070),
.A2(n_489),
.B1(n_1126),
.B2(n_1100),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1088),
.B(n_869),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1100),
.B(n_869),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1100),
.B(n_869),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1066),
.A2(n_955),
.B(n_804),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_996),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1018),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1018),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1060),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1061),
.B(n_1074),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1079),
.B(n_693),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1014),
.B(n_496),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1088),
.B(n_900),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1070),
.B(n_722),
.Y(n_1244)
);

BUFx4_ASAP7_75t_SL g1245 ( 
.A(n_1081),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1088),
.B(n_900),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1089),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1066),
.A2(n_955),
.B(n_804),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1037),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1066),
.A2(n_955),
.B(n_804),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1018),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1097),
.A2(n_1112),
.B(n_988),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1088),
.B(n_869),
.Y(n_1255)
);

O2A1O1Ixp5_ASAP7_75t_L g1256 ( 
.A1(n_1068),
.A2(n_654),
.B(n_957),
.C(n_819),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_SL g1257 ( 
.A1(n_984),
.A2(n_1051),
.B(n_1031),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1127),
.A2(n_819),
.B(n_654),
.C(n_909),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1019),
.B(n_654),
.C(n_909),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1061),
.B(n_1074),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1261)
);

NAND3x1_ASAP7_75t_L g1262 ( 
.A(n_1070),
.B(n_489),
.C(n_676),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1066),
.A2(n_955),
.B(n_804),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1097),
.A2(n_1112),
.B(n_988),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1018),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1100),
.B(n_869),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1088),
.B(n_900),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1088),
.B(n_900),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1270)
);

BUFx8_ASAP7_75t_L g1271 ( 
.A(n_996),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1011),
.A2(n_945),
.B(n_903),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1088),
.B(n_869),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1064),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1066),
.A2(n_955),
.B(n_804),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1018),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_997),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1089),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_R g1279 ( 
.A(n_997),
.B(n_433),
.Y(n_1279)
);

AOI221x1_ASAP7_75t_L g1280 ( 
.A1(n_1127),
.A2(n_1007),
.B1(n_865),
.B2(n_986),
.C(n_819),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1037),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_L g1282 ( 
.A(n_1060),
.B(n_687),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_L g1283 ( 
.A1(n_1127),
.A2(n_1007),
.B1(n_865),
.B2(n_986),
.C(n_819),
.Y(n_1283)
);

AOI221x1_ASAP7_75t_L g1284 ( 
.A1(n_1127),
.A2(n_1007),
.B1(n_865),
.B2(n_986),
.C(n_819),
.Y(n_1284)
);

O2A1O1Ixp5_ASAP7_75t_L g1285 ( 
.A1(n_1068),
.A2(n_654),
.B(n_957),
.C(n_819),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1066),
.A2(n_955),
.B(n_804),
.Y(n_1286)
);

O2A1O1Ixp5_ASAP7_75t_L g1287 ( 
.A1(n_1068),
.A2(n_654),
.B(n_957),
.C(n_819),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1259),
.A2(n_1158),
.B1(n_1230),
.B2(n_1255),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1190),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1215),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1258),
.A2(n_1259),
.B(n_1253),
.C(n_1265),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1169),
.B(n_1163),
.Y(n_1293)
);

OR2x2_ASAP7_75t_SL g1294 ( 
.A(n_1241),
.B(n_1227),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1137),
.B(n_1196),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1155),
.A2(n_1265),
.B1(n_1253),
.B2(n_1167),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1157),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1254),
.A2(n_1264),
.B(n_1261),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1216),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1141),
.A2(n_1164),
.B(n_1280),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1161),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1156),
.A2(n_1160),
.B(n_1243),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1236),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1244),
.A2(n_1170),
.B1(n_1262),
.B2(n_1243),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1271),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1155),
.A2(n_1167),
.B1(n_1183),
.B2(n_1229),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1270),
.A2(n_1272),
.B(n_1153),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1187),
.A2(n_1240),
.B1(n_1199),
.B2(n_1282),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1138),
.A2(n_1165),
.B(n_1172),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1271),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1276),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1190),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1171),
.A2(n_1233),
.B(n_1286),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1249),
.A2(n_1275),
.B(n_1263),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1283),
.A2(n_1284),
.B(n_1191),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1197),
.A2(n_1184),
.B(n_1285),
.C(n_1287),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1251),
.A2(n_1140),
.B(n_1175),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1208),
.A2(n_1257),
.B(n_1209),
.Y(n_1318)
);

AOI222xp33_ASAP7_75t_L g1319 ( 
.A1(n_1273),
.A2(n_1232),
.B1(n_1231),
.B2(n_1267),
.C1(n_1183),
.C2(n_1211),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1194),
.A2(n_1256),
.B(n_1246),
.C(n_1269),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1166),
.B(n_1188),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1250),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1136),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1178),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1180),
.A2(n_1213),
.B(n_1151),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1207),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1235),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1193),
.A2(n_1268),
.B(n_1139),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1252),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1198),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1213),
.A2(n_1151),
.B(n_1217),
.Y(n_1331)
);

CKINVDCx12_ASAP7_75t_R g1332 ( 
.A(n_1168),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1172),
.A2(n_1146),
.B(n_1135),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1266),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1190),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1152),
.A2(n_1149),
.B(n_1219),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1179),
.A2(n_1223),
.A3(n_1143),
.B(n_1205),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1150),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1179),
.A2(n_1202),
.B(n_1221),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1234),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1152),
.A2(n_1149),
.B(n_1223),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1142),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1203),
.A2(n_1159),
.B1(n_1174),
.B2(n_1201),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1174),
.A2(n_1204),
.B1(n_1162),
.B2(n_1195),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1182),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1206),
.A2(n_1225),
.B(n_1212),
.Y(n_1346)
);

AO32x2_ASAP7_75t_L g1347 ( 
.A1(n_1218),
.A2(n_1143),
.A3(n_1192),
.B1(n_1274),
.B2(n_1200),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1248),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1181),
.A2(n_1238),
.B(n_1226),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1250),
.B(n_1281),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1281),
.B(n_1148),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1279),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1143),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1177),
.B(n_1186),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1240),
.A2(n_1218),
.B1(n_1278),
.B2(n_1248),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1238),
.B(n_1181),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1154),
.A2(n_1277),
.B1(n_1173),
.B2(n_1248),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1154),
.A2(n_1277),
.B1(n_1218),
.B2(n_1210),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1189),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1147),
.A2(n_1176),
.B(n_1144),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1220),
.A2(n_1185),
.B1(n_1278),
.B2(n_1228),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1189),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1214),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1278),
.A2(n_1210),
.B1(n_1224),
.B2(n_1222),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1147),
.A2(n_1176),
.B(n_1189),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1214),
.A2(n_1224),
.B1(n_1222),
.B2(n_1192),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1214),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1147),
.A2(n_1176),
.B(n_1145),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1145),
.A2(n_1144),
.B(n_1200),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1222),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1224),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1192),
.A2(n_1242),
.B(n_1237),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1245),
.A2(n_654),
.B(n_1259),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1259),
.A2(n_1043),
.B1(n_1046),
.B2(n_865),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1190),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1244),
.B(n_686),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1215),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1215),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1259),
.A2(n_654),
.B(n_1258),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1259),
.A2(n_654),
.B(n_1258),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1215),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1259),
.A2(n_654),
.B(n_1258),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1280),
.A2(n_1068),
.A3(n_1284),
.B(n_1283),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1279),
.Y(n_1384)
);

BUFx2_ASAP7_75t_R g1385 ( 
.A(n_1220),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1386)
);

BUFx2_ASAP7_75t_R g1387 ( 
.A(n_1220),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1158),
.B(n_1169),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1194),
.A2(n_1011),
.B(n_1233),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1215),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_L g1392 ( 
.A(n_1190),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1239),
.B(n_1260),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1259),
.A2(n_654),
.B(n_1258),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1215),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1259),
.A2(n_909),
.B1(n_865),
.B2(n_1052),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1158),
.B(n_1169),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1258),
.A2(n_1105),
.B(n_819),
.C(n_1007),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1190),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1250),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1259),
.A2(n_654),
.B(n_1258),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1141),
.A2(n_1164),
.B(n_1280),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1141),
.A2(n_1164),
.B(n_1280),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1236),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1237),
.A2(n_1247),
.B(n_1242),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1258),
.A2(n_1127),
.B(n_1259),
.C(n_819),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1137),
.B(n_1109),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1215),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1259),
.A2(n_654),
.B(n_1258),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1215),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1244),
.A2(n_909),
.B1(n_1158),
.B2(n_1070),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1156),
.A2(n_900),
.B(n_1164),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1323),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1292),
.A2(n_1380),
.B(n_1379),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1333),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1347),
.B(n_1296),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1323),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1392),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1376),
.A2(n_1400),
.B1(n_1296),
.B2(n_1306),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1321),
.B(n_1293),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1302),
.A2(n_1416),
.B(n_1292),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1327),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1415),
.A2(n_1304),
.B(n_1373),
.C(n_1394),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1327),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1389),
.B(n_1401),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1347),
.B(n_1306),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1347),
.B(n_1337),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1347),
.B(n_1337),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1329),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1392),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1376),
.A2(n_1400),
.B1(n_1294),
.B2(n_1308),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1337),
.B(n_1328),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1343),
.B(n_1290),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1382),
.A2(n_1405),
.B(n_1413),
.C(n_1410),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1365),
.A2(n_1372),
.B(n_1318),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1354),
.A2(n_1343),
.B1(n_1358),
.B2(n_1374),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1318),
.A2(n_1360),
.B(n_1368),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1337),
.B(n_1353),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1353),
.B(n_1358),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1324),
.Y(n_1444)
);

O2A1O1Ixp5_ASAP7_75t_L g1445 ( 
.A1(n_1288),
.A2(n_1374),
.B(n_1320),
.C(n_1339),
.Y(n_1445)
);

AOI211xp5_ASAP7_75t_L g1446 ( 
.A1(n_1288),
.A2(n_1355),
.B(n_1316),
.C(n_1402),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1340),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1300),
.A2(n_1406),
.B(n_1407),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_L g1449 ( 
.A(n_1384),
.B(n_1301),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1334),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1320),
.A2(n_1414),
.B(n_1412),
.C(n_1377),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_SL g1452 ( 
.A1(n_1393),
.A2(n_1355),
.B(n_1387),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1299),
.B(n_1378),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1402),
.A2(n_1354),
.B(n_1381),
.C(n_1391),
.Y(n_1454)
);

AOI21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1393),
.A2(n_1385),
.B(n_1295),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1396),
.B(n_1345),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1368),
.A2(n_1314),
.B(n_1397),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1344),
.A2(n_1404),
.B1(n_1322),
.B2(n_1351),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1314),
.A2(n_1388),
.B(n_1399),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1408),
.B(n_1369),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1319),
.B(n_1351),
.Y(n_1461)
);

O2A1O1Ixp5_ASAP7_75t_L g1462 ( 
.A1(n_1390),
.A2(n_1362),
.B(n_1359),
.C(n_1364),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1346),
.A2(n_1366),
.B(n_1344),
.C(n_1311),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1303),
.A2(n_1407),
.B(n_1406),
.C(n_1300),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1386),
.A2(n_1397),
.B(n_1398),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1338),
.B(n_1370),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1363),
.B(n_1289),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1384),
.A2(n_1411),
.B(n_1357),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1300),
.A2(n_1406),
.B(n_1310),
.C(n_1305),
.Y(n_1469)
);

O2A1O1Ixp5_ASAP7_75t_L g1470 ( 
.A1(n_1289),
.A2(n_1312),
.B(n_1403),
.C(n_1375),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1315),
.A2(n_1309),
.B(n_1313),
.Y(n_1471)
);

OAI31xp33_ASAP7_75t_L g1472 ( 
.A1(n_1361),
.A2(n_1411),
.A3(n_1312),
.B(n_1375),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_L g1473 ( 
.A(n_1403),
.B(n_1367),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1367),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1332),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1352),
.A2(n_1366),
.B1(n_1335),
.B2(n_1330),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1356),
.A2(n_1348),
.B(n_1315),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1349),
.B(n_1371),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1348),
.B(n_1383),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1356),
.A2(n_1348),
.B(n_1315),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1352),
.A2(n_1335),
.B1(n_1330),
.B2(n_1348),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1383),
.B(n_1325),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1383),
.B(n_1325),
.Y(n_1483)
);

AOI221x1_ASAP7_75t_SL g1484 ( 
.A1(n_1297),
.A2(n_1335),
.B1(n_1325),
.B2(n_1331),
.C(n_1341),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1336),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1331),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1297),
.B(n_1331),
.Y(n_1487)
);

OA22x2_ASAP7_75t_L g1488 ( 
.A1(n_1317),
.A2(n_1307),
.B1(n_1298),
.B2(n_1291),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1317),
.B(n_1307),
.Y(n_1489)
);

CKINVDCx6p67_ASAP7_75t_R g1490 ( 
.A(n_1386),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1388),
.A2(n_1395),
.B1(n_1398),
.B2(n_1399),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1395),
.A2(n_1365),
.B(n_1416),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1409),
.B(n_1323),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1323),
.B(n_1326),
.Y(n_1494)
);

AND2x2_ASAP7_75t_SL g1495 ( 
.A(n_1296),
.B(n_1306),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1323),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1347),
.B(n_1296),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1376),
.A2(n_909),
.B1(n_1400),
.B2(n_1296),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1323),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1294),
.B(n_1345),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1415),
.A2(n_1258),
.B(n_1304),
.C(n_722),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1376),
.A2(n_909),
.B1(n_1400),
.B2(n_1296),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1323),
.B(n_1326),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1323),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1350),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1342),
.Y(n_1506)
);

AOI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1415),
.A2(n_909),
.B1(n_1296),
.B2(n_865),
.C(n_1288),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1505),
.B(n_1438),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1493),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1471),
.A2(n_1448),
.B(n_1425),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1486),
.A2(n_1445),
.B(n_1462),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1483),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1485),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1423),
.B(n_1498),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1460),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1483),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1442),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1438),
.B(n_1437),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1465),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1436),
.B(n_1430),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1436),
.B(n_1430),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1490),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1420),
.B(n_1497),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1465),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1424),
.B(n_1433),
.Y(n_1525)
);

INVx4_ASAP7_75t_L g1526 ( 
.A(n_1478),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1420),
.B(n_1497),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1507),
.A2(n_1501),
.B(n_1451),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1418),
.A2(n_1491),
.B(n_1464),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1463),
.A2(n_1451),
.B(n_1469),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1488),
.A2(n_1419),
.B(n_1457),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1489),
.B(n_1427),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1504),
.B(n_1429),
.Y(n_1534)
);

OAI31xp33_ASAP7_75t_L g1535 ( 
.A1(n_1502),
.A2(n_1435),
.A3(n_1440),
.B(n_1461),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1489),
.B(n_1463),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1495),
.B(n_1444),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1479),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1417),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1421),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1431),
.A2(n_1432),
.B(n_1487),
.Y(n_1541)
);

AOI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1488),
.A2(n_1439),
.B(n_1459),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1441),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1494),
.B(n_1503),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1446),
.B(n_1495),
.C(n_1454),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1450),
.B(n_1503),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1428),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1496),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1499),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1517),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1519),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1513),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1547),
.B(n_1439),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1508),
.B(n_1503),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1519),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1528),
.A2(n_1453),
.B(n_1492),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1426),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1519),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1512),
.B(n_1457),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1517),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1510),
.A2(n_1443),
.B(n_1476),
.Y(n_1563)
);

NAND4xp25_ASAP7_75t_L g1564 ( 
.A(n_1535),
.B(n_1458),
.C(n_1472),
.D(n_1500),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1541),
.B(n_1457),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1509),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1541),
.B(n_1492),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1519),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1516),
.B(n_1459),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1516),
.B(n_1459),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1524),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1516),
.B(n_1426),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1552),
.Y(n_1574)
);

OAI211xp5_ASAP7_75t_L g1575 ( 
.A1(n_1564),
.A2(n_1535),
.B(n_1545),
.C(n_1514),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1564),
.A2(n_1514),
.B1(n_1545),
.B2(n_1533),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1564),
.A2(n_1533),
.B1(n_1518),
.B2(n_1537),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1569),
.B(n_1571),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1556),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1563),
.A2(n_1533),
.B1(n_1518),
.B2(n_1537),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1567),
.A2(n_1532),
.B(n_1543),
.Y(n_1581)
);

A2O1A1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1558),
.A2(n_1449),
.B(n_1522),
.C(n_1481),
.Y(n_1582)
);

OAI31xp33_ASAP7_75t_L g1583 ( 
.A1(n_1554),
.A2(n_1475),
.A3(n_1447),
.B(n_1506),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1553),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1554),
.A2(n_1546),
.B1(n_1534),
.B2(n_1525),
.C(n_1531),
.Y(n_1585)
);

NAND5xp2_ASAP7_75t_L g1586 ( 
.A(n_1558),
.B(n_1468),
.C(n_1452),
.D(n_1455),
.E(n_1456),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1552),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1556),
.B(n_1520),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_SL g1589 ( 
.A(n_1563),
.B(n_1531),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1551),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1559),
.A2(n_1533),
.B1(n_1530),
.B2(n_1536),
.Y(n_1591)
);

AND4x1_ASAP7_75t_L g1592 ( 
.A(n_1563),
.B(n_1470),
.C(n_1467),
.D(n_1466),
.Y(n_1592)
);

AOI33xp33_ASAP7_75t_L g1593 ( 
.A1(n_1555),
.A2(n_1515),
.A3(n_1540),
.B1(n_1539),
.B2(n_1548),
.B3(n_1550),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1566),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1567),
.B(n_1534),
.C(n_1525),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1569),
.B(n_1541),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1553),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1569),
.B(n_1541),
.Y(n_1599)
);

OAI211xp5_ASAP7_75t_L g1600 ( 
.A1(n_1567),
.A2(n_1538),
.B(n_1511),
.C(n_1549),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1563),
.A2(n_1542),
.B(n_1543),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1559),
.B(n_1474),
.Y(n_1602)
);

INVx5_ASAP7_75t_L g1603 ( 
.A(n_1570),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1551),
.B(n_1541),
.Y(n_1604)
);

NAND4xp25_ASAP7_75t_SL g1605 ( 
.A(n_1565),
.B(n_1521),
.C(n_1520),
.D(n_1523),
.Y(n_1605)
);

OAI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1570),
.A2(n_1533),
.B(n_1536),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1570),
.A2(n_1533),
.B1(n_1531),
.B2(n_1536),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1570),
.A2(n_1531),
.B1(n_1536),
.B2(n_1529),
.Y(n_1608)
);

NAND4xp25_ASAP7_75t_SL g1609 ( 
.A(n_1565),
.B(n_1521),
.C(n_1523),
.D(n_1527),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1544),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1562),
.A2(n_1522),
.B(n_1422),
.C(n_1434),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1584),
.Y(n_1612)
);

AOI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1592),
.A2(n_1568),
.B(n_1572),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1581),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1603),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1603),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1584),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1594),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

NOR2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1579),
.B(n_1474),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1604),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1606),
.B(n_1530),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1598),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1598),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1600),
.A2(n_1532),
.B(n_1543),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_SL g1627 ( 
.A(n_1604),
.B(n_1530),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1593),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1589),
.A2(n_1582),
.B(n_1586),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1574),
.Y(n_1630)
);

AOI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1592),
.A2(n_1560),
.B(n_1557),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1587),
.Y(n_1632)
);

CKINVDCx16_ASAP7_75t_R g1633 ( 
.A(n_1591),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1601),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1585),
.B(n_1526),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1628),
.B(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1617),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1617),
.Y(n_1639)
);

NOR2xp67_ASAP7_75t_L g1640 ( 
.A(n_1615),
.B(n_1605),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1628),
.B(n_1596),
.Y(n_1641)
);

OAI211xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1629),
.A2(n_1575),
.B(n_1583),
.C(n_1576),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1621),
.B(n_1597),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1621),
.B(n_1599),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1620),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1635),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1615),
.B(n_1616),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1629),
.A2(n_1635),
.B1(n_1633),
.B2(n_1580),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1620),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1618),
.B(n_1599),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1625),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1625),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1612),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1616),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1612),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1618),
.B(n_1622),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1633),
.B(n_1583),
.C(n_1577),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1623),
.A2(n_1606),
.B1(n_1586),
.B2(n_1607),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1627),
.B(n_1578),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1619),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1627),
.B(n_1578),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1616),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_1603),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1603),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1615),
.B(n_1611),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1615),
.B(n_1603),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1623),
.B(n_1603),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1615),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1619),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1614),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1622),
.B(n_1588),
.Y(n_1672)
);

OAI31xp33_ASAP7_75t_L g1673 ( 
.A1(n_1613),
.A2(n_1591),
.A3(n_1608),
.B(n_1609),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_R g1674 ( 
.A(n_1623),
.B(n_1530),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1623),
.B(n_1569),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1571),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1613),
.B(n_1588),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1631),
.B(n_1571),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1624),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1646),
.B(n_1602),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1653),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1654),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1642),
.B(n_1610),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1641),
.B(n_1631),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1643),
.B(n_1631),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1654),
.B(n_1662),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1648),
.A2(n_1536),
.B1(n_1626),
.B2(n_1636),
.C(n_1634),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1641),
.B(n_1624),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1643),
.B(n_1595),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1660),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1644),
.B(n_1640),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.B(n_1595),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1670),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1670),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1640),
.B(n_1595),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1665),
.B(n_1595),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1654),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1638),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1638),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1669),
.B(n_1632),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1637),
.B(n_1571),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1647),
.Y(n_1709)
);

INVxp33_ASAP7_75t_L g1710 ( 
.A(n_1657),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1639),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_L g1712 ( 
.A(n_1657),
.B(n_1636),
.C(n_1634),
.D(n_1422),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1637),
.B(n_1561),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1639),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1645),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1695),
.B(n_1647),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1693),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1695),
.B(n_1709),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.B(n_1647),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1647),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

CKINVDCx16_ASAP7_75t_R g1722 ( 
.A(n_1710),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1693),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1683),
.B(n_1659),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1710),
.A2(n_1658),
.B1(n_1668),
.B2(n_1677),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1694),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1683),
.B(n_1659),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1684),
.B(n_1666),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_L g1729 ( 
.A(n_1712),
.B(n_1669),
.C(n_1662),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1703),
.B(n_1661),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1691),
.B(n_1650),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1703),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1694),
.Y(n_1733)
);

NAND2x1p5_ASAP7_75t_L g1734 ( 
.A(n_1707),
.B(n_1669),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1702),
.B(n_1669),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1661),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1663),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1691),
.B(n_1650),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1690),
.A2(n_1663),
.B1(n_1664),
.B2(n_1667),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1681),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1722),
.B(n_1680),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1716),
.B(n_1701),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1725),
.A2(n_1673),
.B1(n_1687),
.B2(n_1674),
.C(n_1711),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1729),
.A2(n_1673),
.B1(n_1705),
.B2(n_1664),
.C(n_1667),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1734),
.Y(n_1745)
);

AOI21xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1722),
.A2(n_1714),
.B(n_1704),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1716),
.B(n_1701),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1719),
.Y(n_1748)
);

OAI332xp33_ASAP7_75t_L g1749 ( 
.A1(n_1732),
.A2(n_1715),
.A3(n_1714),
.B1(n_1704),
.B2(n_1682),
.B3(n_1686),
.C1(n_1698),
.C2(n_1685),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1728),
.A2(n_1715),
.B1(n_1688),
.B2(n_1702),
.C(n_1699),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1718),
.B(n_1688),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1692),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1739),
.A2(n_1713),
.B1(n_1708),
.B2(n_1696),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1734),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1692),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1720),
.B(n_1679),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1717),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1696),
.Y(n_1758)
);

NAND2x1_ASAP7_75t_SL g1759 ( 
.A(n_1735),
.B(n_1678),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1757),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1741),
.B(n_1721),
.Y(n_1761)
);

AND2x2_ASAP7_75t_SL g1762 ( 
.A(n_1741),
.B(n_1721),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1756),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1742),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1756),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.B(n_1724),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1746),
.B(n_1737),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1732),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1747),
.B(n_1724),
.Y(n_1769)
);

OAI222xp33_ASAP7_75t_L g1770 ( 
.A1(n_1743),
.A2(n_1734),
.B1(n_1738),
.B2(n_1731),
.C1(n_1737),
.C2(n_1727),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1744),
.B(n_1750),
.Y(n_1771)
);

AOI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1763),
.A2(n_1749),
.B1(n_1765),
.B2(n_1767),
.C(n_1761),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1762),
.B(n_1751),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1764),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1763),
.A2(n_1765),
.B1(n_1768),
.B2(n_1766),
.C(n_1769),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1762),
.A2(n_1759),
.B(n_1745),
.C(n_1754),
.Y(n_1776)
);

O2A1O1Ixp33_ASAP7_75t_L g1777 ( 
.A1(n_1760),
.A2(n_1745),
.B(n_1754),
.C(n_1740),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1766),
.A2(n_1752),
.B(n_1758),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1769),
.A2(n_1740),
.B1(n_1747),
.B2(n_1727),
.C(n_1730),
.Y(n_1779)
);

NOR4xp25_ASAP7_75t_L g1780 ( 
.A(n_1770),
.B(n_1717),
.C(n_1723),
.D(n_1726),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1772),
.A2(n_1771),
.B1(n_1778),
.B2(n_1773),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1780),
.A2(n_1753),
.B1(n_1738),
.B2(n_1731),
.C(n_1730),
.Y(n_1782)
);

AO22x2_ASAP7_75t_L g1783 ( 
.A1(n_1774),
.A2(n_1723),
.B1(n_1726),
.B2(n_1733),
.Y(n_1783)
);

XNOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1775),
.B(n_1755),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1776),
.A2(n_1777),
.B(n_1779),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1771),
.A2(n_1755),
.B1(n_1735),
.B2(n_1736),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1783),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1784),
.B(n_1735),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_SL g1789 ( 
.A(n_1785),
.B(n_1434),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1786),
.B(n_1735),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1782),
.B(n_1697),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1781),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1783),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1792),
.A2(n_1736),
.B1(n_1733),
.B2(n_1706),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1787),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1788),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_R g1797 ( 
.A(n_1793),
.B(n_1697),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1790),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1795),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1798),
.B(n_1791),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_SL g1801 ( 
.A(n_1796),
.B(n_1789),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1799),
.B(n_1796),
.Y(n_1802)
);

AOI32xp33_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1801),
.A3(n_1800),
.B1(n_1794),
.B2(n_1797),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1706),
.B1(n_1652),
.B2(n_1651),
.C(n_1649),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1805),
.Y(n_1806)
);

NAND2x1_ASAP7_75t_SL g1807 ( 
.A(n_1804),
.B(n_1645),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1806),
.B(n_1651),
.C(n_1649),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1652),
.B1(n_1679),
.B2(n_1671),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1808),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1809),
.B(n_1671),
.Y(n_1811)
);

NAND2x1p5_ASAP7_75t_L g1812 ( 
.A(n_1811),
.B(n_1473),
.Y(n_1812)
);

AO221x2_ASAP7_75t_L g1813 ( 
.A1(n_1812),
.A2(n_1671),
.B1(n_1634),
.B2(n_1636),
.C(n_1672),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1636),
.B1(n_1634),
.B2(n_1678),
.C(n_1675),
.Y(n_1814)
);

AOI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1676),
.B(n_1675),
.C(n_1614),
.Y(n_1815)
);


endmodule