module fake_jpeg_2754_n_676 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_676);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_676;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_583;
wire n_56;
wire n_240;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_60),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_11),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_62),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_63),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_65),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_22),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_27),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_89),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_106),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_19),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_18),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_28),
.B(n_10),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

BUFx12f_ASAP7_75t_SL g111 ( 
.A(n_23),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_111),
.Y(n_152)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_118),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_33),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_50),
.B(n_10),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_125),
.Y(n_177)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_23),
.Y(n_127)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_37),
.B(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_131),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_23),
.Y(n_130)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_34),
.B(n_8),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_32),
.B1(n_47),
.B2(n_53),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_139),
.A2(n_165),
.B1(n_25),
.B2(n_1),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_34),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_147),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_153),
.B(n_154),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_63),
.B(n_57),
.Y(n_154)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_157),
.Y(n_243)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_162),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_98),
.A2(n_47),
.B1(n_55),
.B2(n_53),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_34),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_65),
.B(n_37),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_169),
.B(n_170),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_68),
.A2(n_57),
.B(n_44),
.C(n_46),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_88),
.B(n_51),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_180),
.B(n_194),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_109),
.A2(n_44),
.B1(n_46),
.B2(n_51),
.Y(n_183)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_55),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_101),
.B(n_55),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_196),
.B(n_210),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_87),
.A2(n_39),
.B1(n_53),
.B2(n_55),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_203),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_270)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_204),
.Y(n_303)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_129),
.B(n_53),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_167),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_64),
.A2(n_25),
.B1(n_34),
.B2(n_39),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_117),
.B(n_39),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_212),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_102),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_107),
.B(n_12),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_66),
.B(n_12),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_223),
.Y(n_235)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_73),
.B(n_18),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_82),
.Y(n_226)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_230),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_168),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_232),
.B(n_242),
.Y(n_360)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_147),
.B(n_96),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_233),
.Y(n_317)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_152),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_236),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_1),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_237),
.B(n_239),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_132),
.B(n_1),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_241),
.B(n_301),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_25),
.B(n_2),
.C(n_3),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_156),
.B(n_95),
.C(n_93),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_247),
.B(n_164),
.C(n_186),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_168),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_248),
.B(n_268),
.Y(n_316)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_249),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_179),
.A2(n_91),
.B1(n_90),
.B2(n_86),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_250),
.A2(n_149),
.B1(n_276),
.B2(n_291),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_134),
.B(n_84),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_251),
.B(n_253),
.Y(n_321)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_134),
.B(n_83),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_141),
.B(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_259),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_159),
.Y(n_258)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_141),
.B(n_1),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_177),
.B(n_2),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_261),
.B(n_272),
.Y(n_340)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_263),
.Y(n_359)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_5),
.Y(n_265)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_265),
.B(n_218),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_133),
.A2(n_25),
.B1(n_6),
.B2(n_7),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_266),
.A2(n_287),
.B1(n_289),
.B2(n_292),
.Y(n_322)
);

BUFx4f_ASAP7_75t_SL g267 ( 
.A(n_136),
.Y(n_267)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_267),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_5),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_270),
.A2(n_139),
.B1(n_165),
.B2(n_166),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_135),
.B(n_8),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_275),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_177),
.B(n_8),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_155),
.Y(n_273)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_178),
.B(n_13),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_18),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_276),
.A2(n_151),
.B(n_202),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_190),
.B(n_13),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_278),
.B(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_180),
.B(n_206),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_281),
.B(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

CKINVDCx9p33_ASAP7_75t_R g283 ( 
.A(n_182),
.Y(n_283)
);

BUFx4f_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_175),
.Y(n_284)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_174),
.Y(n_286)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_144),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_163),
.Y(n_288)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_137),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_181),
.Y(n_290)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_137),
.A2(n_15),
.B1(n_18),
.B2(n_198),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_171),
.B(n_15),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_195),
.Y(n_294)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_150),
.A2(n_158),
.B1(n_138),
.B2(n_148),
.Y(n_296)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_185),
.B(n_187),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_297),
.B(n_184),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_155),
.Y(n_298)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_213),
.B(n_198),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_211),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_146),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_136),
.B(n_161),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_304),
.B(n_205),
.Y(n_358)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_200),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_305),
.Y(n_313)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_220),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_142),
.Y(n_350)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_164),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_307),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_136),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_308),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_245),
.A2(n_229),
.B1(n_281),
.B2(n_297),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_309),
.A2(n_311),
.B1(n_243),
.B2(n_285),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_237),
.A2(n_176),
.B1(n_201),
.B2(n_197),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_315),
.B(n_327),
.Y(n_388)
);

AO22x2_ASAP7_75t_SL g319 ( 
.A1(n_250),
.A2(n_176),
.B1(n_201),
.B2(n_197),
.Y(n_319)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_319),
.A2(n_296),
.B1(n_257),
.B2(n_231),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_324),
.A2(n_267),
.B1(n_306),
.B2(n_305),
.Y(n_389)
);

O2A1O1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_242),
.A2(n_172),
.B(n_218),
.C(n_151),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_336),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_241),
.A2(n_184),
.B1(n_192),
.B2(n_191),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_283),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_334),
.B(n_351),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_228),
.A2(n_140),
.B1(n_166),
.B2(n_143),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_339),
.B1(n_349),
.B2(n_366),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_235),
.A2(n_140),
.B1(n_143),
.B2(n_186),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_241),
.A2(n_227),
.B1(n_265),
.B2(n_246),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_265),
.A2(n_218),
.B1(n_205),
.B2(n_202),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_233),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_228),
.A2(n_191),
.B1(n_192),
.B2(n_142),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_260),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_365),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_233),
.B(n_149),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_364),
.B(n_246),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_260),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_369),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_348),
.A2(n_302),
.B1(n_235),
.B2(n_279),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_373),
.A2(n_381),
.B1(n_389),
.B2(n_406),
.Y(n_425)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_377),
.Y(n_454)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_362),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_379),
.Y(n_450)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_380),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_348),
.A2(n_276),
.B1(n_247),
.B2(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_360),
.A2(n_261),
.B(n_272),
.C(n_259),
.Y(n_384)
);

OAI31xp33_ASAP7_75t_L g438 ( 
.A1(n_384),
.A2(n_399),
.A3(n_415),
.B(n_314),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_385),
.B(n_325),
.Y(n_446)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_386),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_316),
.B(n_340),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_387),
.B(n_404),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_277),
.C(n_239),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_315),
.C(n_340),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_361),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_402),
.Y(n_419)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_392),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_366),
.A2(n_254),
.B1(n_296),
.B2(n_307),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_409),
.Y(n_424)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_395),
.Y(n_456)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_334),
.A2(n_238),
.B1(n_252),
.B2(n_231),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_397),
.A2(n_405),
.B1(n_413),
.B2(n_357),
.Y(n_445)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_308),
.B(n_267),
.Y(n_399)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_400),
.Y(n_449)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_329),
.Y(n_402)
);

CKINVDCx12_ASAP7_75t_R g404 ( 
.A(n_342),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_317),
.A2(n_276),
.B1(n_286),
.B2(n_282),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_321),
.B(n_301),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_350),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_412),
.Y(n_428)
);

AO22x1_ASAP7_75t_SL g411 ( 
.A1(n_364),
.A2(n_284),
.B1(n_257),
.B2(n_285),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_411),
.A2(n_319),
.B(n_405),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_350),
.Y(n_412)
);

INVx13_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_354),
.A2(n_269),
.B1(n_230),
.B2(n_262),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_315),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_372),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_352),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_423),
.C(n_446),
.Y(n_458)
);

OAI32xp33_ASAP7_75t_L g421 ( 
.A1(n_370),
.A2(n_352),
.A3(n_321),
.B1(n_320),
.B2(n_354),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_421),
.Y(n_467)
);

AOI22x1_ASAP7_75t_SL g422 ( 
.A1(n_370),
.A2(n_326),
.B1(n_349),
.B2(n_337),
.Y(n_422)
);

AO21x1_ASAP7_75t_L g486 ( 
.A1(n_422),
.A2(n_406),
.B(n_415),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_312),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_376),
.A2(n_328),
.B1(n_327),
.B2(n_364),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_431),
.A2(n_388),
.B1(n_416),
.B2(n_408),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_336),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_436),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_312),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_440),
.Y(n_480)
);

OAI32xp33_ASAP7_75t_L g440 ( 
.A1(n_376),
.A2(n_314),
.A3(n_325),
.B1(n_318),
.B2(n_333),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_347),
.Y(n_443)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_443),
.Y(n_461)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_378),
.A2(n_313),
.B1(n_351),
.B2(n_365),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_448),
.A2(n_453),
.B(n_455),
.Y(n_482)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_416),
.A2(n_325),
.B(n_322),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g455 ( 
.A1(n_388),
.A2(n_407),
.A3(n_373),
.B1(n_378),
.B2(n_393),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_450),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_473),
.Y(n_507)
);

INVx13_ASAP7_75t_L g459 ( 
.A(n_449),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_459),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_466),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_488),
.Y(n_496)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_463),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_464),
.A2(n_471),
.B1(n_488),
.B2(n_492),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_384),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_402),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_468),
.B(n_470),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_417),
.B(n_408),
.CI(n_399),
.CON(n_469),
.SN(n_469)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_469),
.B(n_440),
.CI(n_425),
.CON(n_504),
.SN(n_504)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_419),
.B(n_335),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_433),
.A2(n_372),
.B1(n_388),
.B2(n_412),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_369),
.C(n_410),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_472),
.B(n_494),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_439),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_435),
.B(n_375),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_477),
.Y(n_502)
);

OR2x4_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_427),
.Y(n_478)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_333),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_479),
.B(n_481),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_335),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_443),
.B(n_374),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_483),
.B(n_451),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_421),
.B(n_369),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_484),
.B(n_432),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_439),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_489),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_486),
.A2(n_453),
.B(n_429),
.Y(n_511)
);

OAI22x1_ASAP7_75t_SL g487 ( 
.A1(n_433),
.A2(n_394),
.B1(n_371),
.B2(n_411),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_487),
.A2(n_491),
.B1(n_418),
.B2(n_431),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_424),
.A2(n_394),
.B1(n_371),
.B2(n_392),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_428),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_427),
.Y(n_490)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_490),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_424),
.A2(n_394),
.B1(n_319),
.B2(n_411),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_425),
.A2(n_394),
.B1(n_319),
.B2(n_396),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_444),
.A2(n_377),
.B1(n_414),
.B2(n_331),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_493),
.A2(n_391),
.B1(n_430),
.B2(n_454),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_428),
.B(n_313),
.C(n_310),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_496),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_498),
.A2(n_457),
.B1(n_430),
.B2(n_442),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_503),
.B(n_506),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_504),
.A2(n_512),
.B(n_480),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_483),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_429),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_513),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_511),
.A2(n_522),
.B(n_526),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_447),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_461),
.B(n_377),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_514),
.B(n_525),
.C(n_531),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_462),
.A2(n_422),
.B1(n_418),
.B2(n_452),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_516),
.A2(n_487),
.B1(n_491),
.B2(n_477),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_463),
.Y(n_517)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_517),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_489),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_518),
.A2(n_527),
.B1(n_528),
.B2(n_529),
.Y(n_553)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_519),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_437),
.Y(n_521)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_521),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_482),
.A2(n_454),
.B(n_456),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_437),
.Y(n_523)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_524),
.B(n_497),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_461),
.B(n_395),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_482),
.A2(n_451),
.B(n_432),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_474),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_467),
.A2(n_456),
.B1(n_441),
.B2(n_442),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_530),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_467),
.B(n_398),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_532),
.B(n_501),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_534),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_536),
.A2(n_541),
.B1(n_548),
.B2(n_557),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_472),
.C(n_460),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_537),
.B(n_543),
.C(n_544),
.Y(n_569)
);

XNOR2x1_ASAP7_75t_SL g540 ( 
.A(n_497),
.B(n_484),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_540),
.B(n_499),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_516),
.A2(n_480),
.B1(n_465),
.B2(n_486),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_502),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_542),
.B(n_506),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_505),
.B(n_466),
.C(n_464),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_513),
.B(n_475),
.C(n_469),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_475),
.C(n_469),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_549),
.C(n_554),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_520),
.A2(n_492),
.B1(n_465),
.B2(n_476),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_503),
.B(n_490),
.C(n_478),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_551),
.A2(n_555),
.B1(n_558),
.B2(n_562),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_332),
.C(n_355),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_498),
.A2(n_527),
.B1(n_502),
.B2(n_518),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_496),
.A2(n_331),
.B1(n_426),
.B2(n_383),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_496),
.A2(n_426),
.B1(n_459),
.B2(n_386),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_332),
.C(n_355),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_560),
.B(n_563),
.C(n_363),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_310),
.B(n_401),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_561),
.A2(n_508),
.B(n_507),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_526),
.A2(n_367),
.B1(n_298),
.B2(n_273),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_355),
.C(n_359),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_547),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_572),
.Y(n_604)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_538),
.Y(n_566)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_566),
.Y(n_591)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_553),
.Y(n_568)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_582),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_533),
.B(n_507),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_573),
.A2(n_577),
.B1(n_586),
.B2(n_561),
.Y(n_598)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_555),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_574),
.B(n_575),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_539),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_556),
.A2(n_511),
.B(n_508),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_576),
.A2(n_556),
.B(n_557),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_550),
.A2(n_504),
.B1(n_517),
.B2(n_515),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_515),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_578),
.B(n_581),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_585),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_548),
.A2(n_504),
.B1(n_519),
.B2(n_495),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_580),
.A2(n_379),
.B1(n_359),
.B2(n_345),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_559),
.B(n_509),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_544),
.B(n_509),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_583),
.B(n_368),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_537),
.B(n_528),
.C(n_499),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_584),
.B(n_546),
.C(n_554),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_535),
.A2(n_500),
.B1(n_495),
.B2(n_368),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_546),
.B(n_500),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_587),
.B(n_234),
.C(n_303),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_552),
.B(n_367),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_589),
.B(n_552),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_590),
.B(n_595),
.Y(n_627)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_592),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_565),
.A2(n_558),
.B1(n_551),
.B2(n_562),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_609),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_543),
.C(n_545),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_540),
.C(n_563),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_596),
.Y(n_617)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_598),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_571),
.B(n_569),
.C(n_578),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_600),
.C(n_603),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_532),
.C(n_560),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_588),
.B(n_536),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_601),
.Y(n_615)
);

OAI21x1_ASAP7_75t_SL g621 ( 
.A1(n_602),
.A2(n_572),
.B(n_589),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_587),
.B(n_541),
.C(n_363),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_575),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_611),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_574),
.A2(n_345),
.B1(n_338),
.B2(n_356),
.Y(n_609)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_614),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g616 ( 
.A1(n_605),
.A2(n_568),
.B(n_580),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_616),
.B(n_567),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_599),
.B(n_577),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_619),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_590),
.B(n_582),
.C(n_585),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_575),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_623),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_621),
.A2(n_623),
.B(n_607),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_600),
.B(n_576),
.C(n_567),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_595),
.B(n_579),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_629),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_603),
.B(n_610),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_626),
.B(n_611),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_604),
.B(n_566),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_631),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_SL g631 ( 
.A1(n_628),
.A2(n_597),
.B(n_570),
.C(n_593),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_612),
.A2(n_610),
.B(n_594),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_635),
.A2(n_638),
.B(n_356),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_596),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_636),
.B(n_639),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_594),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_616),
.Y(n_639)
);

AOI31xp67_ASAP7_75t_L g647 ( 
.A1(n_640),
.A2(n_619),
.A3(n_622),
.B(n_625),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_641),
.B(n_642),
.Y(n_654)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_616),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_615),
.B(n_591),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_643),
.B(n_634),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_613),
.B(n_586),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_644),
.B(n_249),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_632),
.B(n_613),
.C(n_627),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_645),
.B(n_649),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_630),
.A2(n_622),
.B1(n_609),
.B2(n_626),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_646),
.B(n_648),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_647),
.A2(n_651),
.B(n_652),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_633),
.A2(n_625),
.B1(n_264),
.B2(n_263),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_637),
.B(n_338),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_655),
.A2(n_635),
.B1(n_631),
.B2(n_641),
.Y(n_659)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_659),
.Y(n_668)
);

BUFx4f_ASAP7_75t_SL g660 ( 
.A(n_647),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_660),
.A2(n_662),
.B(n_663),
.Y(n_666)
);

AOI322xp5_ASAP7_75t_L g661 ( 
.A1(n_650),
.A2(n_631),
.A3(n_380),
.B1(n_400),
.B2(n_413),
.C1(n_290),
.C2(n_256),
.Y(n_661)
);

BUFx24_ASAP7_75t_SL g667 ( 
.A(n_661),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_645),
.B(n_295),
.C(n_234),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_303),
.C(n_240),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_657),
.B(n_654),
.Y(n_664)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_664),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_658),
.C(n_659),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_665),
.B(n_660),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_669),
.B(n_671),
.C(n_668),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_666),
.B(n_646),
.Y(n_671)
);

AOI322xp5_ASAP7_75t_L g673 ( 
.A1(n_672),
.A2(n_670),
.A3(n_667),
.B1(n_649),
.B2(n_290),
.C1(n_244),
.C2(n_243),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_673),
.B(n_240),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_244),
.Y(n_675)
);

BUFx24_ASAP7_75t_SL g676 ( 
.A(n_675),
.Y(n_676)
);


endmodule