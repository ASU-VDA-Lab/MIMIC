module fake_jpeg_1332_n_534 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_52),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_14),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_6),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_60),
.Y(n_114)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_81),
.Y(n_159)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_91),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_23),
.B(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_10),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_46),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_154),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_117),
.B(n_118),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_121),
.B(n_123),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_55),
.B(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_135),
.Y(n_164)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_70),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g197 ( 
.A(n_130),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_74),
.B(n_28),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_85),
.B(n_47),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_138),
.B(n_140),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_57),
.B(n_47),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_48),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_63),
.A2(n_56),
.B1(n_32),
.B2(n_43),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_22),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_57),
.A2(n_19),
.B(n_18),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_45),
.B(n_107),
.C(n_30),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_62),
.B(n_46),
.Y(n_154)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_24),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_167),
.B(n_171),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_169),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_24),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_174),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_114),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_194),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_65),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_192),
.Y(n_238)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_126),
.A2(n_149),
.B1(n_157),
.B2(n_73),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_204),
.B1(n_27),
.B2(n_81),
.Y(n_220)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_183),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_28),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_189),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_196),
.Y(n_235)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_98),
.B1(n_97),
.B2(n_67),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_36),
.B1(n_43),
.B2(n_127),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_104),
.A2(n_58),
.B1(n_89),
.B2(n_86),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_42),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_19),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_78),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_201),
.Y(n_244)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_87),
.B1(n_83),
.B2(n_76),
.Y(n_204)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_101),
.B(n_79),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_209),
.B1(n_105),
.B2(n_59),
.Y(n_218)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_212),
.A2(n_215),
.B1(n_220),
.B2(n_229),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_248),
.C(n_197),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_182),
.A2(n_161),
.B1(n_122),
.B2(n_103),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_161),
.B1(n_103),
.B2(n_122),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_152),
.B1(n_128),
.B2(n_139),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_234),
.A2(n_241),
.B1(n_245),
.B2(n_246),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_152),
.B1(n_156),
.B2(n_93),
.Y(n_241)
);

AOI32xp33_ASAP7_75t_L g243 ( 
.A1(n_175),
.A2(n_104),
.A3(n_160),
.B1(n_131),
.B2(n_136),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_170),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_190),
.A2(n_127),
.B1(n_139),
.B2(n_128),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_165),
.B1(n_211),
.B2(n_184),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_164),
.B(n_133),
.C(n_160),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_191),
.B(n_197),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_249),
.Y(n_288)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_250),
.A2(n_258),
.B1(n_262),
.B2(n_263),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_223),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_256),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_166),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_259),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_158),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_173),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_172),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_269),
.Y(n_295)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_179),
.B1(n_205),
.B2(n_202),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_209),
.C(n_188),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_277),
.C(n_159),
.Y(n_289)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_219),
.Y(n_303)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_212),
.A2(n_137),
.B1(n_163),
.B2(n_108),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_279),
.B1(n_248),
.B2(n_232),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_169),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_235),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_271),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_170),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_215),
.A2(n_199),
.B1(n_178),
.B2(n_187),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_273),
.B1(n_263),
.B2(n_255),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_220),
.A2(n_178),
.B1(n_203),
.B2(n_176),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_198),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_183),
.C(n_180),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_133),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_245),
.A2(n_243),
.B1(n_236),
.B2(n_234),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_253),
.B(n_214),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_280),
.B(n_303),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_292),
.B1(n_301),
.B2(n_305),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_289),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_214),
.B1(n_232),
.B2(n_237),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_256),
.B1(n_254),
.B2(n_271),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_237),
.B1(n_221),
.B2(n_239),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_230),
.C(n_223),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_304),
.C(n_136),
.Y(n_338)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_228),
.A3(n_240),
.B1(n_219),
.B2(n_233),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_300),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_240),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_221),
.B1(n_239),
.B2(n_231),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_252),
.A2(n_168),
.B1(n_181),
.B2(n_200),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_307),
.B1(n_268),
.B2(n_256),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_230),
.C(n_228),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_221),
.B1(n_231),
.B2(n_247),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_233),
.B(n_224),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_306),
.A2(n_257),
.B(n_260),
.C(n_284),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_137),
.B1(n_247),
.B2(n_108),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_224),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_276),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_310),
.B(n_278),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_259),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_312),
.B(n_316),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_290),
.B(n_264),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_325),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_249),
.B(n_271),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_314),
.A2(n_273),
.B(n_272),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_296),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_315),
.A2(n_328),
.B1(n_342),
.B2(n_344),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_254),
.B1(n_271),
.B2(n_256),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_322),
.A2(n_333),
.B1(n_308),
.B2(n_306),
.Y(n_353)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_299),
.B(n_264),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_277),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_331),
.Y(n_361)
);

INVx13_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_294),
.C(n_308),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_277),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_332),
.A2(n_343),
.B(n_344),
.C(n_342),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_249),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_334),
.A2(n_308),
.B(n_292),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_254),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_289),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_307),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_176),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_339),
.B(n_341),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_300),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_343),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_208),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_283),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_332),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_338),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_356),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_333),
.B1(n_336),
.B2(n_301),
.Y(n_347)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_294),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_354),
.B(n_363),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_302),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_317),
.A2(n_305),
.B1(n_306),
.B2(n_285),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_369),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_329),
.C(n_321),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_313),
.B(n_311),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_375),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_357),
.B(n_377),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_335),
.B(n_42),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_44),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_366),
.B(n_370),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_317),
.A2(n_306),
.B1(n_258),
.B2(n_250),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_44),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_340),
.B(n_267),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_371),
.B(n_14),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_319),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_374),
.Y(n_397)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_336),
.A2(n_306),
.B1(n_258),
.B2(n_250),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_331),
.B(n_326),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_314),
.B(n_30),
.Y(n_377)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_329),
.A2(n_267),
.B1(n_262),
.B2(n_36),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_378),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_382),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_369),
.B1(n_374),
.B2(n_378),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_385),
.A2(n_147),
.B(n_58),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_404),
.Y(n_430)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_334),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_394),
.B(n_407),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_318),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_336),
.C(n_328),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_400),
.C(n_360),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_350),
.C(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_402),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_405),
.Y(n_434)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_336),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_406),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_262),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_373),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_408),
.B(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_398),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_410),
.B(n_415),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_425),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_387),
.B(n_348),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_412),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_391),
.A2(n_355),
.B1(n_367),
.B2(n_352),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_380),
.B(n_359),
.C(n_375),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_393),
.A2(n_347),
.B1(n_353),
.B2(n_355),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_418),
.A2(n_397),
.B1(n_396),
.B2(n_381),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_419),
.A2(n_422),
.B1(n_428),
.B2(n_119),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_361),
.C(n_377),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_420),
.B(n_396),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_361),
.B1(n_362),
.B2(n_364),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_390),
.A2(n_376),
.B1(n_43),
.B2(n_36),
.Y(n_423)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

XNOR2x1_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_116),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_392),
.B(n_64),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_431),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_390),
.A2(n_43),
.B1(n_36),
.B2(n_89),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_382),
.B(n_400),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_432),
.A2(n_405),
.B(n_404),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_393),
.A2(n_395),
.B1(n_406),
.B2(n_385),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_397),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_429),
.A2(n_383),
.B(n_395),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_435),
.B(n_439),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_388),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_438),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_379),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_399),
.C(n_394),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_440),
.B(n_445),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_384),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_443),
.B(n_449),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_407),
.C(n_403),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_414),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_431),
.C(n_411),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_434),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_451),
.A2(n_427),
.B1(n_428),
.B2(n_425),
.Y(n_466)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_453),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_12),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_119),
.C(n_147),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_426),
.Y(n_471)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_422),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_461),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_435),
.A2(n_418),
.B(n_417),
.Y(n_459)
);

AOI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_459),
.A2(n_10),
.B(n_14),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_433),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_453),
.A2(n_413),
.B(n_419),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_466),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_468),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_448),
.A2(n_432),
.B(n_423),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_475),
.Y(n_485)
);

NOR2x1_ASAP7_75t_SL g474 ( 
.A(n_452),
.B(n_11),
.Y(n_474)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_474),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_22),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_22),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_454),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_469),
.A2(n_444),
.B(n_439),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_491),
.B(n_9),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_450),
.C(n_440),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_482),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_460),
.A2(n_455),
.B1(n_446),
.B2(n_441),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_481),
.B(n_490),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_470),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_441),
.C(n_446),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_488),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_455),
.C(n_456),
.Y(n_488)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_472),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_472),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_459),
.Y(n_495)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_493),
.B(n_494),
.Y(n_507)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_473),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_495),
.B(n_496),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_478),
.Y(n_496)
);

NOR3xp33_ASAP7_75t_SL g498 ( 
.A(n_487),
.B(n_462),
.C(n_467),
.Y(n_498)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

AO221x1_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_464),
.B1(n_465),
.B2(n_468),
.C(n_20),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_499),
.B(n_503),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_464),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_478),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_504),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_487),
.A2(n_27),
.B1(n_9),
.B2(n_14),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_505),
.B(n_508),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_11),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_488),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_516),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_481),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_501),
.C(n_502),
.Y(n_521)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_498),
.B(n_491),
.CI(n_483),
.CON(n_516),
.SN(n_516)
);

AOI322xp5_ASAP7_75t_L g517 ( 
.A1(n_506),
.A2(n_485),
.A3(n_9),
.B1(n_26),
.B2(n_4),
.C1(n_0),
.C2(n_2),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_517),
.A2(n_0),
.B(n_1),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_507),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_522),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_523),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_504),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_505),
.B(n_26),
.Y(n_523)
);

AOI221xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_518),
.B1(n_509),
.B2(n_520),
.C(n_516),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_0),
.Y(n_529)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_520),
.A2(n_515),
.B(n_517),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_1),
.B(n_2),
.Y(n_530)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_530),
.A3(n_526),
.B1(n_2),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_528),
.C(n_4),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_1),
.C(n_5),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_5),
.Y(n_534)
);


endmodule