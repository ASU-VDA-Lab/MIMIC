module fake_jpeg_15436_n_288 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_15),
.B1(n_29),
.B2(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_49),
.B1(n_15),
.B2(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_40),
.B(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_15),
.B1(n_27),
.B2(n_29),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_54),
.B(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_47),
.Y(n_95)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_70),
.B1(n_21),
.B2(n_28),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_27),
.B1(n_29),
.B2(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_75),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_43),
.B1(n_41),
.B2(n_19),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_88),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_48),
.B1(n_17),
.B2(n_22),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_94),
.B1(n_97),
.B2(n_105),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_88)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_20),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_33),
.B1(n_46),
.B2(n_44),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_44),
.B1(n_38),
.B2(n_28),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_61),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_108),
.Y(n_148)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_74),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_35),
.C(n_68),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_132),
.C(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_20),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_128),
.Y(n_143)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_68),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_20),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_91),
.B1(n_56),
.B2(n_66),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_127),
.B(n_23),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_80),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_24),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_83),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_68),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_121),
.Y(n_152)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_102),
.B1(n_91),
.B2(n_98),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_38),
.C(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_83),
.B1(n_94),
.B2(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_155),
.B1(n_131),
.B2(n_23),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_99),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_151),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_96),
.B(n_99),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_144),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_147),
.B(n_152),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_125),
.B(n_111),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_125),
.B(n_122),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_158),
.B(n_159),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_90),
.C(n_106),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_60),
.B(n_0),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_5),
.B(n_9),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_81),
.B1(n_60),
.B2(n_25),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_10),
.B1(n_14),
.B2(n_2),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_7),
.B1(n_14),
.B2(n_2),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_23),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_32),
.B(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_25),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_108),
.B1(n_117),
.B2(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_178),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_171),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_126),
.B1(n_123),
.B2(n_32),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_126),
.B1(n_1),
.B2(n_0),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_16),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_160),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_173),
.Y(n_209)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_16),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_186),
.Y(n_193)
);

AO21x2_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_16),
.B1(n_1),
.B2(n_3),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_159),
.B(n_162),
.Y(n_206)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_185),
.B(n_190),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_1),
.B(n_4),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_137),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_147),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_141),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_151),
.C(n_142),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_199),
.C(n_203),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_190),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_183),
.B(n_178),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_144),
.B(n_153),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_148),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_214),
.C(n_197),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_164),
.C(n_168),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_183),
.B1(n_182),
.B2(n_178),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_225),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_187),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_229),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_228),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_200),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_187),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_193),
.B1(n_207),
.B2(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_177),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_178),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_236),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_198),
.B1(n_182),
.B2(n_193),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_189),
.B1(n_165),
.B2(n_176),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_166),
.B1(n_204),
.B2(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_240),
.C(n_241),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_202),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_195),
.C(n_210),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_239),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_214),
.C(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_216),
.B1(n_222),
.B2(n_215),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_185),
.B1(n_173),
.B2(n_154),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_161),
.B1(n_231),
.B2(n_155),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_255),
.B(n_231),
.Y(n_260)
);

AOI321xp33_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_200),
.A3(n_217),
.B1(n_189),
.B2(n_185),
.C(n_208),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_253),
.A2(n_249),
.B(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_167),
.C(n_139),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_140),
.Y(n_264)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_219),
.B(n_236),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_251),
.B(n_253),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_240),
.CI(n_245),
.CON(n_259),
.SN(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_254),
.C(n_251),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_262),
.B1(n_169),
.B2(n_196),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_9),
.C(n_10),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_245),
.C(n_158),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_143),
.C(n_181),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_261),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_10),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_273),
.B(n_271),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_276),
.B1(n_265),
.B2(n_14),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_279),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_11),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_12),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_12),
.Y(n_288)
);


endmodule