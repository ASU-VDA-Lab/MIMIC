module fake_jpeg_5914_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_30),
.Y(n_49)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_19),
.Y(n_38)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_14),
.B1(n_13),
.B2(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_46),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_45),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_53),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_44),
.B1(n_51),
.B2(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_34),
.B1(n_28),
.B2(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_29),
.C(n_31),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_61),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_42),
.B1(n_52),
.B2(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_61),
.B1(n_67),
.B2(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_67),
.C(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_15),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_21),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_90),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_95),
.C(n_77),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_78),
.B1(n_77),
.B2(n_70),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_54),
.B(n_63),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_69),
.B(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_73),
.B(n_75),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_94),
.A3(n_99),
.B1(n_97),
.B2(n_93),
.C1(n_26),
.C2(n_20),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_114),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_113),
.C(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_70),
.B1(n_30),
.B2(n_56),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_115),
.B1(n_71),
.B2(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_14),
.B1(n_25),
.B2(n_19),
.Y(n_113)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_56),
.B(n_48),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_43),
.B1(n_35),
.B2(n_31),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_48),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_129),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_91),
.B1(n_95),
.B2(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_128),
.C(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_104),
.B(n_101),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_112),
.B1(n_107),
.B2(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_58),
.A3(n_20),
.B1(n_53),
.B2(n_48),
.C1(n_43),
.C2(n_35),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_71),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_102),
.B(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_136),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_134),
.C(n_13),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_101),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_114),
.B(n_110),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_139),
.B(n_142),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_21),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_141),
.A2(n_117),
.B1(n_127),
.B2(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_146),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_148),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_123),
.B1(n_124),
.B2(n_12),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_18),
.B1(n_58),
.B2(n_21),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_47),
.B1(n_18),
.B2(n_3),
.Y(n_156)
);

AOI31xp33_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_13),
.A3(n_21),
.B(n_10),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_21),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_18),
.B(n_2),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_13),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_47),
.C(n_13),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_142),
.C(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.C(n_158),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_149),
.B1(n_152),
.B2(n_151),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_1),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_1),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_18),
.B(n_2),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_3),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_164),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_4),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_154),
.C(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_5),
.C(n_7),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_160),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_5),
.B(n_8),
.Y(n_174)
);

AOI31xp67_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_4),
.A3(n_5),
.B(n_7),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_167),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.C(n_168),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);


endmodule