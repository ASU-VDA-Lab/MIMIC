module real_aes_8393_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_0), .A2(n_235), .B1(n_348), .B2(n_352), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_1), .A2(n_110), .B1(n_355), .B2(n_361), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_2), .A2(n_248), .B1(n_419), .B2(n_422), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_3), .A2(n_91), .B1(n_379), .B2(n_584), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_4), .B(n_402), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_5), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_6), .A2(n_27), .B1(n_444), .B2(n_558), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_7), .A2(n_268), .B1(n_404), .B2(n_452), .C(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_8), .A2(n_206), .B1(n_433), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_9), .A2(n_102), .B1(n_312), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_10), .A2(n_170), .B1(n_429), .B2(n_518), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_11), .A2(n_166), .B1(n_584), .B2(n_585), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g486 ( .A1(n_12), .A2(n_487), .B(n_488), .C(n_493), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_13), .A2(n_129), .B1(n_405), .B2(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_14), .Y(n_877) );
XOR2x2_ASAP7_75t_L g878 ( .A(n_14), .B(n_851), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_15), .Y(n_669) );
OA22x2_ASAP7_75t_L g785 ( .A1(n_16), .A2(n_786), .B1(n_787), .B2(n_810), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_16), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_17), .A2(n_183), .B1(n_563), .B2(n_586), .Y(n_853) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_18), .A2(n_255), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_19), .A2(n_124), .B1(n_518), .B2(n_593), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_20), .A2(n_217), .B1(n_367), .B2(n_371), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_21), .A2(n_147), .B1(n_327), .B2(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_22), .A2(n_145), .B1(n_500), .B2(n_501), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_23), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g779 ( .A1(n_24), .A2(n_131), .B1(n_163), .B2(n_459), .C1(n_514), .C2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_25), .A2(n_189), .B1(n_500), .B2(n_659), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_26), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_28), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_29), .A2(n_232), .B1(n_429), .B2(n_484), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_30), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_31), .A2(n_40), .B1(n_445), .B2(n_592), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_32), .A2(n_261), .B1(n_328), .B2(n_415), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_33), .A2(n_176), .B1(n_348), .B2(n_375), .Y(n_447) );
AO22x2_ASAP7_75t_L g294 ( .A1(n_34), .A2(n_86), .B1(n_295), .B2(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g845 ( .A(n_34), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_35), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_36), .A2(n_39), .B1(n_460), .B2(n_474), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_37), .A2(n_68), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_38), .A2(n_99), .B1(n_441), .B2(n_584), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_41), .A2(n_42), .B1(n_452), .B2(n_809), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_43), .A2(n_577), .B1(n_615), .B2(n_616), .Y(n_576) );
INVx1_ASAP7_75t_L g615 ( .A(n_43), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_44), .A2(n_62), .B1(n_544), .B2(n_545), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_45), .A2(n_262), .B1(n_411), .B2(n_514), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_46), .A2(n_132), .B1(n_196), .B2(n_393), .C1(n_544), .C2(n_545), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_47), .A2(n_125), .B1(n_355), .B2(n_797), .Y(n_796) );
AO22x2_ASAP7_75t_L g298 ( .A1(n_48), .A2(n_89), .B1(n_295), .B2(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g846 ( .A(n_48), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_49), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_50), .A2(n_234), .B1(n_369), .B2(n_377), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_51), .A2(n_70), .B1(n_415), .B2(n_455), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_52), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_53), .A2(n_157), .B1(n_212), .B2(n_457), .C1(n_458), .C2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_54), .A2(n_104), .B1(n_445), .B2(n_557), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_55), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_56), .A2(n_191), .B1(n_379), .B2(n_581), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_57), .B(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_58), .A2(n_270), .B1(n_380), .B2(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_59), .Y(n_309) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_60), .A2(n_80), .B1(n_409), .B2(n_413), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_61), .Y(n_548) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_63), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_64), .A2(n_238), .B1(n_571), .B2(n_582), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_65), .A2(n_388), .B1(n_389), .B2(n_435), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_65), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_66), .A2(n_144), .B1(n_411), .B2(n_415), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_67), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_69), .A2(n_241), .B1(n_431), .B2(n_770), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_71), .A2(n_190), .B1(n_349), .B2(n_659), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_72), .B(n_405), .Y(n_821) );
INVx1_ASAP7_75t_L g866 ( .A(n_73), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_74), .A2(n_165), .B1(n_503), .B2(n_589), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_75), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_76), .A2(n_158), .B1(n_421), .B2(n_501), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_77), .A2(n_260), .B1(n_313), .B2(n_329), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_78), .A2(n_750), .B1(n_781), .B2(n_782), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_78), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_79), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_81), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_82), .A2(n_207), .B1(n_416), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_83), .A2(n_161), .B1(n_592), .B2(n_594), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_84), .A2(n_133), .B1(n_483), .B2(n_503), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_85), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_87), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_88), .A2(n_137), .B1(n_581), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_90), .A2(n_209), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_92), .A2(n_181), .B1(n_741), .B2(n_743), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_93), .Y(n_755) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_94), .A2(n_272), .B(n_280), .C(n_847), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_95), .A2(n_254), .B1(n_482), .B2(n_484), .Y(n_481) );
AND2x2_ASAP7_75t_L g278 ( .A(n_96), .B(n_279), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_97), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_98), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_100), .A2(n_116), .B1(n_442), .B2(n_555), .Y(n_623) );
INVx1_ASAP7_75t_L g275 ( .A(n_101), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_103), .A2(n_188), .B1(n_421), .B2(n_501), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_105), .B(n_361), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_106), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_107), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_108), .A2(n_167), .B1(n_401), .B2(n_405), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_109), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_111), .A2(n_139), .B1(n_473), .B2(n_474), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_112), .A2(n_149), .B1(n_444), .B2(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_113), .A2(n_114), .B1(n_361), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_115), .A2(n_143), .B1(n_313), .B2(n_411), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_117), .A2(n_213), .B1(n_553), .B2(n_555), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_118), .A2(n_150), .B1(n_473), .B2(n_474), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_119), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_120), .A2(n_231), .B1(n_479), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_121), .A2(n_128), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_122), .A2(n_221), .B1(n_401), .B2(n_405), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_123), .A2(n_164), .B1(n_500), .B2(n_625), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_126), .Y(n_777) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_127), .A2(n_216), .B1(n_353), .B2(n_357), .Y(n_814) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_130), .A2(n_179), .B1(n_482), .B2(n_553), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_134), .B(n_327), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_135), .A2(n_219), .B1(n_478), .B2(n_585), .Y(n_651) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_136), .B(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_138), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_140), .A2(n_214), .B1(n_375), .B2(n_379), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_141), .Y(n_336) );
XNOR2x2_ASAP7_75t_L g437 ( .A(n_142), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g279 ( .A(n_146), .Y(n_279) );
XOR2xp5_ASAP7_75t_L g848 ( .A(n_148), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g712 ( .A(n_151), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_152), .B(n_402), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_153), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_154), .A2(n_264), .B1(n_557), .B2(n_558), .Y(n_556) );
AND2x6_ASAP7_75t_L g274 ( .A(n_155), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_155), .Y(n_839) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_156), .A2(n_224), .B1(n_295), .B2(n_299), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_159), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_160), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_162), .A2(n_252), .B1(n_328), .B2(n_415), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_168), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_169), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_171), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_172), .A2(n_211), .B1(n_314), .B2(n_411), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_173), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_174), .B(n_702), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_175), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_177), .A2(n_269), .B1(n_511), .B2(n_862), .Y(n_861) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_178), .A2(n_240), .B1(n_295), .B2(n_296), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_180), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_182), .A2(n_267), .B1(n_349), .B2(n_444), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_184), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_185), .A2(n_220), .B1(n_349), .B2(n_367), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_186), .B(n_401), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_187), .A2(n_253), .B1(n_855), .B2(n_856), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_192), .A2(n_215), .B1(n_433), .B2(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_193), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_194), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_195), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_197), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_198), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g477 ( .A1(n_199), .A2(n_236), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_200), .A2(n_201), .B1(n_431), .B2(n_433), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_202), .A2(n_265), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_203), .A2(n_237), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_204), .A2(n_205), .B1(n_653), .B2(n_655), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_208), .B(n_402), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_210), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_218), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_222), .Y(n_537) );
AOI22x1_ASAP7_75t_L g663 ( .A1(n_223), .A2(n_664), .B1(n_689), .B2(n_690), .Y(n_663) );
INVx1_ASAP7_75t_L g689 ( .A(n_223), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_224), .B(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_225), .Y(n_286) );
OA22x2_ASAP7_75t_L g639 ( .A1(n_226), .A2(n_640), .B1(n_641), .B2(n_661), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_226), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_227), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_228), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_229), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_230), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_233), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_239), .Y(n_818) );
INVx1_ASAP7_75t_L g842 ( .A(n_240), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_242), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_243), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_244), .B(n_398), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_245), .Y(n_394) );
OA22x2_ASAP7_75t_L g529 ( .A1(n_246), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_246), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_247), .B(n_404), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_249), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_250), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_251), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_256), .Y(n_604) );
INVx1_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_257), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_258), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_259), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_263), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_266), .Y(n_644) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_275), .Y(n_838) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_276), .A2(n_837), .B(n_876), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_716), .B1(n_717), .B2(n_833), .C(n_834), .Y(n_280) );
INVxp67_ASAP7_75t_L g833 ( .A(n_281), .Y(n_833) );
XOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_524), .Y(n_281) );
AOI22xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_461), .B1(n_462), .B2(n_523), .Y(n_282) );
INVx1_ASAP7_75t_L g523 ( .A(n_283), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_382), .B2(n_383), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
XNOR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_345), .Y(n_287) );
NOR3xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_310), .C(n_332), .Y(n_288) );
OAI22xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_305), .B1(n_306), .B2(n_309), .Y(n_289) );
INVx1_ASAP7_75t_L g536 ( .A(n_290), .Y(n_536) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g598 ( .A(n_291), .Y(n_598) );
INVx2_ASAP7_75t_L g724 ( .A(n_291), .Y(n_724) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_300), .Y(n_291) );
INVx2_ASAP7_75t_L g370 ( .A(n_292), .Y(n_370) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_298), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_293), .B(n_298), .Y(n_308) );
AND2x2_ASAP7_75t_L g351 ( .A(n_293), .B(n_317), .Y(n_351) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g318 ( .A(n_294), .B(n_304), .Y(n_318) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_298), .Y(n_322) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_297), .Y(n_299) );
INVx2_ASAP7_75t_L g317 ( .A(n_298), .Y(n_317) );
INVx1_ASAP7_75t_L g363 ( .A(n_298), .Y(n_363) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_301), .B(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g381 ( .A(n_301), .B(n_351), .Y(n_381) );
AND2x6_ASAP7_75t_L g402 ( .A(n_301), .B(n_308), .Y(n_402) );
AND2x4_ASAP7_75t_L g407 ( .A(n_301), .B(n_370), .Y(n_407) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g316 ( .A(n_302), .Y(n_316) );
INVx1_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
INVx1_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_302), .B(n_304), .Y(n_364) );
AND2x2_ASAP7_75t_L g323 ( .A(n_303), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g360 ( .A(n_304), .B(n_343), .Y(n_360) );
BUFx3_ASAP7_75t_L g538 ( .A(n_306), .Y(n_538) );
INVx2_ASAP7_75t_L g727 ( .A(n_306), .Y(n_727) );
BUFx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g601 ( .A(n_307), .Y(n_601) );
AND2x4_ASAP7_75t_L g353 ( .A(n_308), .B(n_323), .Y(n_353) );
AND2x2_ASAP7_75t_L g359 ( .A(n_308), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_308), .B(n_360), .Y(n_491) );
OAI222xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_319), .B1(n_320), .B2(n_325), .C1(n_326), .C2(n_331), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_314), .Y(n_398) );
BUFx2_ASAP7_75t_L g458 ( .A(n_314), .Y(n_458) );
BUFx4f_ASAP7_75t_SL g514 ( .A(n_314), .Y(n_514) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_314), .Y(n_606) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g330 ( .A(n_316), .Y(n_330) );
INVx1_ASAP7_75t_L g335 ( .A(n_317), .Y(n_335) );
AND2x4_ASAP7_75t_L g329 ( .A(n_318), .B(n_330), .Y(n_329) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_318), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g411 ( .A(n_318), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
BUFx3_ASAP7_75t_L g457 ( .A(n_321), .Y(n_457) );
INVx4_ASAP7_75t_L g507 ( .A(n_321), .Y(n_507) );
INVx2_ASAP7_75t_L g667 ( .A(n_321), .Y(n_667) );
AND2x6_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g340 ( .A(n_322), .Y(n_340) );
AND2x4_ASAP7_75t_L g416 ( .A(n_322), .B(n_342), .Y(n_416) );
AND2x2_ASAP7_75t_L g350 ( .A(n_323), .B(n_351), .Y(n_350) );
AND2x6_ASAP7_75t_L g369 ( .A(n_323), .B(n_370), .Y(n_369) );
OAI222xp33_ASAP7_75t_L g643 ( .A1(n_326), .A2(n_603), .B1(n_605), .B2(n_644), .C1(n_645), .C2(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx4f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx12f_ASAP7_75t_L g460 ( .A(n_329), .Y(n_460) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_329), .Y(n_470) );
INVx1_ASAP7_75t_L g804 ( .A(n_329), .Y(n_804) );
OAI22xp5_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_336), .B1(n_337), .B2(n_344), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp33_ASAP7_75t_SL g547 ( .A1(n_334), .A2(n_337), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx4_ASAP7_75t_L g613 ( .A(n_334), .Y(n_613) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_334), .Y(n_736) );
AND2x2_ASAP7_75t_L g501 ( .A(n_335), .B(n_373), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_337), .A2(n_611), .B1(n_612), .B2(n_614), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_337), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g677 ( .A(n_338), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g778 ( .A(n_339), .Y(n_778) );
OR2x6_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_365), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_354), .Y(n_346) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_349), .Y(n_428) );
BUFx3_ASAP7_75t_L g584 ( .A(n_349), .Y(n_584) );
INVx3_ASAP7_75t_L g742 ( .A(n_349), .Y(n_742) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_SL g487 ( .A(n_350), .Y(n_487) );
INVx2_ASAP7_75t_L g554 ( .A(n_350), .Y(n_554) );
BUFx2_ASAP7_75t_SL g770 ( .A(n_350), .Y(n_770) );
AND2x4_ASAP7_75t_L g372 ( .A(n_351), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_360), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_351), .B(n_360), .Y(n_567) );
INVx1_ASAP7_75t_L g688 ( .A(n_352), .Y(n_688) );
BUFx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx6_ASAP7_75t_L g434 ( .A(n_353), .Y(n_434) );
BUFx3_ASAP7_75t_L g478 ( .A(n_353), .Y(n_478) );
BUFx3_ASAP7_75t_L g518 ( .A(n_353), .Y(n_518) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_357), .Y(n_557) );
INVx4_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g425 ( .A(n_358), .Y(n_425) );
INVx3_ASAP7_75t_L g444 ( .A(n_358), .Y(n_444) );
INVx5_ASAP7_75t_L g593 ( .A(n_358), .Y(n_593) );
INVx1_ASAP7_75t_L g654 ( .A(n_358), .Y(n_654) );
INVx2_ASAP7_75t_L g855 ( .A(n_358), .Y(n_855) );
INVx8_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g445 ( .A(n_362), .Y(n_445) );
INVx6_ASAP7_75t_SL g559 ( .A(n_362), .Y(n_559) );
INVx1_ASAP7_75t_SL g797 ( .A(n_362), .Y(n_797) );
OR2x6_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g412 ( .A(n_363), .Y(n_412) );
INVx1_ASAP7_75t_L g373 ( .A(n_364), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_374), .Y(n_365) );
INVx1_ASAP7_75t_L g793 ( .A(n_367), .Y(n_793) );
INVx5_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g449 ( .A(n_368), .Y(n_449) );
INVx2_ASAP7_75t_SL g517 ( .A(n_368), .Y(n_517) );
INVx2_ASAP7_75t_L g555 ( .A(n_368), .Y(n_555) );
INVx1_ASAP7_75t_L g658 ( .A(n_368), .Y(n_658) );
INVx11_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx11_ASAP7_75t_L g432 ( .A(n_369), .Y(n_432) );
BUFx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g422 ( .A(n_372), .Y(n_422) );
BUFx3_ASAP7_75t_L g442 ( .A(n_372), .Y(n_442) );
INVx1_ASAP7_75t_L g485 ( .A(n_372), .Y(n_485) );
BUFx3_ASAP7_75t_L g503 ( .A(n_372), .Y(n_503) );
BUFx3_ASAP7_75t_L g659 ( .A(n_372), .Y(n_659) );
BUFx2_ASAP7_75t_SL g743 ( .A(n_372), .Y(n_743) );
BUFx3_ASAP7_75t_L g757 ( .A(n_372), .Y(n_757) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx4f_ASAP7_75t_SL g429 ( .A(n_377), .Y(n_429) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g480 ( .A(n_378), .Y(n_480) );
BUFx3_ASAP7_75t_L g500 ( .A(n_378), .Y(n_500) );
BUFx3_ASAP7_75t_L g586 ( .A(n_378), .Y(n_586) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
BUFx3_ASAP7_75t_L g483 ( .A(n_381), .Y(n_483) );
BUFx3_ASAP7_75t_L g571 ( .A(n_381), .Y(n_571) );
INVx2_ASAP7_75t_L g590 ( .A(n_381), .Y(n_590) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_436), .B2(n_437), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
NAND3x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_417), .C(n_426), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_399), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_395), .Y(n_391) );
OAI21xp5_ASAP7_75t_SL g467 ( .A1(n_392), .A2(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g800 ( .A(n_393), .Y(n_800) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g544 ( .A(n_398), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .C(n_408), .Y(n_399) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g453 ( .A(n_402), .Y(n_453) );
BUFx4f_ASAP7_75t_L g862 ( .A(n_402), .Y(n_862) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx5_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g511 ( .A(n_406), .Y(n_511) );
INVx2_ASAP7_75t_L g702 ( .A(n_406), .Y(n_702) );
INVx2_ASAP7_75t_L g809 ( .A(n_406), .Y(n_809) );
INVx4_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g473 ( .A(n_411), .Y(n_473) );
BUFx3_ASAP7_75t_L g864 ( .A(n_411), .Y(n_864) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .Y(n_417) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx4_ASAP7_75t_L g441 ( .A(n_420), .Y(n_441) );
INVx4_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .Y(n_426) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_432), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g581 ( .A(n_432), .Y(n_581) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g563 ( .A(n_434), .Y(n_563) );
INVx3_ASAP7_75t_L g582 ( .A(n_434), .Y(n_582) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND4xp75_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .C(n_450), .D(n_456), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .Y(n_439) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
BUFx4f_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g546 ( .A(n_460), .Y(n_546) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OAI22x1_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_495), .B1(n_521), .B2(n_522), .Y(n_463) );
INVx1_ASAP7_75t_L g521 ( .A(n_464), .Y(n_521) );
NAND3x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .C(n_486), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
BUFx2_ASAP7_75t_L g609 ( .A(n_470), .Y(n_609) );
BUFx3_ASAP7_75t_L g731 ( .A(n_470), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g754 ( .A(n_482), .Y(n_754) );
BUFx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_485), .A2(n_569), .B1(n_570), .B2(n_572), .Y(n_568) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_492), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_490), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
BUFx2_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g522 ( .A(n_495), .Y(n_522) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_520), .Y(n_496) );
NAND3x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .C(n_515), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .Y(n_498) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
BUFx2_ASAP7_75t_L g603 ( .A(n_507), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_507), .A2(n_818), .B(n_819), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .C(n_513), .Y(n_509) );
INVx1_ASAP7_75t_L g802 ( .A(n_514), .Y(n_802) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_637), .B2(n_715), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_573), .B2(n_574), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_550), .Y(n_532) );
NOR3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_540), .C(n_547), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_537), .B1(n_538), .B2(n_539), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI21xp33_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_542), .B(n_543), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g865 ( .A1(n_541), .A2(n_866), .B(n_867), .Y(n_865) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_560), .C(n_568), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g625 ( .A(n_554), .Y(n_625) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx4f_ASAP7_75t_SL g594 ( .A(n_559), .Y(n_594) );
BUFx2_ASAP7_75t_L g655 ( .A(n_559), .Y(n_655) );
BUFx2_ASAP7_75t_L g856 ( .A(n_559), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B1(n_564), .B2(n_565), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_562), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g772 ( .A(n_566), .Y(n_772) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_617), .B1(n_618), .B2(n_636), .Y(n_575) );
INVx1_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
INVx1_ASAP7_75t_SL g616 ( .A(n_577), .Y(n_616) );
AND2x2_ASAP7_75t_SL g577 ( .A(n_578), .B(n_595), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_587), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g765 ( .A(n_581), .Y(n_765) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_602), .C(n_610), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_598), .A2(n_600), .B1(n_672), .B2(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g628 ( .A(n_601), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_605), .B2(n_607), .C(n_608), .Y(n_602) );
INVx1_ASAP7_75t_L g780 ( .A(n_603), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_605), .A2(n_667), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_612), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
INVx3_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g776 ( .A(n_613), .Y(n_776) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
XOR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_635), .Y(n_620) );
NAND4xp75_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .C(n_631), .D(n_634), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
OA211x2_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_629), .C(n_630), .Y(n_626) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g715 ( .A(n_637), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_662), .B2(n_714), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g661 ( .A(n_641), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_650), .C(n_656), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g761 ( .A(n_655), .Y(n_761) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
INVx2_ASAP7_75t_L g682 ( .A(n_659), .Y(n_682) );
INVx1_ASAP7_75t_L g714 ( .A(n_662), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_691), .B1(n_692), .B2(n_713), .Y(n_662) );
INVx1_ASAP7_75t_L g713 ( .A(n_663), .Y(n_713) );
INVx2_ASAP7_75t_SL g690 ( .A(n_664), .Y(n_690) );
AND2x4_ASAP7_75t_L g664 ( .A(n_665), .B(n_678), .Y(n_664) );
NOR3xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_671), .C(n_674), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_667), .A2(n_698), .B(n_699), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_667), .A2(n_729), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_728) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_684), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
XOR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_712), .Y(n_694) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_696), .B(n_705), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .C(n_704), .Y(n_700) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_748), .B1(n_831), .B2(n_832), .Y(n_717) );
INVx2_ASAP7_75t_L g831 ( .A(n_718), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_738), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_728), .C(n_734), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_725), .B2(n_726), .Y(n_721) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_745), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_744), .Y(n_739) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g832 ( .A(n_748), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_783), .B1(n_829), .B2(n_830), .Y(n_748) );
INVx1_ASAP7_75t_L g830 ( .A(n_749), .Y(n_830) );
INVx1_ASAP7_75t_L g782 ( .A(n_750), .Y(n_782) );
AND4x1_ASAP7_75t_L g750 ( .A(n_751), .B(n_762), .C(n_773), .D(n_779), .Y(n_750) );
NOR2xp33_ASAP7_75t_SL g751 ( .A(n_752), .B(n_758), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_752) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B1(n_771), .B2(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_774) );
INVx2_ASAP7_75t_L g829 ( .A(n_783), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_811), .B2(n_828), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g810 ( .A(n_787), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_798), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_794), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_806), .Y(n_798) );
OAI222xp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B1(n_802), .B2(n_803), .C1(n_804), .C2(n_805), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx3_ASAP7_75t_L g828 ( .A(n_811), .Y(n_828) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_827), .Y(n_811) );
NAND3x1_ASAP7_75t_SL g812 ( .A(n_813), .B(n_816), .C(n_824), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_820), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .C(n_823), .Y(n_820) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
INVx1_ASAP7_75t_SL g834 ( .A(n_835), .Y(n_834) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_836), .B(n_840), .Y(n_835) );
OR2x2_ASAP7_75t_SL g879 ( .A(n_836), .B(n_841), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_839), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_837), .Y(n_869) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_838), .B(n_873), .Y(n_876) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_839), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
OAI322xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_868), .A3(n_870), .B1(n_874), .B2(n_877), .C1(n_878), .C2(n_879), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR4xp75_ASAP7_75t_L g851 ( .A(n_852), .B(n_857), .C(n_860), .D(n_865), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g852 ( .A(n_853), .B(n_854), .Y(n_852) );
NAND2xp5_ASAP7_75t_SL g857 ( .A(n_858), .B(n_859), .Y(n_857) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_861), .B(n_863), .Y(n_860) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx16_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
endmodule