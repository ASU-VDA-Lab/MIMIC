module fake_jpeg_25477_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_53),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_29),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_19),
.B(n_25),
.C(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_31),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_43),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_84),
.Y(n_95)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g96 ( 
.A(n_68),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_42),
.B1(n_37),
.B2(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_73),
.B(n_88),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_32),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_75),
.C(n_2),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_32),
.B(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_47),
.B1(n_64),
.B2(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_33),
.B1(n_27),
.B2(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_51),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_30),
.B1(n_21),
.B2(n_17),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_21),
.B1(n_39),
.B2(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_64),
.B1(n_55),
.B2(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_59),
.B1(n_51),
.B2(n_52),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_0),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_106),
.B(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_1),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_21),
.B1(n_63),
.B2(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_2),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_81),
.B1(n_68),
.B2(n_78),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_95),
.B1(n_90),
.B2(n_108),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_74),
.B(n_84),
.C(n_87),
.D(n_81),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_105),
.B(n_91),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_125),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_74),
.B1(n_87),
.B2(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_100),
.B1(n_94),
.B2(n_109),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_92),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_69),
.B1(n_72),
.B2(n_82),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_132),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_72),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_148),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_151),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_146),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_99),
.B(n_93),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_144),
.B(n_120),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_147),
.B1(n_112),
.B2(n_113),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_106),
.B1(n_103),
.B2(n_69),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_152),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_121),
.C(n_122),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_123),
.C(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_4),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_159),
.B1(n_168),
.B2(n_166),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_119),
.B(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_119),
.C(n_114),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_125),
.B1(n_124),
.B2(n_7),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_167),
.B1(n_152),
.B2(n_6),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_39),
.C(n_66),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_136),
.C(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_143),
.B1(n_142),
.B2(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_4),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_170),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_184),
.C(n_7),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_135),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_133),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_181),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_140),
.C(n_136),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_165),
.C(n_163),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_186),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_140),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_149),
.B1(n_153),
.B2(n_145),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_163),
.B(n_154),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_6),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_7),
.Y(n_197)
);

NAND4xp25_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_169),
.C(n_174),
.D(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_194),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_162),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_193),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_184),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_181),
.B(n_178),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_200),
.A2(n_196),
.B(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_205),
.Y(n_211)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_173),
.B1(n_185),
.B2(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_8),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_209),
.B(n_208),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_203),
.A2(n_190),
.B1(n_196),
.B2(n_11),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_8),
.B(n_10),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_11),
.A3(n_12),
.B(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_212),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_198),
.C(n_14),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_14),
.B1(n_15),
.B2(n_216),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_15),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_15),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_222),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_218),
.Y(n_225)
);


endmodule