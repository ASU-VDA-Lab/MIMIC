module fake_jpeg_16264_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_0),
.A2(n_5),
.B1(n_1),
.B2(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_29),
.B1(n_27),
.B2(n_17),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_15),
.B1(n_12),
.B2(n_19),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_23),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_34),
.B1(n_33),
.B2(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx10_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_38),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_32),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_34),
.C(n_16),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.C(n_21),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_36),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_41),
.A3(n_19),
.B1(n_11),
.B2(n_21),
.C1(n_28),
.C2(n_9),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_21),
.C2(n_39),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_9),
.B(n_11),
.Y(n_50)
);


endmodule