module fake_jpeg_22775_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_45),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_32),
.Y(n_66)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_63),
.B1(n_74),
.B2(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_64),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_71),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_79),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_17),
.B1(n_37),
.B2(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_28),
.B1(n_33),
.B2(n_35),
.Y(n_81)
);

OAI22x1_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_82),
.B1(n_30),
.B2(n_38),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_1),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_33),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_108),
.C(n_30),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_33),
.B1(n_35),
.B2(n_32),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_91),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_31),
.B1(n_42),
.B2(n_36),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_93),
.A2(n_100),
.B(n_102),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_83),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_103),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_22),
.B(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_42),
.B1(n_24),
.B2(n_20),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_49),
.B1(n_34),
.B2(n_30),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_104),
.A2(n_117),
.B1(n_119),
.B2(n_34),
.Y(n_153)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_107),
.Y(n_146)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_55),
.B(n_49),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_115),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_107),
.B1(n_105),
.B2(n_119),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_76),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_61),
.A2(n_30),
.B1(n_38),
.B2(n_19),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_120),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_92),
.B1(n_112),
.B2(n_87),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_89),
.B1(n_114),
.B2(n_103),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_43),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_134),
.C(n_89),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_127),
.A2(n_129),
.B1(n_154),
.B2(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_130),
.Y(n_166)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_132),
.B(n_136),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_50),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_142),
.B(n_116),
.Y(n_170)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_38),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_60),
.B1(n_54),
.B2(n_38),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_149),
.B1(n_121),
.B2(n_5),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_98),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_34),
.B1(n_19),
.B2(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_10),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_152),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_91),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_91),
.B1(n_34),
.B2(n_19),
.Y(n_172)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_164),
.B1(n_179),
.B2(n_183),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_120),
.B1(n_88),
.B2(n_86),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_167),
.B(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_116),
.B(n_88),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_175),
.B(n_7),
.Y(n_216)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_174),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_19),
.Y(n_175)
);

AOI22x1_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_10),
.B1(n_16),
.B2(n_3),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_4),
.Y(n_195)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_1),
.B(n_2),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_185),
.B1(n_190),
.B2(n_125),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_125),
.B(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_134),
.B1(n_133),
.B2(n_137),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

AO21x2_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_2),
.B(n_4),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_189),
.Y(n_194)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_216),
.B1(n_215),
.B2(n_185),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_208),
.B1(n_213),
.B2(n_164),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_130),
.C(n_132),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_207),
.C(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_128),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_157),
.C(n_151),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_169),
.B1(n_173),
.B2(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_145),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_210),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_173),
.A2(n_126),
.B1(n_5),
.B2(n_7),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_126),
.C(n_5),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_4),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_176),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_7),
.B(n_8),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_12),
.C(n_13),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_180),
.C(n_158),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_12),
.B(n_13),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_182),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_232),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_233),
.B1(n_219),
.B2(n_216),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_162),
.B1(n_178),
.B2(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_178),
.B1(n_185),
.B2(n_190),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_197),
.B1(n_201),
.B2(n_213),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_166),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_239),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_241),
.B(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_189),
.C(n_188),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_192),
.C(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_196),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_227),
.B1(n_229),
.B2(n_241),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_255),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_204),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_262),
.B(n_229),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_214),
.B1(n_194),
.B2(n_192),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_221),
.B(n_218),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_240),
.C(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_238),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_187),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_232),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_260),
.B1(n_248),
.B2(n_262),
.Y(n_289)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_276),
.C(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_212),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_259),
.B(n_224),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_235),
.C(n_228),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_249),
.Y(n_288)
);

AO22x1_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_233),
.B1(n_230),
.B2(n_223),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_184),
.B(n_254),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_263),
.C(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_209),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_222),
.B1(n_209),
.B2(n_167),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_284),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_224),
.C(n_226),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_250),
.C(n_168),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_295),
.C(n_297),
.Y(n_302)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_293),
.B(n_199),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_258),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_269),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_200),
.B(n_160),
.C(n_193),
.D(n_199),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_278),
.B1(n_276),
.B2(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_283),
.B1(n_272),
.B2(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_269),
.C(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_289),
.B1(n_298),
.B2(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_292),
.B1(n_291),
.B2(n_287),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_294),
.C(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_306),
.B(n_295),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_193),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_318),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_312),
.A2(n_309),
.B(n_296),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_322),
.B(n_313),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_288),
.B(n_279),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_311),
.C(n_314),
.Y(n_326)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.A3(n_325),
.B1(n_314),
.B2(n_320),
.C(n_212),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_315),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_14),
.B(n_15),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_14),
.B(n_15),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_14),
.CI(n_15),
.CON(n_331),
.SN(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_16),
.B(n_329),
.Y(n_332)
);


endmodule