module fake_ariane_745_n_1806 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1806);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1806;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_206;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_77),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_28),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_97),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_82),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_38),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_83),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_43),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_7),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_16),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_4),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_112),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_115),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_70),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_78),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_49),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_55),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_28),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_52),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_55),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_19),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_45),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_25),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_106),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_20),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_41),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_136),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_4),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_68),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_56),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_42),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_21),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_63),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_46),
.Y(n_223)
);

BUFx2_ASAP7_75t_SL g224 ( 
.A(n_131),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_8),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_105),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_100),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_153),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_36),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_31),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_20),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_74),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_42),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_37),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_60),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_51),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_61),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_108),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_113),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_148),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_12),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_36),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_124),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_127),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_130),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_41),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_54),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_35),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_35),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_48),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_99),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_155),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_81),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_123),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_48),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_87),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_90),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_14),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_23),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_62),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_23),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_26),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_140),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_135),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_89),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_94),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_72),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_47),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_54),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_15),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_67),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_128),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_134),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_73),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_49),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_34),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_12),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_102),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_103),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_114),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_75),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_46),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_85),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_39),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_86),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_88),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_66),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_10),
.Y(n_310)
);

CKINVDCx11_ASAP7_75t_R g311 ( 
.A(n_14),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_160),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_310),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_203),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_179),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_215),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_193),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_193),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_196),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_196),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_252),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_255),
.B(n_2),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_269),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_196),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_163),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_196),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_231),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_196),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_248),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_249),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_292),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_166),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_268),
.B(n_2),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_175),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_178),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_196),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_192),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_196),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_219),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_163),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_288),
.B(n_297),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_191),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_190),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_167),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_190),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_197),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_213),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_190),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_239),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_241),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_198),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_190),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_295),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_277),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_190),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_235),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_235),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_175),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_219),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_244),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_187),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_220),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_175),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_238),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_272),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_221),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_297),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_272),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_238),
.B(n_6),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_275),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_275),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_225),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_273),
.Y(n_377)
);

BUFx6f_ASAP7_75t_SL g378 ( 
.A(n_273),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_273),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_281),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_187),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_281),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_281),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_204),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_159),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_204),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_234),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_335),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_338),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_165),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_319),
.B(n_171),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_344),
.B(n_171),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

BUFx8_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_314),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_170),
.Y(n_409)
);

BUFx8_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_184),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_346),
.A2(n_176),
.B(n_172),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_173),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_341),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_368),
.B(n_180),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_325),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_207),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_355),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_381),
.B(n_182),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_330),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_386),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_320),
.B(n_184),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_364),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_369),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_372),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_340),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_368),
.B(n_181),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_402),
.B(n_349),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_406),
.B(n_337),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_454),
.B(n_354),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

BUFx4f_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_388),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_399),
.B(n_382),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_406),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_454),
.B(n_366),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_454),
.B(n_370),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_454),
.B(n_376),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_337),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_422),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_406),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_388),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_379),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_379),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_436),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_400),
.A2(n_336),
.B1(n_324),
.B2(n_314),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_342),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_400),
.A2(n_314),
.B1(n_315),
.B2(n_328),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_422),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_440),
.B(n_387),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_447),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_393),
.B(n_207),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

BUFx4f_ASAP7_75t_L g498 ( 
.A(n_414),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_395),
.B(n_385),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_393),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_326),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_391),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_391),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_438),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_443),
.B(n_371),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_414),
.B(n_212),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_395),
.B(n_347),
.C(n_343),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_392),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_406),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_393),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_417),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_395),
.B(n_373),
.C(n_174),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_406),
.A2(n_279),
.B1(n_243),
.B2(n_276),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_405),
.B(n_188),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_405),
.B(n_157),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_396),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_441),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_374),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_374),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_406),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_436),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_SL g535 ( 
.A(n_394),
.B(n_361),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_405),
.B(n_157),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_406),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_423),
.B(n_353),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_393),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_409),
.A2(n_356),
.B1(n_212),
.B2(n_195),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_407),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_393),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_393),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_446),
.B(n_375),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_442),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_423),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_407),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_389),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_393),
.B(n_169),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_389),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_421),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_394),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_408),
.B(n_158),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_394),
.B(n_334),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_394),
.B(n_158),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_408),
.B(n_367),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_404),
.B(n_169),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_396),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_456),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_402),
.B(n_169),
.Y(n_567)
);

NOR2x1p5_ASAP7_75t_L g568 ( 
.A(n_409),
.B(n_167),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_389),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_389),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_408),
.B(n_161),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_425),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_391),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_446),
.B(n_375),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_400),
.A2(n_304),
.B1(n_310),
.B2(n_298),
.Y(n_575)
);

INVx8_ASAP7_75t_L g576 ( 
.A(n_400),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_400),
.A2(n_223),
.B1(n_303),
.B2(n_287),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_428),
.B(n_224),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_400),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_404),
.B(n_169),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_445),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_411),
.B(n_377),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_428),
.A2(n_174),
.B1(n_306),
.B2(n_304),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_389),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_428),
.B(n_161),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_404),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_428),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_390),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_404),
.B(n_169),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_411),
.B(n_289),
.C(n_186),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_390),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_392),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_445),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_409),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_448),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_409),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_412),
.B(n_162),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_390),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_404),
.B(n_410),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_448),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_411),
.B(n_162),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_421),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_415),
.B(n_186),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_415),
.A2(n_306),
.B1(n_298),
.B2(n_296),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_472),
.B(n_415),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_486),
.B(n_404),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_461),
.B(n_396),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_486),
.B(n_410),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_497),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_486),
.B(n_492),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_461),
.B(n_396),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_482),
.B(n_410),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_415),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_461),
.B(n_498),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_549),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_498),
.B(n_564),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_410),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_499),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_596),
.B(n_419),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_410),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_539),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_508),
.B(n_410),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_499),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_508),
.B(n_410),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_527),
.B(n_412),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_578),
.B(n_419),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_495),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_464),
.B(n_419),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_541),
.A2(n_412),
.B1(n_414),
.B2(n_430),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_502),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_498),
.B(n_396),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_478),
.B(n_589),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_589),
.B(n_201),
.C(n_200),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_539),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_549),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_501),
.A2(n_598),
.B(n_517),
.C(n_523),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_484),
.B(n_425),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_531),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_560),
.B(n_419),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_578),
.B(n_455),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_507),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_531),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_564),
.B(n_396),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_527),
.B(n_412),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_528),
.B(n_458),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_503),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_485),
.A2(n_289),
.B1(n_290),
.B2(n_296),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_543),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_541),
.A2(n_412),
.B1(n_414),
.B2(n_430),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_518),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_576),
.A2(n_412),
.B1(n_455),
.B2(n_383),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_R g659 ( 
.A(n_484),
.B(n_317),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_564),
.B(n_401),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_SL g661 ( 
.A(n_556),
.B(n_425),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_537),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_542),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_546),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_528),
.B(n_412),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_576),
.A2(n_455),
.B1(n_380),
.B2(n_432),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_577),
.A2(n_258),
.B1(n_211),
.B2(n_217),
.C(n_218),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_483),
.B(n_401),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_601),
.B(n_402),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_548),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_519),
.B(n_401),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_543),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_576),
.B(n_401),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_578),
.B(n_455),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_547),
.B(n_401),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_568),
.A2(n_432),
.B1(n_293),
.B2(n_299),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_541),
.A2(n_432),
.B1(n_333),
.B2(n_318),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_541),
.A2(n_414),
.B1(n_430),
.B2(n_390),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_533),
.A2(n_403),
.B(n_401),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_550),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_503),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_579),
.A2(n_414),
.B1(n_390),
.B2(n_397),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_547),
.B(n_401),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_559),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_587),
.B(n_403),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_L g686 ( 
.A1(n_522),
.A2(n_290),
.B(n_250),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_574),
.B(n_518),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_574),
.B(n_403),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_518),
.B(n_403),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_599),
.B(n_525),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_578),
.B(n_425),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_558),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_525),
.B(n_403),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_513),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_525),
.B(n_403),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_530),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_559),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_561),
.B(n_259),
.C(n_240),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_583),
.A2(n_579),
.B1(n_488),
.B2(n_459),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_565),
.B(n_403),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_565),
.B(n_413),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_467),
.B(n_230),
.C(n_208),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_565),
.B(n_413),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_536),
.B(n_413),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_557),
.B(n_413),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_579),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_552),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_505),
.B(n_413),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_606),
.A2(n_397),
.B1(n_448),
.B2(n_451),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_505),
.B(n_413),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_530),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_530),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_571),
.B(n_413),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_463),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_603),
.B(n_416),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_562),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_554),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_556),
.B(n_332),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_566),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_513),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_544),
.B(n_446),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_554),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_481),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_544),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_510),
.B(n_416),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_582),
.B(n_416),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_594),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_569),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_595),
.B(n_416),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_605),
.B(n_345),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_SL g733 ( 
.A(n_540),
.B(n_446),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_597),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_602),
.B(n_416),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_468),
.B(n_416),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_569),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_511),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_505),
.B(n_416),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_505),
.B(n_418),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_479),
.A2(n_397),
.B1(n_451),
.B2(n_421),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_505),
.B(n_418),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_489),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_466),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_490),
.A2(n_451),
.B1(n_421),
.B2(n_449),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_493),
.B(n_418),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_555),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_594),
.Y(n_749)
);

CKINVDCx11_ASAP7_75t_R g750 ( 
.A(n_511),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_535),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_555),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_604),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_570),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_604),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_496),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_496),
.B(n_418),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_570),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_584),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_605),
.A2(n_421),
.B1(n_449),
.B2(n_444),
.Y(n_760)
);

BUFx6f_ASAP7_75t_SL g761 ( 
.A(n_553),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_500),
.B(n_418),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_586),
.Y(n_763)
);

O2A1O1Ixp5_ASAP7_75t_L g764 ( 
.A1(n_534),
.A2(n_418),
.B(n_446),
.C(n_424),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_506),
.B(n_418),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_535),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_500),
.B(n_446),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_601),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_532),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_532),
.B(n_446),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_551),
.B(n_439),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_469),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_506),
.B(n_402),
.Y(n_774)
);

INVxp33_ASAP7_75t_L g775 ( 
.A(n_585),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_470),
.Y(n_776)
);

AND2x2_ASAP7_75t_SL g777 ( 
.A(n_567),
.B(n_202),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_515),
.B(n_402),
.Y(n_778)
);

INVxp33_ASAP7_75t_L g779 ( 
.A(n_516),
.Y(n_779)
);

OAI321xp33_ASAP7_75t_L g780 ( 
.A1(n_653),
.A2(n_256),
.A3(n_233),
.B1(n_265),
.B2(n_245),
.C(n_263),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_668),
.A2(n_520),
.B(n_473),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_632),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_659),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_608),
.A2(n_551),
.B(n_439),
.C(n_453),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_608),
.B(n_590),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_775),
.A2(n_439),
.B(n_450),
.C(n_453),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_775),
.B(n_575),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_624),
.B(n_588),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_651),
.A2(n_520),
.B(n_473),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_646),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_764),
.A2(n_509),
.B(n_590),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_R g792 ( 
.A(n_750),
.B(n_350),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_625),
.B(n_352),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_624),
.B(n_613),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_652),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_617),
.B(n_506),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_769),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_633),
.B(n_593),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_610),
.A2(n_636),
.B(n_614),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_610),
.A2(n_520),
.B(n_473),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_614),
.A2(n_572),
.B(n_521),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_636),
.A2(n_572),
.B(n_521),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_639),
.B(n_312),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_779),
.B(n_592),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_696),
.A2(n_509),
.B(n_593),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_633),
.B(n_600),
.Y(n_806)
);

CKINVDCx10_ASAP7_75t_R g807 ( 
.A(n_750),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_648),
.A2(n_660),
.B(n_619),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_616),
.B(n_622),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_L g810 ( 
.A1(n_779),
.A2(n_622),
.B(n_616),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_648),
.A2(n_572),
.B(n_521),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_769),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_727),
.B(n_630),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_660),
.A2(n_457),
.B(n_466),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_631),
.A2(n_457),
.B1(n_529),
.B2(n_538),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_727),
.B(n_600),
.Y(n_816)
);

AOI21x1_ASAP7_75t_L g817 ( 
.A1(n_774),
.A2(n_465),
.B(n_462),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_617),
.A2(n_619),
.B(n_705),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_644),
.A2(n_264),
.B(n_261),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_650),
.B(n_494),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_684),
.B(n_509),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_644),
.A2(n_439),
.B(n_453),
.C(n_450),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_706),
.A2(n_512),
.B(n_476),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_708),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_687),
.A2(n_540),
.B1(n_545),
.B2(n_476),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_714),
.A2(n_529),
.B(n_512),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_665),
.B(n_494),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_700),
.B(n_506),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_710),
.B(n_494),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_649),
.B(n_494),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_717),
.A2(n_538),
.B(n_487),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_673),
.B(n_506),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_637),
.B(n_236),
.Y(n_833)
);

NOR2x2_ASAP7_75t_L g834 ( 
.A(n_645),
.B(n_674),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_698),
.A2(n_260),
.B(n_460),
.C(n_487),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_689),
.A2(n_487),
.B(n_460),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_645),
.B(n_545),
.Y(n_837)
);

OAI321xp33_ASAP7_75t_L g838 ( 
.A1(n_667),
.A2(n_450),
.A3(n_453),
.B1(n_439),
.B2(n_437),
.C(n_435),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_693),
.A2(n_460),
.B(n_573),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_640),
.B(n_236),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_701),
.A2(n_573),
.B(n_465),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_708),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_675),
.A2(n_424),
.B(n_433),
.C(n_453),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_723),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_657),
.B(n_494),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_697),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_641),
.A2(n_450),
.B(n_421),
.C(n_431),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_662),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_690),
.A2(n_474),
.B(n_475),
.C(n_477),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_663),
.B(n_494),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_704),
.A2(n_573),
.B(n_471),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_716),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_664),
.B(n_573),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_715),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_670),
.B(n_573),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_671),
.A2(n_471),
.B(n_462),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_692),
.B(n_718),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_721),
.B(n_450),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_734),
.B(n_421),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_696),
.A2(n_477),
.B(n_475),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_631),
.B(n_620),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_748),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_666),
.B(n_474),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_631),
.B(n_553),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_652),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_623),
.B(n_553),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_702),
.A2(n_688),
.B(n_683),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_618),
.B(n_236),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_723),
.B(n_514),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_626),
.B(n_553),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_629),
.B(n_553),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_757),
.A2(n_514),
.B(n_580),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_716),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_723),
.B(n_656),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_656),
.B(n_685),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_729),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_743),
.A2(n_424),
.B(n_433),
.C(n_437),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_762),
.A2(n_514),
.B(n_580),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_774),
.A2(n_431),
.B(n_435),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_690),
.B(n_553),
.Y(n_880)
);

BUFx4f_ASAP7_75t_SL g881 ( 
.A(n_697),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_638),
.A2(n_433),
.B(n_424),
.C(n_435),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_752),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_702),
.A2(n_514),
.B(n_580),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_685),
.A2(n_588),
.B1(n_280),
.B2(n_580),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_652),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_736),
.A2(n_580),
.B(n_514),
.Y(n_887)
);

NOR2xp67_ASAP7_75t_SL g888 ( 
.A(n_712),
.B(n_480),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_691),
.B(n_480),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_652),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_719),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_658),
.B(n_563),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_756),
.B(n_563),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_770),
.B(n_634),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_655),
.B(n_563),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_747),
.A2(n_491),
.B(n_480),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_728),
.A2(n_491),
.B(n_480),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_719),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_724),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_645),
.A2(n_283),
.B1(n_302),
.B2(n_305),
.Y(n_900)
);

AO22x1_ASAP7_75t_L g901 ( 
.A1(n_732),
.A2(n_591),
.B1(n_581),
.B2(n_563),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_681),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_753),
.A2(n_433),
.B(n_424),
.C(n_437),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_725),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_766),
.B(n_402),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_724),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_681),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_731),
.A2(n_491),
.B(n_480),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_735),
.A2(n_491),
.B(n_402),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_755),
.B(n_563),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_691),
.B(n_491),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_713),
.B(n_563),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_709),
.A2(n_402),
.B(n_567),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_659),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_679),
.A2(n_431),
.B(n_433),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_738),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_686),
.B(n_581),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_720),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_749),
.B(n_444),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_707),
.B(n_581),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_691),
.B(n_402),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_709),
.A2(n_402),
.B(n_417),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_615),
.B(n_676),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_778),
.A2(n_433),
.B(n_424),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_767),
.A2(n_424),
.B(n_433),
.C(n_429),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_711),
.A2(n_417),
.B(n_391),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_674),
.A2(n_417),
.B1(n_251),
.B2(n_246),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_778),
.A2(n_227),
.B(n_291),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_674),
.A2(n_168),
.B1(n_164),
.B2(n_177),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_711),
.A2(n_417),
.B(n_391),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_730),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_609),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_776),
.B(n_444),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_677),
.B(n_444),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_607),
.B(n_417),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_607),
.B(n_417),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_739),
.A2(n_417),
.B(n_391),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_699),
.A2(n_449),
.B(n_444),
.C(n_420),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_739),
.A2(n_429),
.B(n_420),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_773),
.B(n_417),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_740),
.A2(n_417),
.B(n_391),
.Y(n_941)
);

CKINVDCx8_ASAP7_75t_R g942 ( 
.A(n_681),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_733),
.A2(n_300),
.B(n_254),
.C(n_247),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_740),
.A2(n_391),
.B(n_164),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_742),
.A2(n_420),
.B(n_427),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_751),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_703),
.B(n_601),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_612),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_761),
.B(n_601),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_612),
.B(n_581),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_742),
.A2(n_391),
.B(n_168),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_730),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_765),
.A2(n_391),
.B(n_307),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_681),
.B(n_434),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_765),
.B(n_444),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_621),
.B(n_581),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_621),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_771),
.A2(n_185),
.B(n_183),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_SL g959 ( 
.A1(n_772),
.A2(n_232),
.B(n_237),
.C(n_262),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_627),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_611),
.B(n_444),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_627),
.B(n_581),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_737),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_628),
.B(n_591),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_628),
.A2(n_177),
.B(n_185),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_635),
.B(n_591),
.Y(n_966)
);

AOI33xp33_ASAP7_75t_L g967 ( 
.A1(n_760),
.A2(n_420),
.A3(n_427),
.B1(n_429),
.B2(n_294),
.B3(n_284),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_635),
.B(n_643),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_695),
.B(n_434),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_643),
.A2(n_183),
.B(n_283),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_SL g971 ( 
.A(n_792),
.B(n_305),
.C(n_285),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_SL g972 ( 
.A1(n_888),
.A2(n_741),
.B(n_746),
.C(n_680),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_809),
.B(n_744),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_781),
.A2(n_669),
.B(n_733),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_782),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_804),
.A2(n_777),
.B(n_661),
.C(n_682),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_942),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_789),
.A2(n_642),
.B(n_744),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_795),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_804),
.A2(n_777),
.B(n_654),
.C(n_647),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_824),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_793),
.B(n_678),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_805),
.A2(n_768),
.B(n_694),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_813),
.B(n_647),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_946),
.B(n_654),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_810),
.B(n_672),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_857),
.A2(n_672),
.B1(n_680),
.B2(n_694),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_790),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_842),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_787),
.A2(n_677),
.B1(n_763),
.B2(n_754),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_798),
.A2(n_758),
.B1(n_763),
.B2(n_754),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_914),
.B(n_695),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_833),
.B(n_677),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_923),
.A2(n_737),
.B(n_758),
.C(n_429),
.Y(n_994)
);

INVx3_ASAP7_75t_SL g995 ( 
.A(n_916),
.Y(n_995)
);

OAI22x1_ASAP7_75t_L g996 ( 
.A1(n_787),
.A2(n_285),
.B1(n_293),
.B2(n_301),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_876),
.B(n_307),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_848),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_796),
.A2(n_875),
.B(n_832),
.C(n_794),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_L g1000 ( 
.A1(n_796),
.A2(n_768),
.B(n_420),
.C(n_427),
.Y(n_1000)
);

BUFx8_ASAP7_75t_L g1001 ( 
.A(n_803),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_821),
.B(n_695),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_852),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_792),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_873),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_821),
.B(n_695),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_876),
.B(n_308),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_806),
.A2(n_785),
.B1(n_861),
.B2(n_862),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_883),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_904),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_881),
.B(n_722),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_828),
.A2(n_427),
.B(n_429),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_844),
.B(n_863),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_788),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_948),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_819),
.A2(n_427),
.B(n_8),
.C(n_9),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_875),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_818),
.A2(n_591),
.B(n_601),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_918),
.B(n_308),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_891),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_844),
.B(n_722),
.Y(n_1022)
);

INVx3_ASAP7_75t_SL g1023 ( 
.A(n_783),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_863),
.A2(n_761),
.B1(n_444),
.B2(n_449),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_881),
.B(n_309),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_900),
.A2(n_309),
.B(n_189),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_933),
.B(n_722),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_832),
.A2(n_591),
.B(n_601),
.C(n_726),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_932),
.B(n_722),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_780),
.A2(n_11),
.B(n_16),
.C(n_17),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_834),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_795),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_795),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_788),
.B(n_759),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_957),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_919),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_856),
.A2(n_759),
.B(n_745),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_SL g1038 ( 
.A(n_807),
.B(n_958),
.C(n_867),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_960),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_894),
.A2(n_449),
.B1(n_444),
.B2(n_434),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_808),
.A2(n_759),
.B(n_745),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_840),
.A2(n_759),
.B1(n_745),
.B2(n_726),
.Y(n_1042)
);

AOI22x1_ASAP7_75t_L g1043 ( 
.A1(n_799),
.A2(n_745),
.B1(n_726),
.B2(n_434),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_858),
.Y(n_1044)
);

INVx6_ASAP7_75t_L g1045 ( 
.A(n_846),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_795),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_868),
.B(n_444),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_846),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_841),
.A2(n_726),
.B(n_591),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_865),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_932),
.B(n_449),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_786),
.A2(n_449),
.B1(n_434),
.B2(n_426),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_874),
.B(n_449),
.Y(n_1053)
);

NAND3xp33_ASAP7_75t_L g1054 ( 
.A(n_784),
.B(n_786),
.C(n_905),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_929),
.B(n_194),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_865),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_898),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_899),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_837),
.B(n_449),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_794),
.B(n_434),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_851),
.A2(n_253),
.B(n_205),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_837),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_906),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_874),
.B(n_449),
.Y(n_1064)
);

OR2x6_ASAP7_75t_SL g1065 ( 
.A(n_927),
.B(n_199),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_865),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_837),
.B(n_434),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_921),
.A2(n_257),
.B1(n_210),
.B2(n_214),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_940),
.B(n_434),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_931),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_784),
.A2(n_434),
.B1(n_426),
.B2(n_266),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_865),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_797),
.B(n_812),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_860),
.A2(n_801),
.B(n_800),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_952),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_905),
.A2(n_434),
.B(n_426),
.C(n_267),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_921),
.B(n_869),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_963),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_802),
.A2(n_242),
.B(n_222),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_886),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_853),
.A2(n_434),
.B1(n_426),
.B2(n_270),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_968),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_943),
.A2(n_11),
.B(n_17),
.C(n_18),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_811),
.A2(n_229),
.B(n_226),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_886),
.B(n_206),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_940),
.A2(n_426),
.B(n_274),
.C(n_278),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_886),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_816),
.B(n_19),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_886),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_855),
.A2(n_822),
.B1(n_815),
.B2(n_829),
.Y(n_1090)
);

OR2x6_ASAP7_75t_SL g1091 ( 
.A(n_864),
.B(n_228),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_902),
.Y(n_1092)
);

BUFx8_ASAP7_75t_L g1093 ( 
.A(n_934),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_961),
.A2(n_426),
.B(n_271),
.C(n_282),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_839),
.A2(n_286),
.B(n_282),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_961),
.A2(n_426),
.B(n_286),
.C(n_282),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_859),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_838),
.B(n_426),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_836),
.A2(n_286),
.B(n_282),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_822),
.A2(n_426),
.B1(n_286),
.B2(n_282),
.Y(n_1100)
);

O2A1O1Ixp5_ASAP7_75t_SL g1101 ( 
.A1(n_828),
.A2(n_426),
.B(n_286),
.C(n_216),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_831),
.A2(n_216),
.B(n_209),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_897),
.A2(n_216),
.B(n_209),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_902),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_967),
.B(n_22),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_959),
.A2(n_22),
.B(n_24),
.C(n_25),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_965),
.B(n_24),
.C(n_26),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_902),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_959),
.A2(n_27),
.B(n_30),
.C(n_31),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_869),
.B(n_27),
.Y(n_1110)
);

O2A1O1Ixp5_ASAP7_75t_L g1111 ( 
.A1(n_814),
.A2(n_32),
.B(n_33),
.C(n_37),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_892),
.A2(n_216),
.B1(n_209),
.B2(n_39),
.Y(n_1112)
);

OA22x2_ASAP7_75t_L g1113 ( 
.A1(n_889),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_908),
.A2(n_896),
.B(n_849),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_835),
.A2(n_40),
.B(n_43),
.C(n_44),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_939),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_823),
.A2(n_216),
.B(n_209),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_826),
.A2(n_209),
.B(n_101),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_902),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_791),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_890),
.B(n_907),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_890),
.B(n_50),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_976),
.A2(n_820),
.B(n_827),
.C(n_830),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1009),
.A2(n_825),
.B(n_924),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1009),
.A2(n_920),
.B(n_938),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1114),
.A2(n_817),
.B(n_945),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1074),
.A2(n_911),
.B(n_889),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_995),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_974),
.A2(n_911),
.B(n_880),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1055),
.A2(n_947),
.B1(n_885),
.B2(n_907),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1030),
.A2(n_845),
.B(n_850),
.C(n_938),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_977),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_1014),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1013),
.A2(n_879),
.B(n_941),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1005),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1017),
.A2(n_866),
.B(n_870),
.C(n_871),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_978),
.A2(n_909),
.B(n_935),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_986),
.A2(n_928),
.B(n_980),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_977),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_999),
.A2(n_955),
.B(n_843),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1011),
.B(n_955),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_L g1142 ( 
.A(n_971),
.B(n_882),
.C(n_847),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1011),
.B(n_970),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_983),
.A2(n_936),
.B(n_935),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_997),
.B(n_53),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_982),
.B(n_901),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1023),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1008),
.B(n_947),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_984),
.A2(n_1054),
.B(n_1069),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_984),
.A2(n_936),
.B(n_878),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1054),
.A2(n_872),
.B(n_887),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_988),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_977),
.B(n_847),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1025),
.B(n_912),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1024),
.A2(n_895),
.B(n_917),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_998),
.B(n_969),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_1100),
.A2(n_893),
.B(n_910),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1024),
.A2(n_1118),
.B(n_1090),
.Y(n_1159)
);

CKINVDCx14_ASAP7_75t_R g1160 ( 
.A(n_1003),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_973),
.A2(n_972),
.B(n_1088),
.C(n_1110),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1065),
.A2(n_903),
.B1(n_877),
.B2(n_969),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_SL g1163 ( 
.A1(n_1105),
.A2(n_966),
.B(n_964),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_1062),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1010),
.B(n_954),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_SL g1166 ( 
.A(n_979),
.B(n_962),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1090),
.A2(n_915),
.B(n_913),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1100),
.A2(n_925),
.B(n_884),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1115),
.A2(n_944),
.B1(n_953),
.B2(n_951),
.C(n_926),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1051),
.A2(n_937),
.B(n_930),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_L g1171 ( 
.A(n_1048),
.B(n_922),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_1056),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1107),
.B(n_956),
.C(n_950),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_1001),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_SL g1175 ( 
.A(n_1045),
.B(n_949),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1077),
.A2(n_954),
.B1(n_57),
.B2(n_65),
.Y(n_1176)
);

BUFx2_ASAP7_75t_R g1177 ( 
.A(n_1091),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1000),
.A2(n_57),
.B(n_59),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1026),
.A2(n_1106),
.B(n_1109),
.C(n_1018),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1087),
.B(n_71),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1040),
.A2(n_80),
.A3(n_84),
.B(n_92),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1019),
.A2(n_93),
.B(n_109),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1045),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1098),
.A2(n_111),
.B(n_117),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1020),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1102),
.A2(n_120),
.B(n_126),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1001),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_985),
.B(n_149),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1031),
.B(n_137),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1085),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1016),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1062),
.B(n_138),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1040),
.A2(n_139),
.A3(n_146),
.B(n_991),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1035),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1015),
.B(n_990),
.Y(n_1195)
);

CKINVDCx11_ASAP7_75t_R g1196 ( 
.A(n_979),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1015),
.B(n_1082),
.Y(n_1197)
);

NAND3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1083),
.B(n_1038),
.C(n_1112),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_1050),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_993),
.B(n_1047),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1073),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1039),
.B(n_1063),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_1122),
.A2(n_1105),
.B(n_1060),
.C(n_1086),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1042),
.B(n_1002),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_1050),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1076),
.A2(n_1081),
.B(n_1094),
.Y(n_1206)
);

AO32x2_ASAP7_75t_L g1207 ( 
.A1(n_1052),
.A2(n_1071),
.A3(n_991),
.B1(n_987),
.B2(n_1081),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_989),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1044),
.A2(n_986),
.B(n_1029),
.C(n_1097),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1019),
.A2(n_1117),
.B(n_1099),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1052),
.A2(n_1041),
.B(n_1037),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_994),
.A2(n_1111),
.B(n_1022),
.C(n_1096),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1095),
.A2(n_1103),
.B(n_1049),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1012),
.B(n_1121),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_996),
.A2(n_1113),
.B1(n_1059),
.B2(n_1067),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1116),
.A2(n_987),
.A3(n_1071),
.B(n_1058),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1004),
.A2(n_1057),
.A3(n_1006),
.B(n_1075),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1043),
.A2(n_1120),
.B(n_1028),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1080),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1021),
.A2(n_1070),
.A3(n_1078),
.B(n_1027),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1101),
.A2(n_1007),
.B(n_1064),
.Y(n_1221)
);

AOI211x1_ASAP7_75t_L g1222 ( 
.A1(n_1053),
.A2(n_1084),
.B(n_1079),
.C(n_992),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1036),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1061),
.A2(n_1113),
.A3(n_1093),
.B(n_1089),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1067),
.B(n_1059),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1034),
.A2(n_1068),
.B(n_1092),
.C(n_1089),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_979),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1093),
.A2(n_1104),
.B1(n_1046),
.B2(n_1033),
.Y(n_1228)
);

INVx8_ASAP7_75t_L g1229 ( 
.A(n_1032),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1032),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1033),
.A2(n_1066),
.B(n_1072),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1046),
.B(n_1104),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1033),
.A2(n_1066),
.B1(n_1072),
.B2(n_1108),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1066),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1119),
.A2(n_1072),
.B(n_1108),
.C(n_804),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_1108),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1119),
.A2(n_484),
.B1(n_511),
.B2(n_436),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1114),
.A2(n_1074),
.B(n_1013),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1062),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1040),
.A2(n_928),
.A3(n_991),
.B(n_1090),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1055),
.A2(n_775),
.B1(n_809),
.B2(n_700),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_995),
.B(n_484),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_995),
.B(n_484),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1040),
.A2(n_928),
.A3(n_991),
.B(n_1090),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_977),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1114),
.A2(n_1074),
.B(n_1013),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1055),
.A2(n_775),
.B1(n_809),
.B2(n_700),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1114),
.A2(n_1074),
.B(n_1013),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1114),
.A2(n_1074),
.B(n_1013),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1055),
.A2(n_775),
.B(n_492),
.C(n_810),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1062),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_982),
.A2(n_677),
.B1(n_732),
.B2(n_594),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1009),
.A2(n_1074),
.B(n_974),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1011),
.B(n_625),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1040),
.A2(n_928),
.A3(n_991),
.B(n_1090),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_981),
.Y(n_1256)
);

OAI22x1_ASAP7_75t_L g1257 ( 
.A1(n_1055),
.A2(n_787),
.B1(n_594),
.B2(n_484),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1114),
.A2(n_1074),
.B(n_1013),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_977),
.B(n_1011),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1115),
.A2(n_653),
.B1(n_1083),
.B2(n_1018),
.C(n_575),
.Y(n_1260)
);

INVx5_ASAP7_75t_L g1261 ( 
.A(n_977),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_976),
.A2(n_804),
.B(n_787),
.C(n_810),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_977),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_976),
.A2(n_804),
.B(n_787),
.C(n_810),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_975),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_973),
.A2(n_809),
.B(n_875),
.C(n_972),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1011),
.B(n_625),
.Y(n_1267)
);

AO32x2_ASAP7_75t_L g1268 ( 
.A1(n_1009),
.A2(n_1090),
.A3(n_1040),
.B1(n_1100),
.B2(n_1052),
.Y(n_1268)
);

AO21x1_ASAP7_75t_L g1269 ( 
.A1(n_1009),
.A2(n_923),
.B(n_1100),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_975),
.Y(n_1270)
);

NAND3x1_ASAP7_75t_L g1271 ( 
.A(n_993),
.B(n_787),
.C(n_732),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1011),
.B(n_625),
.Y(n_1272)
);

OAI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1215),
.A2(n_1185),
.B1(n_1237),
.B2(n_1145),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_SL g1274 ( 
.A(n_1228),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1133),
.B(n_1201),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1149),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1241),
.A2(n_1247),
.B1(n_1189),
.B2(n_1148),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1196),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1261),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1128),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1153),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1252),
.A2(n_1198),
.B1(n_1257),
.B2(n_1269),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1141),
.B(n_1272),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1189),
.A2(n_1195),
.B1(n_1223),
.B2(n_1124),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1259),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1187),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1265),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1125),
.A2(n_1176),
.B1(n_1206),
.B2(n_1177),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1155),
.A2(n_1190),
.B1(n_1242),
.B2(n_1243),
.Y(n_1289)
);

BUFx8_ASAP7_75t_L g1290 ( 
.A(n_1245),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1225),
.B(n_1164),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1147),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1270),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1135),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1174),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1191),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1262),
.A2(n_1264),
.B1(n_1250),
.B2(n_1179),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1194),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1146),
.A2(n_1256),
.B1(n_1208),
.B2(n_1200),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1130),
.A2(n_1154),
.B1(n_1192),
.B2(n_1143),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1172),
.A2(n_1159),
.B1(n_1184),
.B2(n_1162),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1217),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1142),
.A2(n_1138),
.B1(n_1267),
.B2(n_1254),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1197),
.A2(n_1192),
.B1(n_1204),
.B2(n_1158),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1160),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1245),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1228),
.A2(n_1188),
.B1(n_1178),
.B2(n_1150),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1168),
.A2(n_1173),
.B1(n_1245),
.B2(n_1263),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1230),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1263),
.A2(n_1140),
.B1(n_1175),
.B2(n_1271),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1172),
.A2(n_1167),
.B1(n_1214),
.B2(n_1253),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1263),
.B(n_1132),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1268),
.A2(n_1207),
.B1(n_1182),
.B2(n_1260),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1219),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1157),
.A2(n_1165),
.B1(n_1139),
.B2(n_1132),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1220),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1226),
.A2(n_1212),
.B1(n_1227),
.B2(n_1171),
.Y(n_1317)
);

INVx6_ASAP7_75t_L g1318 ( 
.A(n_1205),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1139),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1180),
.A2(n_1164),
.B1(n_1127),
.B2(n_1183),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1183),
.A2(n_1239),
.B1(n_1251),
.B2(n_1199),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1229),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1229),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1164),
.A2(n_1239),
.B1(n_1251),
.B2(n_1268),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1205),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1199),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1268),
.A2(n_1218),
.B1(n_1151),
.B2(n_1234),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1236),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1207),
.A2(n_1233),
.B1(n_1232),
.B2(n_1129),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1209),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1266),
.A2(n_1235),
.B1(n_1161),
.B2(n_1203),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1231),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1216),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1224),
.Y(n_1334)
);

INVx5_ASAP7_75t_L g1335 ( 
.A(n_1166),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1207),
.A2(n_1210),
.B1(n_1144),
.B2(n_1221),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1224),
.B(n_1255),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1152),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1216),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1224),
.B(n_1255),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1163),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1170),
.A2(n_1186),
.B1(n_1211),
.B2(n_1193),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1240),
.B(n_1255),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1238),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1137),
.A2(n_1134),
.B1(n_1126),
.B2(n_1213),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1181),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1193),
.A2(n_1244),
.B1(n_1240),
.B2(n_1181),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1193),
.A2(n_1244),
.B1(n_1240),
.B2(n_1181),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1244),
.A2(n_1131),
.B1(n_1156),
.B2(n_1249),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1246),
.A2(n_1248),
.B1(n_1258),
.B2(n_1123),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1222),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1136),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1169),
.A2(n_677),
.B1(n_541),
.B2(n_1241),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1174),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1241),
.A2(n_1247),
.B1(n_775),
.B2(n_809),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1202),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1202),
.Y(n_1357)
);

OAI21xp33_ASAP7_75t_L g1358 ( 
.A1(n_1241),
.A2(n_775),
.B(n_1055),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1202),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_1247),
.B2(n_541),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_1247),
.B2(n_541),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1202),
.Y(n_1362)
);

BUFx8_ASAP7_75t_L g1363 ( 
.A(n_1187),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1133),
.B(n_1201),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1174),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1196),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1128),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_1247),
.B2(n_541),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1261),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_541),
.B2(n_1247),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1241),
.A2(n_1247),
.B1(n_775),
.B2(n_809),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1128),
.Y(n_1372)
);

BUFx8_ASAP7_75t_SL g1373 ( 
.A(n_1128),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1227),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1133),
.B(n_1201),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1145),
.B(n_1225),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1174),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1133),
.B(n_1201),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1261),
.B(n_1175),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_1247),
.B2(n_541),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1145),
.B(n_1225),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1128),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1261),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_541),
.B2(n_1247),
.Y(n_1384)
);

INVx4_ASAP7_75t_SL g1385 ( 
.A(n_1224),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1241),
.A2(n_1247),
.B1(n_775),
.B2(n_809),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1225),
.B(n_1062),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1202),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1241),
.A2(n_677),
.B1(n_1247),
.B2(n_541),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1174),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1128),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1196),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1252),
.A2(n_677),
.B1(n_1247),
.B2(n_1241),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1261),
.B(n_1175),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1174),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1202),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1174),
.A2(n_484),
.B1(n_751),
.B2(n_511),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1174),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1202),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_SL g1400 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1289),
.C(n_1358),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1370),
.A2(n_1384),
.B1(n_1389),
.B2(n_1361),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1344),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1316),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1385),
.B(n_1335),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1302),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1346),
.A2(n_1340),
.B(n_1343),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1314),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1385),
.B(n_1335),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_L g1409 ( 
.A(n_1282),
.B(n_1288),
.C(n_1303),
.Y(n_1409)
);

CKINVDCx6p67_ASAP7_75t_R g1410 ( 
.A(n_1392),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1333),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1283),
.B(n_1275),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1337),
.B(n_1364),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1375),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1276),
.B(n_1281),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1339),
.A2(n_1329),
.B(n_1300),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1351),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1342),
.A2(n_1345),
.B(n_1350),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1288),
.A2(n_1371),
.B1(n_1355),
.B2(n_1386),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1296),
.B(n_1298),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1332),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1330),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_SL g1424 ( 
.A(n_1295),
.B(n_1397),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1344),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1329),
.A2(n_1300),
.B(n_1331),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1378),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1352),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1354),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1344),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1277),
.A2(n_1273),
.B1(n_1301),
.B2(n_1317),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1356),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1338),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1370),
.A2(n_1384),
.B1(n_1380),
.B2(n_1361),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1311),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1357),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1359),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1362),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1388),
.B(n_1396),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1348),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1348),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1327),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1327),
.Y(n_1443)
);

CKINVDCx16_ASAP7_75t_R g1444 ( 
.A(n_1372),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1334),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1399),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1341),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1274),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1376),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1291),
.B(n_1306),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1347),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1381),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1274),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1313),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1315),
.A2(n_1342),
.B(n_1313),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1324),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1324),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1350),
.A2(n_1336),
.B(n_1349),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1303),
.B(n_1284),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1315),
.A2(n_1336),
.B(n_1307),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

INVx5_ASAP7_75t_SL g1462 ( 
.A(n_1278),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1304),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1309),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1309),
.Y(n_1465)
);

AO31x2_ASAP7_75t_L g1466 ( 
.A1(n_1353),
.A2(n_1307),
.A3(n_1304),
.B(n_1282),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1299),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1284),
.A2(n_1308),
.B(n_1320),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1308),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1353),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1310),
.Y(n_1471)
);

BUFx12f_ASAP7_75t_L g1472 ( 
.A(n_1377),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1390),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1320),
.A2(n_1310),
.B(n_1321),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1379),
.A2(n_1394),
.B(n_1312),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1379),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1394),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1291),
.B(n_1387),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1360),
.A2(n_1380),
.B(n_1368),
.C(n_1389),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1285),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1360),
.A2(n_1368),
.B1(n_1393),
.B2(n_1328),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1278),
.A2(n_1366),
.B1(n_1286),
.B2(n_1374),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1306),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1279),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1279),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1369),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1404),
.B(n_1278),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1449),
.B(n_1366),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1420),
.A2(n_1366),
.B(n_1383),
.Y(n_1489)
);

AOI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1400),
.A2(n_1366),
.B1(n_1325),
.B2(n_1391),
.C(n_1280),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1452),
.B(n_1294),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1414),
.B(n_1367),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1409),
.A2(n_1383),
.B(n_1305),
.Y(n_1493)
);

INVx5_ASAP7_75t_SL g1494 ( 
.A(n_1410),
.Y(n_1494)
);

AOI211xp5_ASAP7_75t_L g1495 ( 
.A1(n_1431),
.A2(n_1435),
.B(n_1474),
.C(n_1459),
.Y(n_1495)
);

AND2x2_ASAP7_75t_SL g1496 ( 
.A(n_1435),
.B(n_1290),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1426),
.A2(n_1319),
.B1(n_1326),
.B2(n_1365),
.Y(n_1497)
);

AO22x2_ASAP7_75t_L g1498 ( 
.A1(n_1440),
.A2(n_1322),
.B1(n_1323),
.B2(n_1382),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_SL g1499 ( 
.A1(n_1447),
.A2(n_1322),
.B(n_1373),
.C(n_1363),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1433),
.B(n_1290),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1404),
.B(n_1363),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1426),
.A2(n_1318),
.B1(n_1292),
.B2(n_1395),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1408),
.B(n_1398),
.Y(n_1503)
);

NAND2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1429),
.B(n_1473),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1427),
.B(n_1436),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1415),
.B(n_1418),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1426),
.A2(n_1468),
.B(n_1455),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1433),
.B(n_1413),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1479),
.A2(n_1454),
.B(n_1463),
.C(n_1434),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1471),
.A2(n_1463),
.B1(n_1454),
.B2(n_1470),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1469),
.A2(n_1461),
.B(n_1468),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1412),
.B(n_1442),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1418),
.B(n_1421),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1421),
.B(n_1478),
.Y(n_1514)
);

OAI211xp5_ASAP7_75t_L g1515 ( 
.A1(n_1401),
.A2(n_1481),
.B(n_1468),
.C(n_1442),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1444),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1478),
.B(n_1464),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1447),
.A2(n_1484),
.B(n_1485),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1443),
.A2(n_1441),
.B1(n_1440),
.B2(n_1469),
.C(n_1461),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1443),
.B(n_1417),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1464),
.B(n_1462),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1419),
.A2(n_1458),
.B(n_1441),
.Y(n_1523)
);

AO32x1_ASAP7_75t_L g1524 ( 
.A1(n_1471),
.A2(n_1428),
.A3(n_1423),
.B1(n_1470),
.B2(n_1417),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1462),
.A2(n_1482),
.B1(n_1457),
.B2(n_1456),
.Y(n_1525)
);

AO21x1_ASAP7_75t_L g1526 ( 
.A1(n_1428),
.A2(n_1423),
.B(n_1432),
.Y(n_1526)
);

O2A1O1Ixp33_ASAP7_75t_SL g1527 ( 
.A1(n_1465),
.A2(n_1483),
.B(n_1407),
.C(n_1486),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_1460),
.B2(n_1467),
.C(n_1424),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1439),
.B(n_1446),
.Y(n_1529)
);

AND3x1_ASAP7_75t_L g1530 ( 
.A(n_1472),
.B(n_1410),
.C(n_1429),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1460),
.A2(n_1455),
.B1(n_1476),
.B2(n_1477),
.Y(n_1531)
);

O2A1O1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1460),
.A2(n_1416),
.B(n_1467),
.C(n_1476),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1422),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1419),
.A2(n_1458),
.B(n_1475),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1448),
.A2(n_1453),
.B(n_1466),
.C(n_1445),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1411),
.B(n_1453),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1520),
.B(n_1416),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1402),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1513),
.B(n_1402),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1514),
.B(n_1425),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1523),
.B(n_1517),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1505),
.B(n_1406),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1508),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1533),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1523),
.B(n_1430),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1528),
.A2(n_1519),
.B1(n_1510),
.B2(n_1490),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1534),
.B(n_1406),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1490),
.A2(n_1448),
.B(n_1450),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1526),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1528),
.A2(n_1466),
.B1(n_1480),
.B2(n_1472),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1519),
.A2(n_1466),
.B1(n_1480),
.B2(n_1445),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1521),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1518),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1498),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1508),
.B(n_1403),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1522),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1524),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1524),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1496),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1536),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1524),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1511),
.B(n_1422),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1511),
.B(n_1405),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1564)
);

NAND4xp25_ASAP7_75t_L g1565 ( 
.A(n_1546),
.B(n_1495),
.C(n_1504),
.D(n_1489),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1544),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1545),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1544),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1553),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1553),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1559),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1553),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1540),
.B(n_1535),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1542),
.B(n_1531),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1492),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_1549),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1547),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1559),
.B(n_1496),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1547),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1560),
.B(n_1529),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1547),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1549),
.A2(n_1532),
.B(n_1557),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1559),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1538),
.B(n_1498),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1547),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1546),
.A2(n_1515),
.B1(n_1509),
.B2(n_1525),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1538),
.B(n_1498),
.Y(n_1590)
);

OAI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1550),
.A2(n_1502),
.B(n_1497),
.C(n_1509),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1557),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1560),
.B(n_1552),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1569),
.Y(n_1595)
);

INVxp33_ASAP7_75t_L g1596 ( 
.A(n_1565),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1593),
.B(n_1588),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1549),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1593),
.B(n_1558),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1566),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1573),
.B(n_1556),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1567),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1559),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1592),
.B(n_1552),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1573),
.B(n_1586),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1558),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1588),
.B(n_1552),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1566),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1568),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1573),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1594),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1567),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1568),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1586),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1567),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1567),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1578),
.B(n_1558),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1573),
.B(n_1556),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1570),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1574),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1568),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1574),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1586),
.B(n_1556),
.Y(n_1626)
);

OAI33xp33_ASAP7_75t_L g1627 ( 
.A1(n_1576),
.A2(n_1561),
.A3(n_1537),
.B1(n_1563),
.B2(n_1555),
.B3(n_1543),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_SL g1628 ( 
.A(n_1565),
.B(n_1548),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1586),
.B(n_1539),
.Y(n_1629)
);

BUFx2_ASAP7_75t_SL g1630 ( 
.A(n_1580),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1613),
.B(n_1577),
.Y(n_1631)
);

OAI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1596),
.A2(n_1589),
.B(n_1578),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1613),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1613),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1571),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1613),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1602),
.B(n_1584),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1617),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1627),
.A2(n_1564),
.B1(n_1584),
.B2(n_1576),
.C(n_1583),
.Y(n_1641)
);

NOR2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1602),
.B(n_1571),
.Y(n_1642)
);

OAI33xp33_ASAP7_75t_L g1643 ( 
.A1(n_1598),
.A2(n_1577),
.A3(n_1594),
.B1(n_1579),
.B2(n_1583),
.B3(n_1587),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1628),
.B(n_1589),
.C(n_1570),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1601),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1630),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1617),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1617),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1621),
.B(n_1584),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1605),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1599),
.B(n_1577),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1621),
.B(n_1584),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1628),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1599),
.B(n_1594),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1610),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1621),
.B(n_1571),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1598),
.B(n_1584),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1607),
.B(n_1584),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1607),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1604),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1599),
.B(n_1582),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1608),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1604),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1611),
.Y(n_1666)
);

AND3x2_ASAP7_75t_L g1667 ( 
.A(n_1607),
.B(n_1503),
.C(n_1493),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1611),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1615),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1608),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1606),
.B(n_1575),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1616),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1663),
.B(n_1608),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1663),
.B(n_1620),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1633),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1633),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1632),
.B(n_1596),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1626),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1632),
.B(n_1644),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_SL g1680 ( 
.A(n_1643),
.B(n_1504),
.C(n_1473),
.Y(n_1680)
);

AOI211x1_ASAP7_75t_L g1681 ( 
.A1(n_1661),
.A2(n_1626),
.B(n_1564),
.C(n_1591),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1655),
.B(n_1606),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_1626),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1671),
.B(n_1620),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1627),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1642),
.B(n_1604),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1645),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1645),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1656),
.B(n_1597),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1646),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1637),
.B(n_1604),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1637),
.B(n_1629),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1638),
.B(n_1516),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1651),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1641),
.A2(n_1564),
.B1(n_1589),
.B2(n_1550),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1664),
.B(n_1564),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1656),
.B(n_1597),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1670),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1634),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1639),
.B(n_1597),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1651),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1650),
.B(n_1575),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1658),
.B(n_1629),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1654),
.A2(n_1585),
.B1(n_1580),
.B2(n_1575),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1660),
.B(n_1575),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1653),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1679),
.A2(n_1591),
.B1(n_1659),
.B2(n_1551),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1677),
.A2(n_1636),
.B(n_1667),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1679),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_SL g1711 ( 
.A(n_1696),
.B(n_1631),
.C(n_1634),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1675),
.Y(n_1712)
);

AOI32xp33_ASAP7_75t_L g1713 ( 
.A1(n_1685),
.A2(n_1652),
.A3(n_1648),
.B1(n_1649),
.B2(n_1640),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1682),
.B(n_1652),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1687),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_SL g1717 ( 
.A1(n_1685),
.A2(n_1638),
.B(n_1662),
.C(n_1665),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1699),
.Y(n_1718)
);

OAI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1680),
.A2(n_1658),
.B(n_1631),
.Y(n_1719)
);

OA21x2_ASAP7_75t_SL g1720 ( 
.A1(n_1681),
.A2(n_1636),
.B(n_1609),
.Y(n_1720)
);

AOI321xp33_ASAP7_75t_L g1721 ( 
.A1(n_1705),
.A2(n_1551),
.A3(n_1532),
.B1(n_1640),
.B2(n_1648),
.C(n_1649),
.Y(n_1721)
);

NAND4xp75_ASAP7_75t_L g1722 ( 
.A(n_1679),
.B(n_1530),
.C(n_1665),
.D(n_1662),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1679),
.B(n_1635),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1673),
.B(n_1684),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1678),
.B(n_1635),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1694),
.A2(n_1585),
.B1(n_1636),
.B2(n_1629),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1703),
.A2(n_1561),
.B1(n_1515),
.B2(n_1581),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1694),
.A2(n_1612),
.B1(n_1590),
.B2(n_1579),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1678),
.B(n_1612),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1674),
.B(n_1614),
.Y(n_1730)
);

AOI31xp33_ASAP7_75t_L g1731 ( 
.A1(n_1686),
.A2(n_1499),
.A3(n_1503),
.B(n_1595),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1688),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1711),
.A2(n_1706),
.B1(n_1701),
.B2(n_1697),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1710),
.B(n_1693),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1715),
.B(n_1674),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_1691),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1729),
.B(n_1683),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1723),
.Y(n_1738)
);

NAND2x1_ASAP7_75t_L g1739 ( 
.A(n_1731),
.B(n_1683),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1712),
.Y(n_1740)
);

XNOR2x1_ASAP7_75t_L g1741 ( 
.A(n_1722),
.B(n_1501),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

OAI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1708),
.A2(n_1548),
.B1(n_1554),
.B2(n_1581),
.Y(n_1743)
);

INVxp33_ASAP7_75t_L g1744 ( 
.A(n_1709),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1724),
.B(n_1689),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1710),
.A2(n_1600),
.B(n_1595),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1727),
.B(n_1689),
.Y(n_1747)
);

OAI33xp33_ASAP7_75t_L g1748 ( 
.A1(n_1732),
.A2(n_1698),
.A3(n_1702),
.B1(n_1707),
.B2(n_1695),
.B3(n_1692),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1731),
.A2(n_1713),
.B1(n_1720),
.B2(n_1719),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1716),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1730),
.A2(n_1698),
.B1(n_1612),
.B2(n_1622),
.Y(n_1751)
);

NAND2xp33_ASAP7_75t_L g1752 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1752)
);

OAI222xp33_ASAP7_75t_L g1753 ( 
.A1(n_1747),
.A2(n_1749),
.B1(n_1743),
.B2(n_1739),
.C1(n_1733),
.C2(n_1721),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1734),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1735),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1744),
.A2(n_1728),
.B(n_1690),
.C(n_1686),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1741),
.A2(n_1726),
.B(n_1700),
.Y(n_1757)
);

XNOR2x1_ASAP7_75t_L g1758 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1740),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1746),
.A2(n_1587),
.B1(n_1583),
.B2(n_1581),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1742),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1750),
.Y(n_1762)
);

NOR2xp67_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1700),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1763),
.B(n_1736),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1758),
.B(n_1737),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1755),
.B(n_1746),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_SL g1767 ( 
.A(n_1754),
.B(n_1751),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1752),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1758),
.Y(n_1769)
);

NOR2x1p5_ASAP7_75t_SL g1770 ( 
.A(n_1759),
.B(n_1748),
.Y(n_1770)
);

NAND4xp75_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1717),
.C(n_1704),
.D(n_1693),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1756),
.Y(n_1772)
);

NAND4xp25_ASAP7_75t_L g1773 ( 
.A(n_1757),
.B(n_1751),
.C(n_1499),
.D(n_1704),
.Y(n_1773)
);

NAND5xp2_ASAP7_75t_L g1774 ( 
.A(n_1769),
.B(n_1765),
.C(n_1768),
.D(n_1764),
.E(n_1756),
.Y(n_1774)
);

NOR4xp25_ASAP7_75t_L g1775 ( 
.A(n_1772),
.B(n_1753),
.C(n_1760),
.D(n_1669),
.Y(n_1775)
);

AOI222xp33_ASAP7_75t_L g1776 ( 
.A1(n_1770),
.A2(n_1669),
.B1(n_1561),
.B2(n_1572),
.C1(n_1600),
.C2(n_1622),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1766),
.A2(n_1572),
.B1(n_1603),
.B2(n_1590),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

OAI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1766),
.A2(n_1615),
.B1(n_1619),
.B2(n_1618),
.C(n_1625),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1775),
.B(n_1773),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1774),
.B(n_1771),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1776),
.A2(n_1672),
.B1(n_1653),
.B2(n_1668),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1778),
.Y(n_1783)
);

OAI211xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1777),
.A2(n_1672),
.B(n_1657),
.C(n_1668),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1779),
.B(n_1657),
.Y(n_1785)
);

OAI22x1_ASAP7_75t_L g1786 ( 
.A1(n_1783),
.A2(n_1666),
.B1(n_1615),
.B2(n_1625),
.Y(n_1786)
);

XOR2xp5_ASAP7_75t_L g1787 ( 
.A(n_1780),
.B(n_1501),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1781),
.A2(n_1666),
.B1(n_1614),
.B2(n_1609),
.C(n_1624),
.Y(n_1788)
);

NOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1784),
.B(n_1494),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1785),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1790),
.Y(n_1791)
);

NAND3x1_ASAP7_75t_L g1792 ( 
.A(n_1789),
.B(n_1494),
.C(n_1782),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1787),
.A2(n_1614),
.B1(n_1494),
.B2(n_1625),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1792),
.A2(n_1788),
.B(n_1786),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1791),
.B1(n_1793),
.B2(n_1615),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1795),
.A2(n_1625),
.B1(n_1623),
.B2(n_1619),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1795),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1797),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1796),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1618),
.B1(n_1623),
.B2(n_1619),
.C(n_1603),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1798),
.B(n_1618),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1801),
.A2(n_1618),
.B1(n_1619),
.B2(n_1623),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1802),
.B(n_1800),
.Y(n_1803)
);

XNOR2xp5_ASAP7_75t_L g1804 ( 
.A(n_1803),
.B(n_1500),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1491),
.B1(n_1500),
.B2(n_1623),
.C(n_1616),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1527),
.B(n_1488),
.C(n_1487),
.Y(n_1806)
);


endmodule