module fake_jpeg_30969_n_451 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_46),
.Y(n_138)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_53),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_54),
.A2(n_21),
.B1(n_37),
.B2(n_23),
.Y(n_114)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_61),
.Y(n_118)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_62),
.A2(n_64),
.B(n_42),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_66),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_70),
.B(n_77),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_25),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_109),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_39),
.B1(n_42),
.B2(n_23),
.Y(n_109)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_126),
.CON(n_144),
.SN(n_144)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_45),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_36),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_36),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_45),
.Y(n_135)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_59),
.A2(n_28),
.B1(n_24),
.B2(n_19),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_53),
.B1(n_61),
.B2(n_46),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_161),
.Y(n_186)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_94),
.A2(n_91),
.B1(n_90),
.B2(n_88),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_158),
.B1(n_159),
.B2(n_166),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_138),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_157),
.Y(n_181)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_102),
.B(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_162),
.Y(n_191)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_95),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_107),
.A2(n_75),
.B1(n_51),
.B2(n_71),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_72),
.B1(n_81),
.B2(n_54),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_141),
.B1(n_57),
.B2(n_105),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_40),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_69),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_169),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_87),
.B1(n_86),
.B2(n_85),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_26),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_26),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_118),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

BUFx4f_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_111),
.A2(n_28),
.B1(n_24),
.B2(n_60),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_104),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_68),
.Y(n_183)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_115),
.A2(n_83),
.B1(n_80),
.B2(n_74),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_140),
.B1(n_112),
.B2(n_96),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_194),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_118),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_198),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_142),
.B(n_76),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_123),
.B1(n_129),
.B2(n_140),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_108),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_143),
.Y(n_230)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_144),
.A2(n_128),
.B1(n_121),
.B2(n_112),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_123),
.B1(n_129),
.B2(n_177),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_144),
.B(n_160),
.C(n_161),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_209),
.A2(n_211),
.B(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_210),
.A2(n_226),
.B1(n_200),
.B2(n_207),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_146),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_222),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_163),
.B(n_179),
.C(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_163),
.B(n_157),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_217),
.A2(n_219),
.B(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_163),
.B1(n_153),
.B2(n_151),
.Y(n_219)
);

AOI32xp33_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_145),
.A3(n_154),
.B1(n_108),
.B2(n_28),
.Y(n_220)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_178),
.B(n_61),
.C(n_46),
.Y(n_222)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_16),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_231),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_147),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_204),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_20),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_172),
.B1(n_92),
.B2(n_122),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_193),
.B1(n_206),
.B2(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_20),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_234),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_195),
.B(n_198),
.C(n_187),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_237),
.B(n_259),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_226),
.B1(n_220),
.B2(n_215),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_247),
.B1(n_249),
.B2(n_252),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_196),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_242),
.B(n_234),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_193),
.B1(n_181),
.B2(n_183),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_243),
.A2(n_234),
.B1(n_215),
.B2(n_213),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_197),
.B(n_181),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_251),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_181),
.B(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_253),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_201),
.B1(n_205),
.B2(n_192),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_201),
.B1(n_199),
.B2(n_119),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_196),
.B(n_190),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_217),
.A2(n_208),
.B(n_185),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_231),
.B(n_182),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_190),
.C(n_185),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_233),
.C(n_213),
.Y(n_268)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_264),
.Y(n_295)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_281),
.B1(n_213),
.B2(n_249),
.Y(n_306)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_288),
.C(n_260),
.Y(n_307)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_225),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_273),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_279),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_211),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_285),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_287),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_188),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_209),
.C(n_213),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_256),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_289),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_209),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_251),
.C(n_281),
.Y(n_296)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_135),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_255),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_307),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_257),
.Y(n_294)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_296),
.B(n_297),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_239),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_254),
.B(n_243),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_298),
.A2(n_313),
.B(n_92),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_255),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_268),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_282),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_305),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_306),
.A2(n_319),
.B1(n_210),
.B2(n_273),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_288),
.B(n_246),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_308),
.B(n_65),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_284),
.A2(n_240),
.B1(n_245),
.B2(n_247),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_265),
.B1(n_270),
.B2(n_279),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_222),
.B(n_241),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_284),
.A2(n_283),
.B1(n_267),
.B2(n_275),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_228),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_323),
.A2(n_333),
.B1(n_312),
.B2(n_299),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_324),
.B(n_340),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_334),
.B1(n_338),
.B2(n_344),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_286),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_329),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_218),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_343),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_316),
.A2(n_263),
.B1(n_222),
.B2(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_304),
.Y(n_332)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_263),
.B1(n_212),
.B2(n_216),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_306),
.A2(n_274),
.B1(n_212),
.B2(n_292),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_176),
.C(n_170),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_326),
.C(n_339),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_337),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_319),
.A2(n_274),
.B1(n_264),
.B2(n_262),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_175),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_298),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_304),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_313),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_39),
.B1(n_20),
.B2(n_122),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_300),
.A2(n_39),
.B1(n_99),
.B2(n_170),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_327),
.B1(n_334),
.B2(n_338),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_296),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_363),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_352),
.B(n_355),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_315),
.B(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_354),
.B(n_357),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_294),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_356),
.A2(n_119),
.B1(n_73),
.B2(n_55),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_314),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_337),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_335),
.A2(n_312),
.B(n_303),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_360),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_321),
.C(n_314),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_367),
.C(n_368),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_321),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_318),
.C(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_325),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_369),
.B(n_11),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_384),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_361),
.A2(n_323),
.B(n_333),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_356),
.B(n_352),
.Y(n_394)
);

OAI321xp33_ASAP7_75t_L g374 ( 
.A1(n_366),
.A2(n_322),
.A3(n_330),
.B1(n_301),
.B2(n_311),
.C(n_299),
.Y(n_374)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_SL g376 ( 
.A1(n_355),
.A2(n_340),
.A3(n_301),
.B1(n_156),
.B2(n_63),
.C1(n_53),
.C2(n_221),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_379),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_152),
.C(n_99),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_382),
.C(n_347),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_223),
.C(n_221),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_369),
.B(n_350),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_383),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_362),
.A2(n_223),
.B1(n_119),
.B2(n_98),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_385),
.A2(n_388),
.B1(n_358),
.B2(n_359),
.Y(n_393)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_31),
.A3(n_63),
.B1(n_22),
.B2(n_12),
.C1(n_16),
.C2(n_15),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_25),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_98),
.B1(n_15),
.B2(n_12),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_365),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_395),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_402),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_396),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_375),
.A2(n_367),
.B1(n_347),
.B2(n_349),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_349),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_399),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_398),
.B(n_381),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_25),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_381),
.A2(n_22),
.B(n_12),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_401),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_11),
.Y(n_402)
);

AOI21x1_ASAP7_75t_L g403 ( 
.A1(n_370),
.A2(n_11),
.B(n_1),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_403),
.A2(n_386),
.B(n_1),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_416),
.B1(n_404),
.B2(n_410),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_380),
.C(n_371),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_408),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_382),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_411),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_386),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_413),
.B(n_389),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_371),
.C(n_373),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_395),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_412),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_418),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_419),
.A2(n_424),
.B1(n_427),
.B2(n_22),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_420),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_426),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_414),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_384),
.B(n_401),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_425),
.A2(n_0),
.B(n_2),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_390),
.Y(n_426)
);

AOI31xp67_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_399),
.A3(n_2),
.B(n_3),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_434),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_421),
.A2(n_0),
.B(n_2),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_430),
.A2(n_4),
.B(n_5),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_5),
.B(n_6),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_423),
.A2(n_2),
.B(n_4),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_433),
.A2(n_435),
.B(n_4),
.Y(n_440)
);

BUFx24_ASAP7_75t_SL g434 ( 
.A(n_417),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_22),
.B(n_38),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_440),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_38),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_441),
.B(n_442),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_443),
.B(n_429),
.Y(n_446)
);

OAI221xp5_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_447),
.B1(n_445),
.B2(n_439),
.C(n_38),
.Y(n_448)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_444),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_5),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_6),
.B1(n_7),
.B2(n_38),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_6),
.C(n_7),
.Y(n_451)
);


endmodule