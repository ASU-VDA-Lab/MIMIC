module real_aes_8625_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_316;
wire n_532;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g537 ( .A(n_1), .Y(n_537) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_3), .A2(n_39), .B1(n_165), .B2(n_479), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g144 ( .A1(n_4), .A2(n_145), .B(n_152), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_5), .B(n_138), .Y(n_528) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_7), .A2(n_244), .B(n_245), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_8), .B(n_41), .Y(n_116) );
INVx1_ASAP7_75t_L g162 ( .A(n_9), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_10), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g143 ( .A(n_11), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_12), .B(n_175), .Y(n_474) );
INVx1_ASAP7_75t_L g250 ( .A(n_13), .Y(n_250) );
INVx1_ASAP7_75t_L g532 ( .A(n_14), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_15), .B(n_139), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_16), .A2(n_748), .B1(n_749), .B2(n_752), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_16), .Y(n_752) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_17), .A2(n_138), .A3(n_172), .B1(n_495), .B2(n_499), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_18), .B(n_165), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_19), .B(n_191), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_20), .B(n_139), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_21), .A2(n_53), .B1(n_165), .B2(n_479), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_22), .B(n_145), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_23), .A2(n_79), .B1(n_165), .B2(n_175), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_24), .B(n_165), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_25), .B(n_136), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_26), .A2(n_248), .B(n_249), .C(n_251), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_27), .A2(n_77), .B1(n_750), .B2(n_751), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_27), .Y(n_751) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_29), .B(n_168), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_160), .Y(n_205) );
INVx1_ASAP7_75t_L g181 ( .A(n_31), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_32), .B(n_168), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_33), .B(n_447), .Y(n_451) );
INVx2_ASAP7_75t_L g148 ( .A(n_34), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_35), .B(n_165), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_36), .B(n_168), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_37), .A2(n_65), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_37), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_38), .A2(n_150), .B(n_155), .C(n_217), .Y(n_216) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_40), .A2(n_454), .B1(n_746), .B2(n_747), .C1(n_753), .C2(n_757), .Y(n_453) );
INVx1_ASAP7_75t_L g179 ( .A(n_42), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_43), .B(n_160), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_44), .A2(n_104), .B1(n_117), .B2(n_761), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_45), .B(n_165), .Y(n_522) );
OAI321xp33_ASAP7_75t_L g123 ( .A1(n_46), .A2(n_124), .A3(n_447), .B1(n_448), .B2(n_449), .C(n_451), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g448 ( .A(n_46), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_47), .A2(n_89), .B1(n_222), .B2(n_479), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_48), .B(n_165), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_49), .B(n_165), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_50), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_51), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_52), .B(n_145), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_54), .A2(n_63), .B1(n_165), .B2(n_175), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_55), .A2(n_155), .B1(n_175), .B2(n_177), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_56), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_57), .B(n_165), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_58), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_59), .B(n_165), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_60), .A2(n_159), .B(n_161), .C(n_164), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_61), .Y(n_268) );
INVx1_ASAP7_75t_L g153 ( .A(n_62), .Y(n_153) );
INVx1_ASAP7_75t_L g151 ( .A(n_64), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_65), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_66), .B(n_165), .Y(n_538) );
INVx1_ASAP7_75t_L g142 ( .A(n_67), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
AO32x2_ASAP7_75t_L g504 ( .A1(n_69), .A2(n_138), .A3(n_230), .B1(n_499), .B2(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g549 ( .A(n_70), .Y(n_549) );
INVx1_ASAP7_75t_L g487 ( .A(n_71), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_SL g190 ( .A1(n_72), .A2(n_164), .B(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g193 ( .A(n_73), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_74), .B(n_175), .Y(n_488) );
INVx1_ASAP7_75t_L g110 ( .A(n_75), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_76), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_77), .Y(n_750) );
INVx1_ASAP7_75t_L g261 ( .A(n_78), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_80), .A2(n_150), .B(n_155), .C(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_81), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_82), .B(n_175), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_83), .B(n_204), .Y(n_218) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_85), .B(n_191), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_86), .B(n_175), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_87), .A2(n_150), .B(n_155), .C(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g112 ( .A(n_88), .B(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g459 ( .A(n_88), .B(n_114), .Y(n_459) );
INVx2_ASAP7_75t_L g462 ( .A(n_88), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_90), .A2(n_102), .B1(n_175), .B2(n_176), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_91), .B(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_92), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_93), .A2(n_150), .B(n_155), .C(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_94), .Y(n_240) );
INVx1_ASAP7_75t_L g189 ( .A(n_95), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_96), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_97), .B(n_204), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_98), .B(n_175), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_99), .B(n_138), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_100), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_101), .A2(n_145), .B(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g762 ( .A(n_107), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g447 ( .A(n_112), .Y(n_447) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_113), .B(n_462), .Y(n_759) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g461 ( .A(n_114), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AO21x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_452), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g760 ( .A(n_121), .Y(n_760) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_124), .B(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_446), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_129), .A2(n_464), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx2_ASAP7_75t_L g446 ( .A(n_130), .Y(n_446) );
AND3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_368), .C(n_413), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_291), .C(n_332), .D(n_349), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_195), .B(n_211), .C(n_253), .Y(n_132) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_169), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_134), .B(n_196), .Y(n_195) );
NOR4xp25_ASAP7_75t_L g315 ( .A(n_134), .B(n_309), .C(n_316), .D(n_322), .Y(n_315) );
AND2x2_ASAP7_75t_L g388 ( .A(n_134), .B(n_277), .Y(n_388) );
AND2x2_ASAP7_75t_L g407 ( .A(n_134), .B(n_353), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_134), .B(n_402), .Y(n_416) );
AND2x2_ASAP7_75t_L g429 ( .A(n_134), .B(n_210), .Y(n_429) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_SL g274 ( .A(n_135), .Y(n_274) );
AND2x2_ASAP7_75t_L g281 ( .A(n_135), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g331 ( .A(n_135), .B(n_170), .Y(n_331) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_135), .B(n_277), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_135), .B(n_170), .Y(n_346) );
AND2x2_ASAP7_75t_L g355 ( .A(n_135), .B(n_280), .Y(n_355) );
BUFx2_ASAP7_75t_L g378 ( .A(n_135), .Y(n_378) );
AND2x2_ASAP7_75t_L g382 ( .A(n_135), .B(n_186), .Y(n_382) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_144), .B(n_167), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_137), .B(n_225), .Y(n_224) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_137), .B(n_499), .C(n_515), .Y(n_514) );
AO21x1_ASAP7_75t_L g552 ( .A1(n_137), .A2(n_515), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_138), .A2(n_187), .B(n_194), .Y(n_186) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_138), .A2(n_520), .B(n_528), .Y(n_519) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_140), .B(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g244 ( .A(n_145), .Y(n_244) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_146), .B(n_150), .Y(n_183) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g527 ( .A(n_147), .Y(n_527) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
INVx1_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx3_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx1_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx4_ASAP7_75t_SL g166 ( .A(n_150), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_150), .A2(n_472), .B(n_476), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_150), .A2(n_486), .B(n_489), .Y(n_485) );
BUFx3_ASAP7_75t_L g499 ( .A(n_150), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_150), .A2(n_521), .B(n_524), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_150), .A2(n_531), .B(n_535), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_158), .C(n_166), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_154), .A2(n_166), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_154), .A2(n_166), .B(n_246), .C(n_247), .Y(n_245) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_156), .Y(n_165) );
BUFx3_ASAP7_75t_L g222 ( .A(n_156), .Y(n_222) );
INVx1_ASAP7_75t_L g479 ( .A(n_156), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_159), .A2(n_477), .B(n_478), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_L g548 ( .A1(n_159), .A2(n_536), .B(n_549), .C(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx4_ASAP7_75t_L g236 ( .A(n_160), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_160), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g505 ( .A1(n_160), .A2(n_163), .B1(n_506), .B2(n_507), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_160), .A2(n_497), .B1(n_516), .B2(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_163), .B(n_193), .Y(n_192) );
INVx5_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_SL g486 ( .A1(n_164), .A2(n_204), .B(n_487), .C(n_488), .Y(n_486) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_165), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_166), .A2(n_174), .B1(n_182), .B2(n_183), .Y(n_173) );
INVx1_ASAP7_75t_L g209 ( .A(n_168), .Y(n_209) );
INVx2_ASAP7_75t_L g230 ( .A(n_168), .Y(n_230) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_168), .A2(n_243), .B(n_252), .Y(n_242) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_168), .A2(n_471), .B(n_480), .Y(n_470) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_168), .A2(n_485), .B(n_492), .Y(n_484) );
OR2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_186), .Y(n_169) );
AND2x2_ASAP7_75t_L g210 ( .A(n_170), .B(n_186), .Y(n_210) );
BUFx2_ASAP7_75t_L g284 ( .A(n_170), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_170), .A2(n_317), .B1(n_319), .B2(n_320), .Y(n_316) );
OR2x2_ASAP7_75t_L g338 ( .A(n_170), .B(n_198), .Y(n_338) );
AND2x2_ASAP7_75t_L g402 ( .A(n_170), .B(n_280), .Y(n_402) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g270 ( .A(n_171), .B(n_198), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_171), .B(n_186), .Y(n_277) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_171), .Y(n_319) );
OR2x2_ASAP7_75t_L g354 ( .A(n_171), .B(n_197), .Y(n_354) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_184), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_172), .B(n_185), .Y(n_184) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_172), .A2(n_199), .B(n_207), .Y(n_198) );
INVx2_ASAP7_75t_L g223 ( .A(n_172), .Y(n_223) );
INVx2_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_177) );
INVx2_ASAP7_75t_L g180 ( .A(n_178), .Y(n_180) );
INVx4_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_183), .A2(n_200), .B(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_183), .A2(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g273 ( .A(n_186), .Y(n_273) );
INVx3_ASAP7_75t_L g282 ( .A(n_186), .Y(n_282) );
BUFx2_ASAP7_75t_L g306 ( .A(n_186), .Y(n_306) );
AND2x2_ASAP7_75t_L g339 ( .A(n_186), .B(n_274), .Y(n_339) );
INVx1_ASAP7_75t_L g475 ( .A(n_191), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_195), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_424) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_210), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_197), .B(n_282), .Y(n_286) );
INVx1_ASAP7_75t_L g314 ( .A(n_197), .Y(n_314) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g280 ( .A(n_198), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
INVx2_ASAP7_75t_L g497 ( .A(n_204), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_204), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_204), .A2(n_546), .B(n_547), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_206), .A2(n_532), .B(n_533), .C(n_534), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_209), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_209), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g292 ( .A(n_210), .Y(n_292) );
NAND2x1_ASAP7_75t_SL g211 ( .A(n_212), .B(n_226), .Y(n_211) );
AND2x2_ASAP7_75t_L g290 ( .A(n_212), .B(n_241), .Y(n_290) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_212), .Y(n_364) );
AND2x2_ASAP7_75t_L g391 ( .A(n_212), .B(n_311), .Y(n_391) );
AND2x2_ASAP7_75t_L g399 ( .A(n_212), .B(n_361), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_212), .B(n_256), .Y(n_426) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g257 ( .A(n_213), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g275 ( .A(n_213), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g296 ( .A(n_213), .Y(n_296) );
INVx1_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_213), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g335 ( .A(n_213), .B(n_259), .Y(n_335) );
OR2x2_ASAP7_75t_L g373 ( .A(n_213), .B(n_328), .Y(n_373) );
AOI32xp33_ASAP7_75t_L g385 ( .A1(n_213), .A2(n_386), .A3(n_389), .B1(n_390), .B2(n_391), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_213), .B(n_361), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_213), .B(n_321), .Y(n_436) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_216), .B(n_223), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_220), .A2(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
INVx1_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_223), .A2(n_530), .B(n_539), .Y(n_529) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_223), .A2(n_544), .B(n_551), .Y(n_543) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g347 ( .A(n_227), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
INVx1_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
AND2x2_ASAP7_75t_L g311 ( .A(n_228), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_228), .B(n_258), .Y(n_328) );
AND2x2_ASAP7_75t_L g361 ( .A(n_228), .B(n_337), .Y(n_361) );
AND2x2_ASAP7_75t_L g398 ( .A(n_228), .B(n_259), .Y(n_398) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_229), .B(n_258), .Y(n_288) );
AND2x2_ASAP7_75t_L g295 ( .A(n_229), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g336 ( .A(n_229), .B(n_337), .Y(n_336) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .Y(n_233) );
INVx2_ASAP7_75t_L g312 ( .A(n_241), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_241), .B(n_258), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_241), .B(n_303), .Y(n_384) );
INVx1_ASAP7_75t_L g406 ( .A(n_241), .Y(n_406) );
INVx1_ASAP7_75t_L g423 ( .A(n_241), .Y(n_423) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g276 ( .A(n_242), .B(n_258), .Y(n_276) );
AND2x2_ASAP7_75t_L g298 ( .A(n_242), .B(n_259), .Y(n_298) );
INVx1_ASAP7_75t_L g337 ( .A(n_242), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_248), .B(n_250), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_248), .A2(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g534 ( .A(n_248), .Y(n_534) );
AOI221x1_ASAP7_75t_SL g253 ( .A1(n_254), .A2(n_269), .B1(n_275), .B2(n_277), .C(n_278), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_254), .A2(n_342), .B1(n_409), .B2(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
AND2x2_ASAP7_75t_L g300 ( .A(n_255), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g395 ( .A(n_255), .B(n_275), .Y(n_395) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g351 ( .A(n_256), .B(n_276), .Y(n_351) );
INVx1_ASAP7_75t_L g363 ( .A(n_257), .Y(n_363) );
AND2x2_ASAP7_75t_L g374 ( .A(n_257), .B(n_361), .Y(n_374) );
AND2x2_ASAP7_75t_L g441 ( .A(n_257), .B(n_336), .Y(n_441) );
INVx2_ASAP7_75t_L g303 ( .A(n_258), .Y(n_303) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_266), .B(n_267), .Y(n_259) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_270), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g393 ( .A(n_270), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_271), .B(n_354), .Y(n_357) );
INVx3_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_272), .A2(n_393), .B(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NOR2xp33_ASAP7_75t_SL g415 ( .A(n_275), .B(n_301), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_276), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g367 ( .A(n_276), .B(n_295), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_276), .B(n_302), .Y(n_444) );
AND2x2_ASAP7_75t_L g313 ( .A(n_277), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g380 ( .A(n_277), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_283), .B(n_287), .Y(n_278) );
NAND2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_280), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g329 ( .A(n_280), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g341 ( .A(n_280), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_280), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g365 ( .A(n_281), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_281), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_281), .B(n_284), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_284), .A2(n_323), .B(n_353), .C(n_355), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_284), .A2(n_371), .B1(n_374), .B2(n_375), .C(n_379), .Y(n_370) );
AND2x2_ASAP7_75t_L g366 ( .A(n_285), .B(n_319), .Y(n_366) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g326 ( .A(n_290), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g397 ( .A(n_290), .B(n_398), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_299), .C(n_324), .Y(n_291) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_292), .B(n_411), .C(n_412), .Y(n_410) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
OR2x2_ASAP7_75t_L g383 ( .A(n_294), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_304), .B1(n_307), .B2(n_313), .C(n_315), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_301), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_301), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_363), .B1(n_364), .B2(n_365), .Y(n_362) );
OR2x2_ASAP7_75t_L g443 ( .A(n_306), .B(n_354), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVxp67_ASAP7_75t_L g417 ( .A(n_309), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_311), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g318 ( .A(n_312), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_314), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_314), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_314), .B(n_381), .Y(n_420) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g434 ( .A(n_323), .B(n_354), .Y(n_434) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g412 ( .A(n_329), .Y(n_412) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI322xp33_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_338), .A3(n_339), .B1(n_340), .B2(n_343), .C1(n_345), .C2(n_347), .Y(n_332) );
OAI322xp33_ASAP7_75t_L g414 ( .A1(n_333), .A2(n_415), .A3(n_416), .B1(n_417), .B2(n_418), .C1(n_419), .C2(n_421), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx4_ASAP7_75t_L g348 ( .A(n_335), .Y(n_348) );
AND2x2_ASAP7_75t_L g409 ( .A(n_335), .B(n_361), .Y(n_409) );
AND2x2_ASAP7_75t_L g422 ( .A(n_335), .B(n_423), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g433 ( .A(n_338), .Y(n_433) );
INVx1_ASAP7_75t_L g411 ( .A(n_339), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g428 ( .A(n_341), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_341), .B(n_382), .Y(n_439) );
OR2x2_ASAP7_75t_L g372 ( .A(n_344), .B(n_373), .Y(n_372) );
INVxp33_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
OAI221xp5_ASAP7_75t_SL g349 ( .A1(n_348), .A2(n_350), .B1(n_352), .B2(n_356), .C(n_358), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_348), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g432 ( .A(n_348), .Y(n_432) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx3_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI322xp5_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_380), .A3(n_397), .B1(n_399), .B2(n_400), .C1(n_403), .C2(n_407), .Y(n_396) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_366), .B2(n_367), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_392), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_385), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_373), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NAND2xp33_ASAP7_75t_SL g390 ( .A(n_376), .B(n_387), .Y(n_390) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
OAI322xp33_ASAP7_75t_L g430 ( .A1(n_378), .A2(n_431), .A3(n_433), .B1(n_434), .B2(n_435), .C1(n_437), .C2(n_440), .Y(n_430) );
AOI21xp33_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_381), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_388), .B(n_436), .Y(n_445) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B(n_396), .C(n_408), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_424), .C(n_430), .D(n_442), .Y(n_413) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_444), .B(n_445), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_446), .A2(n_456), .B1(n_460), .B2(n_463), .Y(n_455) );
INVx1_ASAP7_75t_L g450 ( .A(n_447), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_451), .A2(n_453), .B(n_760), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g755 ( .A(n_459), .Y(n_755) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx6_ASAP7_75t_L g756 ( .A(n_461), .Y(n_756) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_668), .Y(n_464) );
NAND5xp2_ASAP7_75t_L g465 ( .A(n_466), .B(n_587), .C(n_602), .D(n_628), .E(n_650), .Y(n_465) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_467), .B(n_567), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_508), .B1(n_540), .B2(n_556), .C(n_557), .Y(n_467) );
NOR2xp33_ASAP7_75t_SL g468 ( .A(n_469), .B(n_500), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_469), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g744 ( .A(n_469), .Y(n_744) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_481), .Y(n_469) );
INVx1_ASAP7_75t_L g584 ( .A(n_470), .Y(n_584) );
AND2x2_ASAP7_75t_L g586 ( .A(n_470), .B(n_494), .Y(n_586) );
AND2x2_ASAP7_75t_L g596 ( .A(n_470), .B(n_493), .Y(n_596) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_470), .Y(n_614) );
INVx1_ASAP7_75t_L g624 ( .A(n_470), .Y(n_624) );
OR2x2_ASAP7_75t_L g662 ( .A(n_470), .B(n_561), .Y(n_662) );
INVx2_ASAP7_75t_L g712 ( .A(n_470), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_470), .B(n_560), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_475), .Y(n_472) );
NOR2xp67_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_483), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_483), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_SL g644 ( .A(n_483), .B(n_584), .Y(n_644) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_484), .Y(n_502) );
INVx2_ASAP7_75t_L g561 ( .A(n_484), .Y(n_561) );
OR2x2_ASAP7_75t_L g623 ( .A(n_484), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_504), .Y(n_562) );
AND2x2_ASAP7_75t_L g579 ( .A(n_493), .B(n_559), .Y(n_579) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g503 ( .A(n_494), .B(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g582 ( .A(n_494), .Y(n_582) );
AND2x2_ASAP7_75t_L g711 ( .A(n_494), .B(n_712), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_497), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_497), .A2(n_536), .B(n_537), .C(n_538), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_499), .A2(n_545), .B(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
AND2x2_ASAP7_75t_L g674 ( .A(n_501), .B(n_562), .Y(n_674) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g675 ( .A(n_502), .B(n_586), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_503), .A2(n_643), .B(n_645), .C(n_647), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_503), .B(n_643), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_503), .A2(n_573), .B1(n_716), .B2(n_717), .C(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g559 ( .A(n_504), .Y(n_559) );
INVx1_ASAP7_75t_L g595 ( .A(n_504), .Y(n_595) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_504), .Y(n_604) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .Y(n_509) );
AND2x2_ASAP7_75t_L g621 ( .A(n_510), .B(n_566), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_510), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_511), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g713 ( .A(n_511), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g745 ( .A(n_511), .Y(n_745) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
AND2x2_ASAP7_75t_L g601 ( .A(n_512), .B(n_555), .Y(n_601) );
NOR2x1_ASAP7_75t_L g610 ( .A(n_512), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g617 ( .A(n_512), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g553 ( .A(n_513), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_518), .B(n_657), .Y(n_692) );
INVx1_ASAP7_75t_SL g696 ( .A(n_518), .Y(n_696) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
INVx3_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
AND2x2_ASAP7_75t_L g566 ( .A(n_519), .B(n_543), .Y(n_566) );
AND2x2_ASAP7_75t_L g588 ( .A(n_519), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g633 ( .A(n_519), .B(n_627), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_519), .B(n_565), .Y(n_714) );
INVx2_ASAP7_75t_L g536 ( .A(n_527), .Y(n_536) );
AND2x2_ASAP7_75t_L g554 ( .A(n_529), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_529), .B(n_543), .Y(n_590) );
AND2x2_ASAP7_75t_L g626 ( .A(n_529), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_554), .Y(n_541) );
INVx1_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
AND2x2_ASAP7_75t_L g648 ( .A(n_542), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_542), .B(n_569), .Y(n_654) );
AOI21xp5_ASAP7_75t_SL g728 ( .A1(n_542), .A2(n_560), .B(n_583), .Y(n_728) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_552), .Y(n_542) );
OR2x2_ASAP7_75t_L g571 ( .A(n_543), .B(n_552), .Y(n_571) );
AND2x2_ASAP7_75t_L g618 ( .A(n_543), .B(n_555), .Y(n_618) );
INVx2_ASAP7_75t_L g627 ( .A(n_543), .Y(n_627) );
INVx1_ASAP7_75t_L g733 ( .A(n_543), .Y(n_733) );
AND2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_627), .Y(n_657) );
INVx1_ASAP7_75t_L g682 ( .A(n_552), .Y(n_682) );
AND2x2_ASAP7_75t_L g591 ( .A(n_554), .B(n_575), .Y(n_591) );
AND2x2_ASAP7_75t_L g603 ( .A(n_554), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g721 ( .A(n_554), .Y(n_721) );
INVx2_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_555), .B(n_565), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_555), .B(n_733), .Y(n_732) );
OAI21xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_562), .B(n_563), .Y(n_557) );
AND2x2_ASAP7_75t_L g664 ( .A(n_558), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g718 ( .A(n_558), .Y(n_718) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g638 ( .A(n_559), .Y(n_638) );
BUFx2_ASAP7_75t_L g737 ( .A(n_559), .Y(n_737) );
BUFx2_ASAP7_75t_L g608 ( .A(n_560), .Y(n_608) );
AND2x2_ASAP7_75t_L g710 ( .A(n_560), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g693 ( .A(n_561), .Y(n_693) );
AND2x4_ASAP7_75t_L g620 ( .A(n_562), .B(n_583), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_562), .B(n_644), .Y(n_656) );
AOI32xp33_ASAP7_75t_L g580 ( .A1(n_563), .A2(n_581), .A3(n_583), .B1(n_585), .B2(n_586), .Y(n_580) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx3_ASAP7_75t_L g569 ( .A(n_564), .Y(n_569) );
OR2x2_ASAP7_75t_L g705 ( .A(n_564), .B(n_661), .Y(n_705) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_565), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g681 ( .A(n_565), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g573 ( .A(n_566), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g585 ( .A(n_566), .B(n_575), .Y(n_585) );
INVx1_ASAP7_75t_L g706 ( .A(n_566), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_566), .B(n_681), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_572), .B(n_576), .C(n_580), .Y(n_567) );
OAI322xp33_ASAP7_75t_L g676 ( .A1(n_568), .A2(n_613), .A3(n_677), .B1(n_679), .B2(n_683), .C1(n_684), .C2(n_688), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVxp67_ASAP7_75t_L g641 ( .A(n_569), .Y(n_641) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g695 ( .A(n_571), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_571), .B(n_611), .Y(n_742) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
OR2x2_ASAP7_75t_L g720 ( .A(n_575), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_578), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g629 ( .A(n_579), .B(n_608), .Y(n_629) );
AND2x2_ASAP7_75t_L g700 ( .A(n_579), .B(n_613), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_579), .B(n_687), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_581), .A2(n_588), .B1(n_591), .B2(n_592), .C(n_597), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_581), .B(n_594), .Y(n_598) );
AND2x2_ASAP7_75t_L g686 ( .A(n_581), .B(n_687), .Y(n_686) );
AOI32xp33_ASAP7_75t_L g725 ( .A1(n_581), .A2(n_611), .A3(n_726), .B1(n_727), .B2(n_730), .Y(n_725) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_582), .B(n_618), .C(n_641), .Y(n_659) );
AND2x2_ASAP7_75t_L g685 ( .A(n_582), .B(n_678), .Y(n_685) );
INVxp67_ASAP7_75t_L g665 ( .A(n_583), .Y(n_665) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_586), .B(n_638), .Y(n_694) );
INVx2_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_586), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g673 ( .A(n_589), .Y(n_673) );
OR2x2_ASAP7_75t_L g599 ( .A(n_590), .B(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_592), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_595), .Y(n_678) );
AND2x2_ASAP7_75t_L g637 ( .A(n_596), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g683 ( .A(n_596), .Y(n_683) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_598), .A2(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g716 ( .A(n_601), .B(n_626), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B(n_615), .C(n_622), .Y(n_602) );
AND2x2_ASAP7_75t_L g646 ( .A(n_604), .B(n_614), .Y(n_646) );
INVx2_ASAP7_75t_L g661 ( .A(n_604), .Y(n_661) );
OR2x2_ASAP7_75t_L g699 ( .A(n_604), .B(n_662), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_604), .B(n_742), .Y(n_741) );
AOI211xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_607), .B(n_609), .C(n_612), .Y(n_605) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g727 ( .A1(n_609), .A2(n_704), .B(n_728), .C(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_610), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g667 ( .A(n_611), .B(n_657), .Y(n_667) );
INVx1_ASAP7_75t_L g672 ( .A(n_611), .Y(n_672) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVxp33_ASAP7_75t_L g723 ( .A(n_617), .Y(n_723) );
AND2x2_ASAP7_75t_L g702 ( .A(n_618), .B(n_681), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_623), .A2(n_685), .B(n_686), .Y(n_684) );
OAI322xp33_ASAP7_75t_L g703 ( .A1(n_625), .A2(n_704), .A3(n_705), .B1(n_706), .B2(n_707), .C1(n_709), .C2(n_713), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_635), .B2(n_639), .C(n_642), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g680 ( .A(n_633), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g724 ( .A(n_637), .Y(n_724) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_640), .B(n_660), .Y(n_726) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g689 ( .A(n_649), .B(n_657), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_655), .B2(n_657), .C(n_658), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_653), .A2(n_670), .B1(n_674), .B2(n_675), .C(n_676), .Y(n_669) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_657), .B(n_672), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_663), .B2(n_666), .Y(n_658) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx2_ASAP7_75t_SL g687 ( .A(n_662), .Y(n_687) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND5xp2_ASAP7_75t_L g668 ( .A(n_669), .B(n_690), .C(n_715), .D(n_725), .E(n_735), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_673), .Y(n_670) );
NOR4xp25_ASAP7_75t_L g743 ( .A(n_672), .B(n_678), .C(n_744), .D(n_745), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_675), .A2(n_736), .B1(n_738), .B2(n_740), .C(n_743), .Y(n_735) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g734 ( .A(n_681), .Y(n_734) );
OAI322xp33_ASAP7_75t_L g691 ( .A1(n_685), .A2(n_692), .A3(n_693), .B1(n_694), .B2(n_695), .C1(n_697), .C2(n_701), .Y(n_691) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_703), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g736 ( .A(n_711), .B(n_737), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_719) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
endmodule