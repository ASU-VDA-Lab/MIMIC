module real_jpeg_33464_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_578;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_0),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_1),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_138),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_1),
.A2(n_138),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_1),
.A2(n_138),
.B1(n_423),
.B2(n_427),
.Y(n_422)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_73),
.B1(n_197),
.B2(n_202),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_3),
.A2(n_73),
.B1(n_252),
.B2(n_256),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_4),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_4),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_4),
.B(n_140),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g432 ( 
.A1(n_4),
.A2(n_433),
.A3(n_438),
.B1(n_440),
.B2(n_445),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_4),
.A2(n_372),
.B1(n_462),
.B2(n_465),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_4),
.A2(n_40),
.B(n_498),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_5),
.A2(n_49),
.B1(n_244),
.B2(n_247),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_6),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_6),
.A2(n_101),
.B1(n_337),
.B2(n_340),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_6),
.A2(n_101),
.B1(n_234),
.B2(n_456),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_6),
.A2(n_101),
.B1(n_490),
.B2(n_494),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_7),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_9),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_10),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_10),
.A2(n_39),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_11),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_12),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B(n_582),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_13),
.B(n_583),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_14),
.Y(n_169)
);

AOI22x1_ASAP7_75t_L g185 ( 
.A1(n_14),
.A2(n_169),
.B1(n_186),
.B2(n_191),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_14),
.A2(n_169),
.B1(n_208),
.B2(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_14),
.A2(n_169),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_206),
.B1(n_207),
.B2(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_15),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_15),
.A2(n_206),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_15),
.A2(n_206),
.B1(n_449),
.B2(n_452),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_15),
.A2(n_206),
.B1(n_400),
.B2(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_17),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_17),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_17),
.A2(n_91),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_17),
.A2(n_91),
.B1(n_297),
.B2(n_302),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_18),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_18),
.Y(n_120)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_18),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_18),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_279),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_277),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_237),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_25),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_181),
.C(n_222),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_27),
.A2(n_28),
.B1(n_222),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_97),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_29),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_53),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_30),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_30),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_40),
.B1(n_47),
.B2(n_51),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_31),
.A2(n_40),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_35),
.Y(n_546)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_40),
.A2(n_47),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_40),
.A2(n_296),
.B1(n_399),
.B2(n_404),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_40),
.A2(n_489),
.B(n_498),
.Y(n_488)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_41),
.A2(n_196),
.B1(n_295),
.B2(n_305),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_41),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_41),
.A2(n_558),
.B1(n_559),
.B2(n_560),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_45),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_46),
.Y(n_500)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_66),
.B1(n_77),
.B2(n_87),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_54),
.A2(n_77),
.B1(n_87),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_54),
.A2(n_66),
.B1(n_77),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_54),
.A2(n_77),
.B1(n_448),
.B2(n_455),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_54),
.B(n_372),
.Y(n_540)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_55),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_55),
.A2(n_242),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_55),
.B(n_376),
.Y(n_471)
);

AO22x2_ASAP7_75t_SL g485 ( 
.A1(n_55),
.A2(n_242),
.B1(n_376),
.B2(n_486),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_78),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_59),
.Y(n_525)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_74),
.Y(n_529)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_76),
.Y(n_380)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_76),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_77),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_SL g470 ( 
.A1(n_77),
.A2(n_455),
.B(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_79),
.Y(n_191)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_80),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_81),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_81),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_86),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_86),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_86),
.Y(n_517)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_95),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_96),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_141),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_98),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_132),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_100),
.A2(n_110),
.B1(n_140),
.B2(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_105),
.Y(n_371)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_109),
.Y(n_270)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_109),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_110),
.B(n_133),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_110),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_124),
.Y(n_110)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_118),
.B2(n_121),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_113),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_117),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_117),
.Y(n_437)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_119),
.Y(n_255)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_119),
.Y(n_341)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_120),
.Y(n_467)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_123),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_127),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_129),
.Y(n_210)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_132),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_140),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_140),
.B(n_205),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_165),
.B1(n_172),
.B2(n_173),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_142),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_142),
.A2(n_173),
.B1(n_251),
.B2(n_260),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_142),
.A2(n_260),
.B1(n_362),
.B2(n_367),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_142),
.B(n_215),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_145),
.Y(n_249)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_149),
.Y(n_521)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_158),
.B(n_161),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_157),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_157),
.Y(n_327)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_160),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_171),
.Y(n_364)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_172),
.B(n_215),
.Y(n_342)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_182),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_204),
.C(n_211),
.Y(n_182)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_183),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_192),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_184),
.B(n_192),
.Y(n_384)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_185),
.Y(n_375)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_190),
.Y(n_451)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_193),
.Y(n_559)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g404 ( 
.A(n_194),
.Y(n_404)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_200),
.Y(n_403)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_201),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_201),
.Y(n_430)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_201),
.Y(n_497)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_204),
.B(n_212),
.Y(n_286)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_220),
.B2(n_221),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_213),
.A2(n_336),
.B(n_342),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_213),
.A2(n_342),
.B(n_461),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_219),
.Y(n_366)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g395 ( 
.A1(n_220),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_220),
.B(n_372),
.Y(n_487)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_222),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_236),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_265),
.B(n_271),
.Y(n_264)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx4f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_278),
.Y(n_277)
);

XOR2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_273),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_262),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_250),
.B(n_261),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_250),
.Y(n_261)
);

OAI211xp5_ASAP7_75t_L g527 ( 
.A1(n_242),
.A2(n_528),
.B(n_529),
.C(n_530),
.Y(n_527)
);

BUFx4f_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_266),
.B(n_333),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.C(n_276),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_346),
.B(n_579),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_343),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_282),
.B(n_343),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.C(n_291),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_284),
.B(n_352),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_331),
.C(n_334),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_292),
.A2(n_293),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_308),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_294),
.B(n_308),
.Y(n_392)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_301),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_301),
.Y(n_426)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_304),
.Y(n_493)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_320),
.B2(n_324),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx2_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_357)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx8_ASAP7_75t_L g464 ( 
.A(n_339),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_407),
.B(n_573),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_353),
.B(n_385),
.Y(n_349)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_350),
.Y(n_578)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_354),
.B(n_575),
.C(n_578),
.Y(n_574)
);

MAJx2_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.C(n_383),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_355),
.A2(n_356),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_359),
.A2(n_360),
.B1(n_383),
.B2(n_384),
.Y(n_387)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_368),
.C(n_374),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_374),
.Y(n_391)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx4f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_391),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B(n_373),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_372),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_372),
.B(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_372),
.B(n_516),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_372),
.B(n_555),
.Y(n_554)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_386),
.Y(n_577)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_387),
.Y(n_388)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_389),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.C(n_393),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_390),
.B(n_569),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_392),
.A2(n_393),
.B1(n_394),
.B2(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_392),
.Y(n_570)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.C(n_405),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_395),
.B(n_476),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_398),
.A2(n_405),
.B1(n_406),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_399),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

OAI21x1_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_564),
.B(n_571),
.Y(n_408)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_478),
.B(n_563),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_468),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_411),
.B(n_468),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_447),
.C(n_460),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_413),
.B(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_431),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_414),
.B(n_432),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_421),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_420),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_419),
.Y(n_550)
);

OAI21xp33_ASAP7_75t_L g541 ( 
.A1(n_421),
.A2(n_542),
.B(n_547),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_422),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_438),
.Y(n_446)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_460),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_448),
.Y(n_486)
);

BUFx4f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_475),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.Y(n_469)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_470),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_471),
.B(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_472),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_472),
.B(n_473),
.C(n_567),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_501),
.B(n_533),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_534),
.C(n_537),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_483),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.C(n_488),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g532 ( 
.A(n_485),
.B(n_487),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_532),
.Y(n_531)
);

INVxp33_ASAP7_75t_SL g560 ( 
.A(n_489),
.Y(n_560)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

BUFx2_ASAP7_75t_SL g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_494),
.B(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_494),
.Y(n_518)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_504),
.B2(n_531),
.Y(n_501)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_504),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_526),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_505),
.B(n_526),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_514),
.B1(n_518),
.B2(n_519),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_516),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_531),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_536),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_557),
.C(n_561),
.Y(n_537)
);

OA21x2_ASAP7_75t_SL g538 ( 
.A1(n_539),
.A2(n_551),
.B(n_556),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_540),
.B(n_541),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_542),
.Y(n_558)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_544),
.B(n_554),
.Y(n_553)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_548),
.Y(n_555)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_550),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_552),
.B(n_553),
.Y(n_551)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_568),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_568),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_577),
.Y(n_575)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);


endmodule