module real_jpeg_4796_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_1),
.A2(n_57),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_1),
.A2(n_57),
.B1(n_75),
.B2(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_52),
.B1(n_63),
.B2(n_76),
.Y(n_158)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_5),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_5),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_6),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_6),
.A2(n_132),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_6),
.A2(n_132),
.B1(n_304),
.B2(n_307),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_6),
.A2(n_126),
.B1(n_132),
.B2(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_7),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_7),
.Y(n_142)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_67),
.B1(n_83),
.B2(n_200),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_67),
.B1(n_117),
.B2(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_10),
.Y(n_153)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_10),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_83),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_11),
.A2(n_90),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_12),
.A2(n_150),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_12),
.A2(n_150),
.B1(n_166),
.B2(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_12),
.A2(n_150),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_13),
.A2(n_54),
.B1(n_195),
.B2(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_13),
.B(n_260),
.C(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_13),
.B(n_110),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_13),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_13),
.B(n_59),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_13),
.B(n_121),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_14),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_15),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_15),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_15),
.A2(n_119),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_15),
.A2(n_119),
.B1(n_221),
.B2(n_254),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_15),
.A2(n_119),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_16),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_241),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_240),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_214),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_21),
.B(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_156),
.C(n_171),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_22),
.A2(n_23),
.B1(n_156),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_93),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_24),
.B(n_94),
.C(n_155),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_72),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_25),
.B(n_72),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_26),
.A2(n_250),
.B(n_252),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_26),
.A2(n_58),
.B1(n_280),
.B2(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_26),
.A2(n_252),
.B(n_330),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_27),
.A2(n_59),
.B1(n_61),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_27),
.A2(n_59),
.B1(n_158),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_27),
.B(n_253),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_32),
.Y(n_224)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_33),
.Y(n_283)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_33),
.Y(n_349)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_53),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_40),
.Y(n_281)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_41),
.A2(n_280),
.B(n_284),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_45),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_48),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_48),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_50),
.A2(n_58),
.B(n_284),
.Y(n_390)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_56),
.Y(n_221)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_59),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_66),
.Y(n_258)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_71),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_80),
.B1(n_86),
.B2(n_91),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_73),
.Y(n_204)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_79),
.Y(n_268)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_80),
.B(n_272),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_80),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_80),
.A2(n_199),
.B1(n_342),
.B2(n_368),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_82),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_82),
.Y(n_299)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_82),
.Y(n_311)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_84),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_85),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_85),
.Y(n_306)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_87),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_159)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_88),
.Y(n_273)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_89),
.Y(n_262)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_129),
.B1(n_154),
.B2(n_155),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_94),
.Y(n_154)
);

AOI22x1_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_110),
.B1(n_115),
.B2(n_122),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_95),
.A2(n_206),
.B(n_212),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_95),
.A2(n_212),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_95),
.B(n_115),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_96),
.A2(n_123),
.B1(n_213),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_96),
.A2(n_207),
.B1(n_213),
.B2(n_361),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_110),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_101),
.Y(n_346)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_109),
.Y(n_363)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_113),
.Y(n_350)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_116),
.B(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g344 ( 
.A1(n_126),
.A2(n_255),
.A3(n_338),
.B1(n_345),
.B2(n_347),
.Y(n_344)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_143),
.B2(n_148),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_174),
.B(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_134),
.A2(n_148),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_135),
.A2(n_383),
.B(n_387),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_143)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_143),
.B(n_195),
.Y(n_366)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_153),
.Y(n_386)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_156),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_157),
.B(n_159),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_198),
.B1(n_201),
.B2(n_204),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_160),
.A2(n_164),
.B(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_160),
.A2(n_265),
.B(n_269),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_160),
.A2(n_195),
.B(n_269),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_171),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_182),
.C(n_205),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_172),
.A2(n_173),
.B1(n_205),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_175),
.B(n_177),
.Y(n_239)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_182),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_183),
.A2(n_196),
.B1(n_197),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_183),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_186),
.A3(n_187),
.B1(n_190),
.B2(n_194),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g383 ( 
.A1(n_194),
.A2(n_195),
.B(n_384),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_SL g336 ( 
.A1(n_195),
.A2(n_235),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_205),
.Y(n_400)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_213),
.A2(n_361),
.B(n_364),
.Y(n_360)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_214),
.Y(n_415)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.CI(n_230),
.CON(n_214),
.SN(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_225),
.B2(n_229),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_239),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_393),
.B(n_412),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_371),
.B(n_392),
.Y(n_243)
);

AO21x1_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_352),
.B(n_370),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_324),
.B(n_351),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_287),
.B(n_323),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_263),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_248),
.B(n_263),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_249),
.A2(n_256),
.B1(n_257),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_249),
.Y(n_321)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_277),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_264),
.B(n_278),
.C(n_286),
.Y(n_325)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_285),
.B2(n_286),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_315),
.B(n_322),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_301),
.B(n_314),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_300),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_313),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_313),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_309),
.B(n_312),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_311),
.A2(n_312),
.B(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_320),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_326),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_339),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_334),
.B2(n_335),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_334),
.C(n_339),
.Y(n_353)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_353),
.B(n_354),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_359),
.B2(n_369),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_358),
.C(n_369),
.Y(n_372)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_365),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_366),
.C(n_367),
.Y(n_377)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_372),
.B(n_373),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_380),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_374)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_375),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_378),
.C(n_380),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_388),
.B2(n_391),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_389),
.C(n_390),
.Y(n_403)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_388),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_407),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_413),
.B(n_414),
.Y(n_412)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_404),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_401),
.C(n_403),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_410),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_401),
.A2(n_402),
.B1(n_403),
.B2(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_409),
.Y(n_413)
);


endmodule