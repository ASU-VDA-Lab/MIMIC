module real_jpeg_12971_n_16 (n_5, n_4, n_8, n_0, n_12, n_358, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_358;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_68),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_3),
.B(n_82),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_3),
.B(n_63),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_3),
.B(n_46),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_4),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_46),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_4),
.B(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_27),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_4),
.B(n_63),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_7),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_7),
.B(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_7),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_7),
.B(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_7),
.B(n_54),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_68),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_8),
.B(n_63),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_8),
.B(n_46),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_8),
.B(n_27),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_8),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_31),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_12),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_12),
.B(n_68),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_13),
.B(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_63),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_13),
.B(n_68),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_13),
.B(n_82),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_13),
.B(n_46),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_13),
.B(n_31),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_13),
.B(n_35),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_14),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_14),
.B(n_82),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_14),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_14),
.B(n_54),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_14),
.B(n_63),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_14),
.B(n_31),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_31),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_15),
.B(n_27),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_15),
.B(n_54),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_149),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_148),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_20),
.B(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.C(n_108),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_21),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_77),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_22),
.A2(n_23),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_42),
.C(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_26),
.B(n_30),
.C(n_33),
.Y(n_107)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_27),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_34),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_34),
.B(n_50),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_34),
.B(n_206),
.Y(n_277)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_38),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_38),
.B(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_57),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_53),
.C(n_55),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_49),
.A2(n_55),
.B1(n_142),
.B2(n_143),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_51),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_51),
.B(n_92),
.Y(n_295)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_67),
.C(n_71),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_56),
.B1(n_67),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_53),
.A2(n_56),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_53),
.B(n_167),
.Y(n_183)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_54),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_55),
.B(n_142),
.C(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_60),
.A2(n_62),
.B1(n_139),
.B2(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_60),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_61),
.B(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_65),
.B(n_77),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_73),
.C(n_75),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_67),
.A2(n_80),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_67),
.B(n_234),
.Y(n_266)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_69),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_69),
.B(n_206),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_75),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_75),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_118),
.C(n_120),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_100),
.C(n_104),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_74),
.A2(n_75),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_75),
.B(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_83),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_78),
.B(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_81),
.A2(n_83),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_81),
.Y(n_328)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_83),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_84),
.B(n_108),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_96),
.B2(n_97),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_98),
.C(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_95),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_90),
.C(n_93),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_91),
.B(n_163),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_94),
.B(n_165),
.Y(n_273)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_106),
.B2(n_107),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_100),
.A2(n_105),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_100),
.B(n_289),
.C(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_103),
.A2(n_104),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_103),
.A2(n_104),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_104),
.B(n_227),
.C(n_229),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_113),
.C(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_121),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_147),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_136),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_133),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

AOI321xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_335),
.A3(n_345),
.B1(n_349),
.B2(n_354),
.C(n_358),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_280),
.C(n_330),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_251),
.B(n_279),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_221),
.B(n_250),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_190),
.B(n_220),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_169),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_155),
.B(n_169),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_166),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_172),
.B1(n_173),
.B2(n_181),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_217),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.CI(n_159),
.CON(n_156),
.SN(n_156)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_182),
.B2(n_189),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_181),
.C(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_177),
.C(n_180),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_187),
.A2(n_188),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_187),
.B(n_303),
.C(n_306),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_214),
.B(n_219),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_203),
.B(n_213),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_201),
.C(n_202),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_208),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_223),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_236),
.B2(n_237),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_238),
.C(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_232),
.C(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_248),
.B2(n_249),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_244),
.C(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_243),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_253),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_269),
.B2(n_278),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_268),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_268),
.C(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_266),
.C(n_267),
.Y(n_299)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_260),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.CI(n_263),
.CON(n_260),
.SN(n_260)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_269),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.CI(n_275),
.CON(n_269),
.SN(n_269)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_271),
.C(n_275),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_274),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_281),
.A2(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_312),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_312),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_300),
.C(n_311),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_299),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_292),
.C(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_296),
.C(n_298),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_301),
.B1(n_311),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_308),
.C(n_310),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_305),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_329),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_321),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_321),
.C(n_329),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_319),
.C(n_320),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_336),
.A2(n_350),
.B(n_353),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_337),
.B(n_338),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_344),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_341),
.C(n_344),
.Y(n_346)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_347),
.Y(n_354)
);


endmodule