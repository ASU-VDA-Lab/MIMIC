module fake_jpeg_2562_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_68),
.Y(n_80)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_51),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_62),
.B(n_53),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_62),
.C(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_84),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_51),
.B(n_50),
.C(n_58),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_94),
.B(n_95),
.C(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_59),
.B1(n_65),
.B2(n_56),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_57),
.B1(n_61),
.B2(n_54),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_98),
.B1(n_99),
.B2(n_73),
.Y(n_110)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_48),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_55),
.B(n_59),
.C(n_4),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_56),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_97),
.C(n_73),
.Y(n_113)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_61),
.B1(n_60),
.B2(n_4),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_60),
.B1(n_3),
.B2(n_5),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_116),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_107),
.Y(n_130)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_20),
.B1(n_39),
.B2(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_114),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_9),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_43),
.B1(n_21),
.B2(n_23),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_17),
.B(n_29),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_6),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_121),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_126),
.B(n_135),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_7),
.B(n_8),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_24),
.C(n_37),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.C(n_117),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_19),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_136),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_18),
.B1(n_36),
.B2(n_31),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_133),
.A2(n_136),
.B(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_142),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_112),
.C(n_25),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_141),
.C(n_145),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_15),
.C(n_28),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_41),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_11),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_14),
.B1(n_130),
.B2(n_135),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_152),
.A2(n_153),
.B(n_136),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_120),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_151),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_166),
.B1(n_145),
.B2(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_141),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_165),
.B(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_161),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_146),
.A3(n_150),
.B1(n_147),
.B2(n_167),
.C1(n_161),
.C2(n_140),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_160),
.Y(n_177)
);


endmodule