module fake_netlist_1_6129_n_525 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_525);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_525;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_38), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_52), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_50), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_60), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_33), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_75), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_54), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_7), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_70), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_22), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_62), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_36), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_8), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_39), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_41), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_69), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_72), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_63), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_46), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_64), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_67), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_53), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_14), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_48), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_35), .Y(n_111) );
BUFx10_ASAP7_75t_L g112 ( .A(n_82), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_81), .B(n_0), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_84), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_106), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_85), .B(n_0), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_96), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_83), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_108), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
NOR2xp33_ASAP7_75t_R g129 ( .A(n_87), .B(n_29), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_89), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_89), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_95), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_126), .B(n_91), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_114), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_117), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_126), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_114), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_115), .B(n_97), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g144 ( .A1(n_130), .A2(n_91), .B1(n_93), .B2(n_105), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_114), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_119), .B(n_98), .Y(n_147) );
OAI22xp33_ASAP7_75t_SL g148 ( .A1(n_115), .A2(n_93), .B1(n_105), .B2(n_100), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_121), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_122), .B(n_111), .Y(n_151) );
INVx1_ASAP7_75t_SL g152 ( .A(n_123), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_122), .B(n_103), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_121), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_127), .B(n_103), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_149), .B(n_128), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_147), .B(n_134), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_151), .B(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_140), .B(n_118), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_151), .B(n_127), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_135), .B(n_118), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_135), .B(n_118), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_151), .B(n_132), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_138), .A2(n_132), .B(n_131), .Y(n_178) );
NOR2xp33_ASAP7_75t_R g179 ( .A(n_139), .B(n_116), .Y(n_179) );
AND3x1_ASAP7_75t_L g180 ( .A(n_143), .B(n_131), .C(n_113), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_138), .B(n_112), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_143), .B(n_131), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_141), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_152), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_166), .B(n_155), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
NOR2xp67_ASAP7_75t_L g199 ( .A(n_185), .B(n_155), .Y(n_199) );
AOI21x1_ASAP7_75t_L g200 ( .A1(n_178), .A2(n_159), .B(n_153), .Y(n_200) );
INVx4_ASAP7_75t_SL g201 ( .A(n_162), .Y(n_201) );
INVx8_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_148), .B(n_159), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_179), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_188), .B(n_153), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_185), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_161), .A2(n_154), .B(n_156), .Y(n_213) );
OR2x6_ASAP7_75t_SL g214 ( .A(n_193), .B(n_116), .Y(n_214) );
INVx6_ASAP7_75t_L g215 ( .A(n_185), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_179), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_188), .B(n_154), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_163), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_185), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_185), .B(n_136), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_166), .B(n_130), .Y(n_221) );
AO22x1_ASAP7_75t_L g222 ( .A1(n_193), .A2(n_113), .B1(n_80), .B2(n_111), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_165), .Y(n_224) );
INVx5_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_165), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_221), .A2(n_166), .B1(n_194), .B2(n_192), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_221), .A2(n_194), .B1(n_192), .B2(n_187), .Y(n_229) );
NOR2xp33_ASAP7_75t_R g230 ( .A(n_204), .B(n_194), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_202), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_196), .B(n_188), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_196), .B(n_187), .Y(n_235) );
OAI221xp5_ASAP7_75t_L g236 ( .A1(n_216), .A2(n_189), .B1(n_192), .B2(n_164), .C(n_180), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_213), .A2(n_186), .B(n_173), .Y(n_237) );
INVx6_ASAP7_75t_L g238 ( .A(n_225), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_203), .A2(n_178), .B(n_164), .C(n_176), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_213), .A2(n_186), .B(n_176), .Y(n_240) );
AOI21xp33_ASAP7_75t_SL g241 ( .A1(n_222), .A2(n_144), .B(n_189), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_211), .B(n_188), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_202), .Y(n_243) );
NAND2xp33_ASAP7_75t_R g244 ( .A(n_220), .B(n_170), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_202), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_214), .A2(n_144), .B1(n_123), .B2(n_170), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_203), .A2(n_188), .B1(n_180), .B2(n_174), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_220), .A2(n_188), .B1(n_174), .B2(n_175), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_202), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_211), .B(n_170), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_215), .A2(n_175), .B1(n_174), .B2(n_182), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_220), .A2(n_217), .B1(n_199), .B2(n_175), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_214), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_202), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_246), .A2(n_175), .B1(n_174), .B2(n_215), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_231), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_247), .A2(n_175), .B1(n_174), .B2(n_215), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_247), .A2(n_214), .B1(n_174), .B2(n_175), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_231), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_244), .A2(n_217), .B1(n_220), .B2(n_225), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_248), .A2(n_200), .B1(n_220), .B2(n_207), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_233), .B(n_201), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_242), .B(n_190), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_253), .A2(n_236), .B1(n_228), .B2(n_229), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_241), .A2(n_222), .B1(n_148), .B2(n_167), .C(n_156), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_253), .A2(n_215), .B1(n_212), .B2(n_219), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_220), .B1(n_225), .B2(n_202), .Y(n_269) );
OAI221xp5_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_125), .B1(n_124), .B2(n_133), .C(n_167), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_249), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_125), .B1(n_133), .B2(n_124), .C(n_120), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_249), .B(n_190), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_233), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_239), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_275), .Y(n_277) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_258), .B(n_230), .C(n_254), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_261), .A2(n_240), .B(n_237), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_256), .Y(n_280) );
BUFx4f_ASAP7_75t_L g281 ( .A(n_263), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_256), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_261), .A2(n_252), .B(n_207), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_264), .B(n_200), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_275), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_263), .B(n_233), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_259), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_262), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_251), .B1(n_245), .B2(n_243), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_264), .B(n_243), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_255), .A2(n_232), .B1(n_245), .B2(n_238), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_266), .A2(n_238), .B1(n_215), .B2(n_219), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_271), .B(n_195), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_265), .B(n_195), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_265), .B(n_195), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g298 ( .A1(n_276), .A2(n_125), .B(n_133), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_276), .Y(n_300) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_277), .B(n_260), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_284), .B(n_274), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_274), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_272), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_287), .B(n_257), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_290), .A2(n_269), .B1(n_267), .B2(n_275), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_287), .B(n_263), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_278), .B(n_99), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_282), .B(n_263), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_282), .B(n_270), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
BUFx2_ASAP7_75t_SL g314 ( .A(n_277), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_290), .A2(n_270), .B1(n_268), .B2(n_238), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_283), .A2(n_207), .B(n_198), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_289), .B(n_273), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_295), .B(n_137), .Y(n_318) );
AO221x2_ASAP7_75t_L g319 ( .A1(n_293), .A2(n_88), .B1(n_110), .B2(n_109), .C(n_107), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_293), .B(n_88), .Y(n_320) );
AOI33xp33_ASAP7_75t_L g321 ( .A1(n_294), .A2(n_92), .A3(n_90), .B1(n_94), .B2(n_109), .B3(n_110), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_296), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_297), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_277), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_295), .B(n_137), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_285), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_285), .B(n_137), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_327), .B(n_281), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_291), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_304), .B(n_291), .Y(n_331) );
NOR2xp33_ASAP7_75t_R g332 ( .A(n_325), .B(n_281), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_312), .Y(n_333) );
NOR2xp33_ASAP7_75t_R g334 ( .A(n_325), .B(n_281), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_312), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_302), .B(n_297), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_304), .B(n_286), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_306), .B(n_286), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_305), .B(n_286), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_306), .B(n_292), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_315), .A2(n_283), .B(n_279), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_305), .B(n_279), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_308), .B(n_281), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_308), .B(n_90), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_309), .B(n_92), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_300), .B(n_94), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_300), .B(n_104), .Y(n_351) );
OR2x4_ASAP7_75t_L g352 ( .A(n_310), .B(n_104), .Y(n_352) );
NAND4xp75_ASAP7_75t_SL g353 ( .A(n_319), .B(n_1), .C(n_2), .D(n_3), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_319), .A2(n_298), .B1(n_107), .B2(n_101), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_299), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_322), .B(n_298), .Y(n_357) );
NAND2xp33_ASAP7_75t_SL g358 ( .A(n_327), .B(n_129), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_324), .B(n_102), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_310), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_322), .B(n_2), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_314), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_324), .B(n_323), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_319), .B(n_4), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_4), .Y(n_366) );
OR2x6_ASAP7_75t_L g367 ( .A(n_301), .B(n_238), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_311), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_318), .B(n_5), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_333), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_332), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_348), .A2(n_301), .B(n_307), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g376 ( .A(n_348), .B(n_321), .C(n_320), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_352), .A2(n_317), .B1(n_326), .B2(n_328), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
AOI31xp33_ASAP7_75t_L g379 ( .A1(n_362), .A2(n_316), .A3(n_326), .B(n_328), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_332), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_364), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_366), .A2(n_137), .B1(n_201), .B2(n_205), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_368), .B(n_6), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_225), .B1(n_219), .B2(n_212), .Y(n_385) );
AOI321xp33_ASAP7_75t_L g386 ( .A1(n_365), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_9), .C(n_10), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_9), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_330), .B(n_10), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_369), .B(n_11), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_339), .B(n_12), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_331), .B(n_12), .Y(n_391) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_349), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .C1(n_18), .C2(n_19), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_358), .A2(n_206), .B(n_208), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_336), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_351), .A2(n_137), .B1(n_129), .B2(n_168), .C(n_171), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_334), .Y(n_396) );
OA22x2_ASAP7_75t_L g397 ( .A1(n_329), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_342), .A2(n_137), .B1(n_201), .B2(n_223), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_225), .B1(n_212), .B2(n_218), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_358), .A2(n_201), .B1(n_223), .B2(n_198), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_360), .B(n_18), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_340), .B(n_19), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_341), .B(n_346), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_361), .B(n_210), .C(n_197), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_367), .A2(n_225), .B1(n_224), .B2(n_218), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
OAI32xp33_ASAP7_75t_L g408 ( .A1(n_329), .A2(n_20), .A3(n_21), .B1(n_208), .B2(n_206), .Y(n_408) );
AOI32xp33_ASAP7_75t_L g409 ( .A1(n_354), .A2(n_208), .A3(n_197), .B1(n_206), .B2(n_209), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_345), .B(n_23), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_367), .A2(n_225), .B1(n_224), .B2(n_218), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_347), .B(n_26), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_359), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_354), .A2(n_207), .B(n_198), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_355), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_356), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_359), .B(n_27), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_357), .B(n_28), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g419 ( .A1(n_353), .A2(n_201), .B1(n_183), .B2(n_168), .C1(n_171), .C2(n_181), .Y(n_419) );
NAND3xp33_ASAP7_75t_SL g420 ( .A(n_334), .B(n_224), .C(n_161), .Y(n_420) );
OAI21xp33_ASAP7_75t_SL g421 ( .A1(n_353), .A2(n_227), .B(n_197), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_404), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_382), .B(n_344), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_371), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_413), .B(n_31), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_380), .B(n_32), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_403), .B(n_34), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_416), .B(n_415), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_375), .B(n_37), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_372), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_407), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_374), .Y(n_432) );
NAND4xp25_ASAP7_75t_SL g433 ( .A(n_388), .B(n_409), .C(n_421), .D(n_387), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_414), .A2(n_227), .B1(n_209), .B2(n_197), .C(n_210), .Y(n_434) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_420), .B(n_209), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_386), .B(n_198), .C(n_207), .Y(n_436) );
NAND2xp33_ASAP7_75t_SL g437 ( .A(n_381), .B(n_226), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_373), .B(n_40), .Y(n_438) );
NOR4xp25_ASAP7_75t_SL g439 ( .A(n_397), .B(n_42), .C(n_43), .D(n_44), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_394), .B(n_45), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_396), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_378), .Y(n_442) );
OAI322xp33_ASAP7_75t_L g443 ( .A1(n_391), .A2(n_146), .A3(n_150), .B1(n_157), .B2(n_158), .C1(n_142), .C2(n_181), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_397), .Y(n_444) );
AOI321xp33_ASAP7_75t_L g445 ( .A1(n_377), .A2(n_183), .A3(n_172), .B1(n_169), .B2(n_146), .C(n_158), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_379), .B(n_47), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_379), .B(n_49), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_410), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_376), .A2(n_227), .B1(n_210), .B2(n_226), .Y(n_449) );
XNOR2xp5_ASAP7_75t_L g450 ( .A(n_390), .B(n_51), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_408), .A2(n_207), .B(n_198), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_384), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_402), .B(n_55), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_389), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_401), .B(n_56), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_383), .B(n_57), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_398), .B(n_59), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_405), .B(n_61), .Y(n_458) );
AOI321xp33_ASAP7_75t_L g459 ( .A1(n_385), .A2(n_412), .A3(n_417), .B1(n_386), .B2(n_418), .C(n_395), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_376), .B(n_65), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_392), .B(n_66), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_419), .B(n_198), .C(n_207), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_399), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_423), .B(n_411), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_442), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_431), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_442), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_445), .B(n_419), .C(n_400), .Y(n_468) );
XNOR2x1_ASAP7_75t_L g469 ( .A(n_441), .B(n_406), .Y(n_469) );
AOI211xp5_ASAP7_75t_L g470 ( .A1(n_433), .A2(n_393), .B(n_226), .C(n_158), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_452), .B(n_68), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_428), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g473 ( .A1(n_444), .A2(n_226), .B(n_177), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_452), .Y(n_474) );
AOI21xp33_ASAP7_75t_SL g475 ( .A1(n_447), .A2(n_73), .B(n_74), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_424), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g477 ( .A1(n_463), .A2(n_112), .B1(n_226), .B2(n_177), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_422), .B(n_76), .Y(n_478) );
AOI32xp33_ASAP7_75t_L g479 ( .A1(n_432), .A2(n_142), .A3(n_150), .B1(n_157), .B2(n_177), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_454), .Y(n_480) );
AOI31xp33_ASAP7_75t_L g481 ( .A1(n_450), .A2(n_172), .A3(n_169), .B(n_150), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_430), .Y(n_482) );
OA22x2_ASAP7_75t_L g483 ( .A1(n_463), .A2(n_169), .B1(n_177), .B2(n_157), .Y(n_483) );
XOR2xp5_ASAP7_75t_L g484 ( .A(n_427), .B(n_226), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_429), .A2(n_191), .B1(n_112), .B2(n_142), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_448), .B(n_191), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_422), .B(n_191), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_446), .B(n_191), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_466), .B(n_460), .Y(n_489) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_464), .B(n_429), .Y(n_490) );
NOR2xp33_ASAP7_75t_R g491 ( .A(n_480), .B(n_437), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_472), .B(n_434), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_476), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_482), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_474), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_470), .A2(n_449), .B1(n_435), .B2(n_462), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_473), .A2(n_461), .B1(n_436), .B2(n_437), .C1(n_453), .C2(n_425), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_469), .Y(n_498) );
NAND2xp33_ASAP7_75t_R g499 ( .A(n_475), .B(n_439), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_471), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_470), .A2(n_434), .B(n_443), .C(n_455), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_465), .B(n_440), .Y(n_502) );
NAND2xp33_ASAP7_75t_SL g503 ( .A(n_473), .B(n_456), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_467), .B(n_438), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_SL g505 ( .A1(n_479), .A2(n_458), .B(n_426), .C(n_457), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_483), .B(n_451), .Y(n_506) );
AOI21xp33_ASAP7_75t_SL g507 ( .A1(n_481), .A2(n_459), .B(n_451), .Y(n_507) );
AOI21xp33_ASAP7_75t_SL g508 ( .A1(n_468), .A2(n_477), .B(n_484), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_468), .A2(n_182), .B1(n_184), .B2(n_486), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_488), .A2(n_184), .B1(n_487), .B2(n_485), .C(n_478), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_464), .A2(n_444), .B(n_470), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_498), .B(n_495), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_491), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_489), .B(n_490), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_511), .A2(n_503), .B(n_506), .Y(n_515) );
NOR4xp25_ASAP7_75t_L g516 ( .A(n_501), .B(n_500), .C(n_493), .D(n_494), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_512), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_515), .B(n_508), .C(n_507), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_513), .A2(n_490), .B1(n_497), .B2(n_509), .Y(n_519) );
AOI22xp33_ASAP7_75t_R g520 ( .A1(n_517), .A2(n_513), .B1(n_516), .B2(n_512), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_519), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_521), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_520), .A2(n_518), .B1(n_514), .B2(n_492), .Y(n_523) );
AOI322xp5_ASAP7_75t_L g524 ( .A1(n_522), .A2(n_500), .A3(n_496), .B1(n_510), .B2(n_504), .C1(n_502), .C2(n_499), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_524), .A2(n_523), .B(n_505), .Y(n_525) );
endmodule