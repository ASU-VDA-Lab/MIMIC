module fake_jpeg_18997_n_293 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_265;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_23),
.B1(n_31),
.B2(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_19),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_33),
.B(n_27),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_22),
.C(n_20),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_47),
.B1(n_29),
.B2(n_14),
.Y(n_56)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_23),
.B1(n_14),
.B2(n_19),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_29),
.B1(n_23),
.B2(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_60),
.B1(n_66),
.B2(n_46),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_33),
.B(n_34),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_35),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_35),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_32),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_32),
.B1(n_34),
.B2(n_28),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_82),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_59),
.B1(n_52),
.B2(n_62),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_60),
.B1(n_66),
.B2(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_88),
.Y(n_89)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_54),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_65),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_64),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_106),
.B1(n_68),
.B2(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_61),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_123),
.B1(n_115),
.B2(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_115),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_126),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_87),
.C(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_58),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_128),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_68),
.B1(n_87),
.B2(n_56),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_125),
.B1(n_41),
.B2(n_46),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_107),
.Y(n_133)
);

OAI22x1_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_58),
.B1(n_38),
.B2(n_47),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_58),
.B1(n_42),
.B2(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_86),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_42),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_42),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_30),
.B(n_43),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_142),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_155),
.B1(n_159),
.B2(n_129),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_30),
.Y(n_175)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_49),
.B1(n_132),
.B2(n_59),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_149),
.B1(n_153),
.B2(n_158),
.Y(n_179)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_100),
.B(n_98),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_128),
.B(n_1),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_18),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_10),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_92),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_95),
.B1(n_49),
.B2(n_41),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_95),
.B1(n_78),
.B2(n_41),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_22),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_44),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_12),
.B(n_22),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_16),
.B(n_12),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_49),
.B1(n_130),
.B2(n_45),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_114),
.A2(n_45),
.B1(n_34),
.B2(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_116),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_146),
.B(n_118),
.C(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_172),
.B1(n_159),
.B2(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_176),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_140),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_44),
.B(n_45),
.C(n_30),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_44),
.C(n_30),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_185),
.C(n_143),
.Y(n_197)
);

BUFx8_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_20),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_184),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_20),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_44),
.C(n_20),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_136),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_45),
.B1(n_25),
.B2(n_21),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_145),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_175),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_154),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_144),
.B(n_156),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_8),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_204),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_45),
.C(n_25),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_45),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_24),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_8),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_179),
.B1(n_167),
.B2(n_178),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_212),
.B1(n_222),
.B2(n_21),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_167),
.B1(n_172),
.B2(n_170),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_167),
.B1(n_176),
.B2(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_172),
.B(n_174),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_226),
.B(n_194),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_221),
.B(n_191),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_0),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_7),
.B(n_11),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_197),
.C(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_229),
.C(n_235),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_187),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_240),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_187),
.C(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_205),
.B1(n_203),
.B2(n_195),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_232),
.B(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_218),
.B1(n_209),
.B2(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_206),
.C(n_25),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_21),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_24),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_11),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_241),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_218),
.B1(n_208),
.B2(n_220),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_227),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_24),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_221),
.B1(n_225),
.B2(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_228),
.C(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_263),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_260),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_250),
.A2(n_238),
.B1(n_240),
.B2(n_13),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_262),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_273),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_243),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_274),
.C(n_262),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_247),
.C(n_16),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_0),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_271),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_276),
.B(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_2),
.C(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_281),
.A2(n_266),
.B(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_280),
.C(n_5),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_285),
.C(n_5),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_4),
.C(n_5),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_4),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_4),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_6),
.B(n_276),
.Y(n_293)
);


endmodule