module real_jpeg_5245_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_1),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_1),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_1),
.B(n_161),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_2),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_2),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_2),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_2),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_4),
.Y(n_307)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_6),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_6),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_6),
.B(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_7),
.Y(n_335)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_8),
.Y(n_174)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_8),
.Y(n_244)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_10),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_10),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_10),
.B(n_52),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_10),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_10),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_10),
.B(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_11),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_12),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_12),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_12),
.B(n_146),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_12),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_12),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_12),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_13),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_13),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_13),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_13),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_13),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_13),
.B(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_14),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_14),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_14),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_14),
.B(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_15),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_220),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_219),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_177),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_19),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_19),
.B(n_223),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_19),
.B(n_223),
.Y(n_422)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_77),
.CI(n_136),
.CON(n_19),
.SN(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_22),
.B(n_41),
.C(n_62),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.C(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_28),
.Y(n_144)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_29),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_30),
.B(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_35),
.Y(n_268)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_40),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_42),
.A2(n_43),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_43),
.B(n_50),
.C(n_61),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_43),
.B(n_110),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_43),
.B(n_110),
.Y(n_371)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_47),
.Y(n_148)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_61),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_54),
.Y(n_288)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_55),
.Y(n_322)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_60),
.Y(n_295)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_60),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_75),
.B2(n_76),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_63),
.B(n_152),
.C(n_155),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_63),
.B(n_69),
.C(n_72),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_63),
.A2(n_75),
.B1(n_152),
.B2(n_392),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_67),
.Y(n_325)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_72),
.B1(n_82),
.B2(n_87),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_71),
.A2(n_72),
.B1(n_260),
.B2(n_261),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_82),
.C(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_72),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_105),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_78),
.B(n_106),
.C(n_125),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_93),
.C(n_103),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_79),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_88),
.B2(n_92),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_82),
.B(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_82),
.A2(n_87),
.B1(n_241),
.B2(n_242),
.Y(n_365)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_85),
.Y(n_332)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g263 ( 
.A(n_86),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_89),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_90),
.Y(n_293)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_91),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_93),
.B(n_103),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_100),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_100),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_100),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_102),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_125),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_118),
.C(n_121),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_116),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_109),
.A2(n_110),
.B1(n_116),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_112),
.Y(n_312)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_112),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_113),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_113),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_150),
.Y(n_149)
);

OR2x2_ASAP7_75t_SL g183 ( 
.A(n_115),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_116),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_121),
.Y(n_176)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_134),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_128),
.B(n_132),
.C(n_135),
.Y(n_209)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_132),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_132),
.A2(n_134),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_158),
.C(n_175),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_137),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_151),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_138),
.B(n_151),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_140),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_149),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_141),
.A2(n_149),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_145),
.B(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_149),
.Y(n_232)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_152),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_155),
.B(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_156),
.B(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_156),
.B(n_325),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_175),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.C(n_171),
.Y(n_158)
);

FAx1_ASAP7_75t_L g250 ( 
.A(n_159),
.B(n_166),
.CI(n_171),
.CON(n_250),
.SN(n_250)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_159),
.A2(n_160),
.B(n_164),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_172),
.B(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_204),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_192),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_182),
.A2(n_183),
.B1(n_236),
.B2(n_363),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_235),
.C(n_236),
.Y(n_234)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_203),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_251),
.B(n_422),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.C(n_228),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_224),
.B(n_226),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_228),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_245),
.C(n_250),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_229),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.C(n_239),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_230),
.B(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_234),
.A2(n_239),
.B1(n_240),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_234),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_235),
.B(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_236),
.Y(n_363)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_245),
.B(n_250),
.Y(n_408)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g424 ( 
.A(n_250),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_403),
.B(n_418),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_383),
.B(n_402),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_356),
.B(n_382),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_314),
.B(n_355),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_298),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_257),
.B(n_298),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_270),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_258),
.B(n_271),
.C(n_285),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_259),
.B(n_265),
.C(n_269),
.Y(n_369)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_285),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.C(n_282),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_272),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_273),
.B(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_278),
.B1(n_282),
.B2(n_283),
.Y(n_300)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_286),
.B(n_290),
.C(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_313),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_301),
.A2(n_302),
.B1(n_313),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_304),
.B1(n_308),
.B2(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_349),
.B(n_354),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_336),
.B(n_348),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_327),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_327),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_323),
.C(n_326),
.Y(n_350)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_333),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_328),
.A2(n_329),
.B1(n_333),
.B2(n_334),
.Y(n_346)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_344),
.B(n_347),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_345),
.B(n_346),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_351),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_358),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_367),
.B2(n_368),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_369),
.C(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_365),
.C(n_366),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_381),
.Y(n_370)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_377),
.B2(n_380),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_380),
.C(n_381),
.Y(n_387)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_377),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_401),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_401),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_395),
.B2(n_400),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_396),
.C(n_397),
.Y(n_413)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_390),
.C(n_393),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_393),
.B2(n_394),
.Y(n_388)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_390),
.Y(n_394)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_395),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_414),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_413),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_410),
.C(n_411),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_420),
.B(n_421),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_416),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);


endmodule