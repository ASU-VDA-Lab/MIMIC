module real_jpeg_21863_n_17 (n_8, n_0, n_2, n_10, n_9, n_350, n_12, n_349, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_350;
input n_12;
input n_349;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_286;
wire n_166;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_53),
.B1(n_56),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_0),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_0),
.A2(n_72),
.B1(n_73),
.B2(n_96),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_0),
.A2(n_24),
.B1(n_26),
.B2(n_96),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_72),
.B1(n_73),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_1),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_1),
.A2(n_53),
.B1(n_56),
.B2(n_113),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_113),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_113),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_2),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_2),
.A2(n_23),
.B1(n_72),
.B2(n_73),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_2),
.A2(n_23),
.B1(n_53),
.B2(n_56),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_56),
.B(n_68),
.C(n_93),
.D(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_3),
.B(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_52),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_114),
.B(n_116),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_33),
.B(n_49),
.C(n_151),
.D(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_3),
.B(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_37),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_32),
.B(n_34),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_132),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_72),
.B1(n_73),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_4),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_4),
.A2(n_53),
.B1(n_56),
.B2(n_163),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_163),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_163),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_36),
.B1(n_53),
.B2(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_5),
.A2(n_36),
.B1(n_72),
.B2(n_73),
.Y(n_242)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_7),
.B(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_9),
.A2(n_53),
.B1(n_56),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_9),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_9),
.A2(n_72),
.B1(n_73),
.B2(n_108),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_108),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_108),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_10),
.A2(n_53),
.B1(n_56),
.B2(n_65),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_65),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_12),
.A2(n_53),
.B1(n_56),
.B2(n_63),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_63),
.Y(n_269)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_16),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_21),
.B(n_43),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_22),
.A2(n_27),
.B1(n_37),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_24),
.A2(n_29),
.B(n_132),
.C(n_196),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_35),
.B(n_37),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_27),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_27),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_28),
.A2(n_31),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_28),
.A2(n_31),
.B1(n_223),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_28),
.A2(n_214),
.B(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_28),
.A2(n_31),
.B1(n_62),
.B2(n_297),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_31),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_31),
.A2(n_224),
.B(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_37),
.B(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_82),
.B(n_347),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_77),
.C(n_79),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_44),
.A2(n_45),
.B1(n_342),
.B2(n_344),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_60),
.C(n_66),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_46),
.A2(n_47),
.B1(n_66),
.B2(n_322),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_48),
.A2(n_58),
.B1(n_174),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_48),
.A2(n_209),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_48),
.A2(n_57),
.B1(n_58),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_52),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_49),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_49),
.A2(n_52),
.B1(n_250),
.B2(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_49),
.A2(n_52),
.B1(n_269),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_51),
.Y(n_159)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_53),
.B(n_55),
.Y(n_158)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_56),
.A2(n_151),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_58),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_58),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_58),
.A2(n_175),
.B(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_60),
.A2(n_61),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_66),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_66),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_75),
.B(n_76),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_67),
.A2(n_75),
.B1(n_107),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_67),
.A2(n_149),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_67),
.A2(n_75),
.B1(n_206),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_67),
.A2(n_75),
.B1(n_235),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_67),
.A2(n_75),
.B1(n_244),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_68),
.A2(n_71),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

CKINVDCx9p33_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_72),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_73),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_75),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_75),
.A2(n_109),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_76),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_343),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_77),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_340),
.B(n_346),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_313),
.A3(n_333),
.B1(n_338),
.B2(n_339),
.C(n_349),
.Y(n_83)
);

AOI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_261),
.A3(n_301),
.B1(n_307),
.B2(n_312),
.C(n_350),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_217),
.C(n_257),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_189),
.B(n_216),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_168),
.B(n_188),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_143),
.B(n_167),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_119),
.B(n_142),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_101),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_91),
.B(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_106),
.C(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_114),
.B(n_116),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_114),
.A2(n_115),
.B1(n_162),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_114),
.A2(n_165),
.B1(n_179),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_114),
.A2(n_199),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_114),
.A2(n_115),
.B1(n_233),
.B2(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_114),
.A2(n_232),
.B(n_242),
.Y(n_274)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_123),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_132),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_129),
.B(n_141),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_127),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_136),
.B(n_140),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_161),
.B(n_164),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_156),
.B2(n_166),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_155),
.C(n_166),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_170),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_184),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_185),
.C(n_186),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_183),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_180),
.C(n_181),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_191),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_203),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_193),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_202),
.C(n_203),
.Y(n_258)
);

AOI22x1_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_198),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_211),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_218),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_237),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_219),
.B(n_237),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.C(n_236),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_236),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_255),
.B2(n_256),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_245),
.C(n_256),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_243),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_251),
.C(n_254),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_255),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_258),
.B(n_259),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_279),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_262),
.B(n_279),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_272),
.C(n_278),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_272),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_272)
);

AOI22x1_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_274),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_292),
.B(n_296),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_275),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_275),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_299),
.B2(n_300),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_290),
.B2(n_291),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_291),
.C(n_300),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_287),
.B(n_289),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_287),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_288),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_289),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_289),
.A2(n_315),
.B1(n_324),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_298),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_294),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_308),
.B(n_311),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_326),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.C(n_325),
.Y(n_314)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_316),
.A2(n_317),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_322),
.C(n_323),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_328),
.C(n_332),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_320),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_334),
.B(n_335),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_345),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_342),
.Y(n_344)
);


endmodule