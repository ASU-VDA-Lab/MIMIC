module fake_jpeg_12217_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_9),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_71),
.B1(n_53),
.B2(n_70),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_66),
.B1(n_52),
.B2(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_0),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_69),
.Y(n_88)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_73),
.Y(n_100)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_61),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_98),
.B(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_63),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_R g95 ( 
.A(n_77),
.B(n_66),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_49),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_71),
.B1(n_56),
.B2(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_31),
.Y(n_133)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_117),
.Y(n_132)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_109),
.Y(n_121)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_97),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_110),
.C(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_1),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_51),
.A3(n_74),
.B1(n_56),
.B2(n_59),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_1),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_24),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_3),
.Y(n_127)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_51),
.B1(n_4),
.B2(n_6),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_137),
.B1(n_36),
.B2(n_37),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_25),
.C(n_43),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_23),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_7),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_7),
.B(n_8),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_32),
.B(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_21),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_11),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_38),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_137)
);

AOI22x1_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_138)
);

AO21x1_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_118),
.B(n_27),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_126),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_34),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_151),
.C(n_153),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_45),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_128),
.B1(n_139),
.B2(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_140),
.Y(n_163)
);

OAI321xp33_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_164),
.A3(n_165),
.B1(n_159),
.B2(n_151),
.C(n_141),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_148),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_142),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_159),
.C(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_162),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_122),
.C(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_152),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_146),
.Y(n_172)
);


endmodule