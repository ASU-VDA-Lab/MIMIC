module real_jpeg_7494_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_0),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_0),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_0),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_0),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_0),
.B(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_32),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_2),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_2),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_2),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2x1_ASAP7_75t_SL g84 ( 
.A(n_3),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_3),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_3),
.B(n_134),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_3),
.B(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_4),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_4),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_5),
.Y(n_512)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_7),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_7),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_7),
.B(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_8),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_8),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g427 ( 
.A(n_8),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_11),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_11),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_11),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_11),
.B(n_63),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_11),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_11),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_11),
.B(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_13),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_13),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_13),
.B(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_13),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_13),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_13),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_13),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_13),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_14),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_14),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_14),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_14),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_14),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_14),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_15),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_15),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_15),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_15),
.B(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_16),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_17),
.Y(n_171)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_17),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_507),
.B(n_509),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_75),
.B(n_110),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_21),
.B(n_75),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_35),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_24),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_24),
.A2(n_35),
.B1(n_48),
.B2(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_24),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_28),
.Y(n_221)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_29),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_30),
.A2(n_31),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_30),
.A2(n_31),
.B1(n_335),
.B2(n_341),
.Y(n_334)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_31),
.B(n_336),
.C(n_340),
.Y(n_489)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_35),
.A2(n_58),
.B1(n_65),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_35),
.A2(n_58),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_35),
.B(n_155),
.C(n_160),
.Y(n_258)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_37),
.Y(n_280)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_38),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_38),
.Y(n_338)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_38),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_66),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_39),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_39),
.B(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_43),
.A2(n_44),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_43),
.A2(n_44),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_43),
.B(n_349),
.C(n_356),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_44),
.B(n_314),
.C(n_318),
.Y(n_347)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_46),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_48),
.B(n_231),
.C(n_236),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_49),
.A2(n_50),
.B1(n_79),
.B2(n_80),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_65),
.C(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_51),
.Y(n_330)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_52),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.C(n_64),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_55),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_65),
.C(n_69),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_104),
.B1(n_122),
.B2(n_126),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_65),
.B(n_122),
.C(n_127),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_65),
.A2(n_104),
.B1(n_484),
.B2(n_485),
.Y(n_483)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_67),
.Y(n_219)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_67),
.Y(n_380)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_68),
.Y(n_257)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_68),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_70),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_69),
.A2(n_70),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_69),
.B(n_196),
.C(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_74),
.Y(n_208)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_74),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_105),
.C(n_106),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_76),
.B(n_105),
.CI(n_106),
.CON(n_504),
.SN(n_504)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_93),
.C(n_101),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_77),
.B(n_495),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_88),
.C(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_79),
.A2(n_80),
.B1(n_137),
.B2(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_79),
.A2(n_80),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_133),
.C(n_137),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_80),
.B(n_196),
.C(n_329),
.Y(n_488)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_93),
.B(n_101),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_94),
.Y(n_479)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_97),
.A2(n_98),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_98),
.B(n_142),
.C(n_244),
.Y(n_318)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_100),
.B(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_503),
.B(n_506),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_471),
.B(n_500),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_321),
.B(n_357),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_288),
.B(n_320),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_259),
.B(n_287),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_116),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_223),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_117),
.B(n_223),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_175),
.C(n_209),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_118),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_151),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_119),
.B(n_152),
.C(n_162),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_132),
.C(n_140),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_120),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_132),
.A2(n_140),
.B1(n_141),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_132),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_133),
.B(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_142),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_142),
.A2(n_147),
.B1(n_148),
.B2(n_246),
.Y(n_281)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_145),
.Y(n_424)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_146),
.Y(n_368)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_162),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_156),
.B(n_196),
.Y(n_374)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_158),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_162),
.Y(n_516)
);

FAx1_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.CI(n_172),
.CON(n_162),
.SN(n_162)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_164),
.B(n_165),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_163),
.B(n_167),
.C(n_172),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_173),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_175),
.B(n_209),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_191),
.C(n_193),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_176),
.A2(n_191),
.B1(n_192),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_180),
.C(n_184),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_178),
.B(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_178),
.B(n_417),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_190),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_183),
.A2(n_184),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_184),
.B(n_244),
.C(n_303),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_188),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_189),
.Y(n_373)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_193),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.C(n_205),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_194),
.A2(n_195),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_196),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_196),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_196),
.A2(n_296),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_200),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_459)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_203),
.Y(n_404)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_222),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_212),
.C(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_218),
.C(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_218),
.A2(n_336),
.B1(n_339),
.B2(n_340),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_218),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_226),
.C(n_247),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_247),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_240),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_229),
.C(n_240),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_243),
.A2(n_244),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_243),
.A2(n_244),
.B1(n_365),
.B2(n_366),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_244),
.B(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_255),
.C(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_285),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_260),
.B(n_285),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.C(n_282),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_261),
.A2(n_262),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_265),
.B(n_282),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_281),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_266),
.B(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_269),
.B(n_281),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_276),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_270),
.A2(n_271),
.B1(n_276),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_273),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_276),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_277),
.B(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_277),
.B(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_289),
.B(n_321),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_322),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_291),
.B(n_322),
.Y(n_470)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_306),
.CI(n_319),
.CON(n_291),
.SN(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_294),
.B(n_295),
.C(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_302),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_323),
.B(n_325),
.C(n_342),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_342),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_332),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_326),
.B(n_333),
.C(n_334),
.Y(n_480)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_335),
.Y(n_341)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_343),
.B(n_347),
.C(n_348),
.Y(n_490)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

AO22x1_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_353),
.Y(n_356)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

OAI31xp33_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_467),
.A3(n_468),
.B(n_470),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_461),
.B(n_466),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_448),
.B(n_460),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_406),
.B(n_447),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_392),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_362),
.B(n_392),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_375),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_363),
.B(n_376),
.C(n_389),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_364),
.B(n_370),
.C(n_374),
.Y(n_456)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_374),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_389),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_381),
.C(n_386),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_377),
.B(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_381),
.A2(n_382),
.B1(n_386),
.B2(n_387),
.Y(n_394)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_405),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_393),
.B(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_395),
.A2(n_396),
.B1(n_405),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_398),
.B1(n_402),
.B2(n_403),
.Y(n_418)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_401),
.Y(n_432)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_441),
.B(n_446),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_428),
.B(n_440),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_419),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_419),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_418),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_415),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_415),
.C(n_418),
.Y(n_442)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_421),
.B1(n_425),
.B2(n_426),
.Y(n_438)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_436),
.B(n_439),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

INVx5_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_438),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_443),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_450),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_454),
.B2(n_455),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_456),
.C(n_457),
.Y(n_465)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_465),
.Y(n_466)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_496),
.Y(n_471)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_472),
.A2(n_501),
.B(n_502),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_491),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_491),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_481),
.C(n_490),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_481),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_480),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_477),
.C(n_480),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_486),
.B2(n_487),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_488),
.C(n_489),
.Y(n_493)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_499),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_491),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_493),
.CI(n_494),
.CON(n_491),
.SN(n_491)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_493),
.C(n_494),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_498),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_505),
.Y(n_506)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_504),
.Y(n_514)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_508),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_512),
.Y(n_509)
);

BUFx12f_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);


endmodule