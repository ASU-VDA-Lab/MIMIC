module fake_jpeg_23645_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_18),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_18),
.B1(n_29),
.B2(n_26),
.Y(n_48)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_24),
.B(n_15),
.Y(n_54)
);

BUFx12f_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_78),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2x1_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_24),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_53),
.B(n_25),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_58),
.Y(n_91)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_18),
.B1(n_29),
.B2(n_31),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_42),
.B1(n_41),
.B2(n_52),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_101),
.C(n_82),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_102),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_48),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_106),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_63),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_29),
.B1(n_20),
.B2(n_26),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_26),
.B1(n_20),
.B2(n_75),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_57),
.B1(n_52),
.B2(n_40),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_84),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_45),
.B1(n_46),
.B2(n_39),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_111),
.B(n_90),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_64),
.A3(n_78),
.B1(n_65),
.B2(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_37),
.C(n_87),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_68),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

OAI221xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_72),
.B1(n_59),
.B2(n_87),
.C(n_37),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_77),
.B(n_28),
.C(n_23),
.Y(n_154)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_134),
.Y(n_163)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_136),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_109),
.B1(n_100),
.B2(n_104),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_144),
.B1(n_150),
.B2(n_152),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_100),
.A3(n_103),
.B1(n_106),
.B2(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_131),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_102),
.B1(n_111),
.B2(n_57),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_116),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_139),
.B(n_135),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_114),
.B1(n_127),
.B2(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_57),
.B1(n_75),
.B2(n_50),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_75),
.B1(n_72),
.B2(n_93),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_154),
.A2(n_134),
.B(n_96),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_49),
.B1(n_93),
.B2(n_40),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_86),
.B1(n_73),
.B2(n_62),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_105),
.B1(n_86),
.B2(n_94),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_62),
.B1(n_89),
.B2(n_43),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_170),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_185),
.B(n_190),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_189),
.B(n_141),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_176),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_118),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_186),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_129),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_77),
.B(n_96),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_46),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_105),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_151),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_165),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_198),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_147),
.C(n_150),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_206),
.C(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_165),
.B1(n_162),
.B2(n_154),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_213),
.B1(n_39),
.B2(n_36),
.Y(n_237)
);

XOR2x2_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_153),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_204),
.B(n_208),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_185),
.B(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_156),
.C(n_154),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_154),
.B(n_20),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_7),
.B(n_13),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_9),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_171),
.C(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_39),
.C(n_36),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_88),
.C(n_39),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_138),
.B1(n_137),
.B2(n_136),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_176),
.A2(n_15),
.B(n_30),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_180),
.B1(n_19),
.B2(n_21),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_15),
.B(n_30),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_190),
.B1(n_19),
.B2(n_21),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_24),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_215),
.B1(n_213),
.B2(n_202),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_209),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_207),
.B(n_206),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_21),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_113),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_24),
.C(n_36),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_212),
.B1(n_197),
.B2(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_198),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_7),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_250),
.B1(n_222),
.B2(n_227),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_201),
.B1(n_208),
.B2(n_193),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_255),
.C(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_223),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_24),
.C(n_28),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_263),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_218),
.B1(n_233),
.B2(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_221),
.B1(n_236),
.B2(n_2),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_271),
.B(n_238),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_8),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_0),
.C(n_1),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_244),
.C(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_28),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_279),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_255),
.C(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_265),
.C(n_259),
.Y(n_287)
);

BUFx12_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_278),
.B(n_285),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_11),
.B(n_1),
.Y(n_295)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

OAI31xp33_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_250),
.A3(n_249),
.B(n_8),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_5),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_275),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_272),
.C(n_1),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_294),
.B(n_281),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_292),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_5),
.B(n_10),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_0),
.B(n_2),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

AO221x1_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.C(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_11),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_2),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_301),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_306),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_3),
.C(n_4),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_289),
.B(n_298),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_310),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_287),
.B(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_304),
.B(n_277),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_291),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_314),
.B(n_315),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_309),
.B(n_307),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_274),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_278),
.C(n_279),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_302),
.B(n_3),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_4),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_4),
.C(n_229),
.Y(n_324)
);


endmodule