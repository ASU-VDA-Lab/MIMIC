module fake_jpeg_14396_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_40),
.B(n_42),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_61),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_22),
.B(n_4),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_64),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_62),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_71),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_12),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_6),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_12),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_17),
.B(n_6),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_7),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_75),
.A2(n_81),
.B1(n_97),
.B2(n_87),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_20),
.B1(n_34),
.B2(n_31),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_76),
.A2(n_95),
.B1(n_103),
.B2(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_77),
.B(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_108),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_93),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_19),
.C(n_25),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_47),
.C(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_19),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_32),
.B1(n_34),
.B2(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_35),
.B1(n_25),
.B2(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_7),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_27),
.B1(n_17),
.B2(n_52),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_27),
.B1(n_21),
.B2(n_9),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_21),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_104),
.B1(n_102),
.B2(n_96),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_21),
.B1(n_54),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_98),
.B1(n_87),
.B2(n_91),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_115),
.B(n_148),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_10),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_126),
.C(n_134),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

OR2x4_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_136),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_117),
.Y(n_175)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_135),
.B(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_137),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_82),
.C(n_98),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_94),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_143),
.Y(n_171)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_74),
.B(n_83),
.C(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_145),
.Y(n_155)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_92),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_92),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_149),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_99),
.Y(n_149)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_88),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_118),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_146),
.B1(n_119),
.B2(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_174),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_124),
.B(n_116),
.C(n_141),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_154),
.B(n_175),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_127),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_139),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_148),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_126),
.B1(n_134),
.B2(n_125),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_144),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_123),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_196),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_155),
.B(n_160),
.Y(n_201)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_153),
.B(n_123),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_192),
.C(n_198),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_194),
.B(n_165),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_142),
.C(n_150),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_155),
.A2(n_122),
.B1(n_170),
.B2(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_159),
.B1(n_168),
.B2(n_173),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_156),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_164),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_176),
.C(n_160),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_202),
.B(n_194),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_152),
.B(n_165),
.C(n_168),
.D(n_172),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_198),
.C(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_219),
.C(n_223),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_193),
.B1(n_181),
.B2(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_220),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_209),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_203),
.C(n_179),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_197),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_226),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_179),
.C(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_206),
.B(n_188),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_233),
.C(n_221),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_209),
.A3(n_205),
.B1(n_202),
.B2(n_214),
.C1(n_184),
.C2(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_229),
.B(n_232),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_182),
.B(n_205),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_202),
.B(n_182),
.Y(n_234)
);

AOI31xp67_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_207),
.A3(n_208),
.B(n_204),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_219),
.B1(n_223),
.B2(n_216),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_235),
.A2(n_173),
.B1(n_177),
.B2(n_183),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_231),
.A2(n_214),
.B1(n_189),
.B2(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.C(n_230),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_211),
.C(n_208),
.Y(n_238)
);

AOI31xp33_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_227),
.A3(n_183),
.B(n_177),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_204),
.B1(n_195),
.B2(n_207),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_232),
.B(n_233),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_245),
.B(n_246),
.C(n_244),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_246),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_235),
.Y(n_251)
);

NAND2x1p5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_237),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_249),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_249),
.B(n_178),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_167),
.Y(n_255)
);


endmodule