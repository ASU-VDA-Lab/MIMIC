module fake_aes_1987_n_19 (n_1, n_2, n_0, n_19);
input n_1;
input n_2;
input n_0;
output n_19;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_4;
wire n_7;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_0), .B(n_2), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
OAI21xp5_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_4), .B(n_0), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_3), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_7), .Y(n_12) );
AND3x1_ASAP7_75t_L g13 ( .A(n_12), .B(n_9), .C(n_3), .Y(n_13) );
NAND4xp25_ASAP7_75t_SL g14 ( .A(n_11), .B(n_6), .C(n_1), .D(n_2), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_14), .B(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_1), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_2), .B1(n_1), .B2(n_0), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_15), .B(n_18), .Y(n_19) );
endmodule