module real_jpeg_10454_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_32),
.B1(n_36),
.B2(n_42),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_9),
.B(n_55),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_5),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_21),
.B1(n_25),
.B2(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_9),
.B(n_21),
.Y(n_182)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_8),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_11),
.B1(n_43),
.B2(n_69),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_8),
.A2(n_21),
.B1(n_25),
.B2(n_43),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_36),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_11),
.B1(n_45),
.B2(n_69),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_21),
.B1(n_25),
.B2(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_93),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_9),
.B(n_50),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_52),
.B(n_56),
.C(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_24),
.B1(n_36),
.B2(n_42),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_11),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_11),
.B(n_64),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_11),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_11),
.A2(n_45),
.B(n_64),
.C(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_122),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_120),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_99),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_72),
.C(n_81),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_16),
.A2(n_17),
.B1(n_72),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_46),
.B1(n_47),
.B2(n_71),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_33),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_19),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_19),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_25),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_26),
.B(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_28),
.B1(n_87),
.B2(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_28),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_28),
.B(n_45),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_29),
.A2(n_86),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_33),
.A2(n_34),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_33),
.A2(n_34),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_34),
.B(n_136),
.C(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_34),
.B(n_214),
.C(n_220),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_44),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_35),
.A2(n_39),
.B1(n_77),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_35),
.B(n_39),
.Y(n_151)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_36),
.A2(n_45),
.B(n_53),
.Y(n_207)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_39),
.B(n_45),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_40),
.A2(n_42),
.B(n_45),
.C(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_44),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_48),
.A2(n_49),
.B1(n_149),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_48),
.A2(n_49),
.B1(n_88),
.B2(n_89),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_49),
.B(n_61),
.C(n_71),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_49),
.B(n_92),
.C(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_49),
.B(n_89),
.C(n_209),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_57),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_54),
.B1(n_98),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_52),
.B(n_56),
.C(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_56),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_59),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_104),
.C(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_61),
.A2(n_62),
.B1(n_103),
.B2(n_104),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_63),
.B(n_66),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_72),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_74),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_75),
.B(n_87),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_92),
.C(n_95),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_83),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_88),
.A2(n_89),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_89),
.B(n_181),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_127),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_118),
.B2(n_119),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_109),
.B1(n_116),
.B2(n_117),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_108),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_106),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_103),
.A2(n_104),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_168),
.C(n_169),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_141),
.B(n_230),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_124),
.B(n_138),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_130),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_128),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_131),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_189),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_136),
.A2(n_165),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_172),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_157),
.B(n_171),
.Y(n_143)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_154),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.CI(n_152),
.CON(n_145),
.SN(n_145)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_159),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_164),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_169),
.B1(n_185),
.B2(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_179),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_228),
.C(n_229),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_222),
.B(n_227),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_211),
.B(n_221),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_200),
.B(n_210),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_192),
.B(n_199),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_191),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_188),
.B(n_190),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_213),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);


endmodule