module fake_netlist_1_6370_n_741 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_741);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_741;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_76), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_36), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_63), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_44), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
BUFx2_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_80), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_52), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_47), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_5), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_55), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_21), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_10), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_4), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_27), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_77), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_70), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_9), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_3), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_40), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_37), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_20), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_13), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_49), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_59), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_10), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_51), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_22), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_62), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_48), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_46), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_30), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_43), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_6), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_24), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_2), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_130), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_130), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_95), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_134) );
CKINVDCx8_ASAP7_75t_R g135 ( .A(n_116), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_109), .B(n_0), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_130), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_89), .B(n_1), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_89), .B(n_4), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_113), .B(n_129), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_111), .B(n_5), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
NAND2xp33_ASAP7_75t_L g149 ( .A(n_117), .B(n_79), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_81), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_129), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_111), .B(n_7), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_93), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_156) );
NOR2x1_ASAP7_75t_L g157 ( .A(n_87), .B(n_11), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_83), .Y(n_160) );
INVxp33_ASAP7_75t_SL g161 ( .A(n_107), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_93), .B(n_11), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_83), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_128), .B(n_13), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
NAND2xp33_ASAP7_75t_SL g166 ( .A(n_112), .B(n_14), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_90), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_121), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_116), .B(n_14), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_119), .Y(n_171) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_91), .A2(n_42), .B(n_73), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_91), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_121), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_167), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_140), .B(n_125), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_143), .B(n_125), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_144), .B(n_102), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_161), .B(n_84), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_143), .A2(n_96), .B1(n_108), .B2(n_103), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_135), .B(n_94), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_140), .B(n_97), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_146), .B(n_97), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_170), .B(n_106), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_154), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_135), .A2(n_106), .B1(n_101), .B2(n_102), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
OAI22xp33_ASAP7_75t_SL g207 ( .A1(n_142), .A2(n_101), .B1(n_126), .B2(n_105), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
INVxp33_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_146), .B(n_85), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_150), .B(n_114), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_162), .B(n_127), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_160), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_160), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_136), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
CKINVDCx8_ASAP7_75t_R g221 ( .A(n_138), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_160), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_150), .B(n_124), .Y(n_223) );
BUFx4f_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_154), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_163), .Y(n_228) );
AND2x6_ASAP7_75t_L g229 ( .A(n_157), .B(n_127), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_164), .B(n_158), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_163), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_159), .B(n_126), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_159), .B(n_110), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_136), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_131), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_142), .A2(n_110), .B1(n_123), .B2(n_98), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_156), .B(n_92), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_163), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_131), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_165), .B(n_122), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_131), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
INVx5_ASAP7_75t_L g244 ( .A(n_180), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_214), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_176), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_178), .B(n_165), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_175), .B(n_145), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_229), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_189), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_179), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_230), .B(n_145), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_224), .B(n_168), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_183), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_179), .A2(n_155), .B1(n_166), .B2(n_149), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_230), .B(n_173), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_180), .Y(n_258) );
NAND3xp33_ASAP7_75t_SL g259 ( .A(n_238), .B(n_171), .C(n_156), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_214), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_234), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_210), .B(n_173), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_180), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_183), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_187), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_214), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_177), .A2(n_172), .B(n_168), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_224), .B(n_212), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_180), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_183), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_224), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_185), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_209), .B(n_155), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_185), .Y(n_277) );
BUFx12f_ASAP7_75t_SL g278 ( .A(n_197), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_199), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_185), .Y(n_280) );
AND2x6_ASAP7_75t_SL g281 ( .A(n_191), .B(n_197), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_215), .B(n_157), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_190), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_212), .B(n_172), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_185), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_212), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_221), .B(n_153), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_193), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_241), .B(n_153), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_193), .B(n_153), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_193), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_229), .A2(n_174), .B1(n_169), .B2(n_153), .Y(n_294) );
OAI22xp5_ASAP7_75t_SL g295 ( .A1(n_190), .A2(n_134), .B1(n_172), .B2(n_98), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_193), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_196), .B(n_174), .Y(n_297) );
BUFx8_ASAP7_75t_L g298 ( .A(n_229), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_196), .B(n_174), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_236), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_196), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_212), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_229), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_196), .B(n_169), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_204), .A2(n_134), .B1(n_82), .B2(n_169), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_221), .B(n_115), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_207), .A2(n_118), .B(n_100), .C(n_104), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_240), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_177), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_232), .B(n_120), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_181), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_228), .B(n_15), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_181), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_232), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_314), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_261), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_253), .B(n_232), .Y(n_318) );
BUFx12f_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_245), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_249), .A2(n_252), .B1(n_266), .B2(n_253), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_253), .B(n_232), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_244), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_245), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_278), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_276), .B(n_207), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_252), .A2(n_229), .B1(n_233), .B2(n_237), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_260), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_282), .B(n_233), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_280), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_264), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_260), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_223), .B(n_228), .C(n_239), .Y(n_340) );
INVx6_ASAP7_75t_L g341 ( .A(n_244), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_267), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_248), .A2(n_231), .B(n_239), .C(n_233), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_262), .A2(n_200), .B(n_198), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_244), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_251), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_268), .A2(n_198), .B(n_203), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_282), .B(n_233), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_283), .A2(n_229), .B1(n_231), .B2(n_205), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_264), .Y(n_353) );
INVx5_ASAP7_75t_L g354 ( .A(n_244), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_254), .A2(n_205), .B(n_200), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_276), .B(n_202), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_288), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_295), .A2(n_229), .B1(n_202), .B2(n_203), .Y(n_358) );
BUFx2_ASAP7_75t_R g359 ( .A(n_266), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_286), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_302), .A2(n_186), .B1(n_195), .B2(n_99), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_267), .Y(n_362) );
AOI21x1_ASAP7_75t_L g363 ( .A1(n_254), .A2(n_216), .B(n_217), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_302), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g365 ( .A1(n_259), .A2(n_115), .B(n_99), .C(n_123), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_250), .B(n_186), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_244), .B(n_100), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_296), .B(n_186), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_256), .B(n_186), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_289), .B(n_104), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_322), .A2(n_305), .B(n_307), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_365), .B(n_257), .C(n_291), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_324), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_316), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_325), .B(n_315), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_347), .B(n_283), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_320), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_317), .A2(n_290), .B1(n_303), .B2(n_250), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_332), .A2(n_290), .B1(n_303), .B2(n_298), .Y(n_380) );
AOI21x1_ASAP7_75t_L g381 ( .A1(n_363), .A2(n_208), .B(n_213), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_328), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_325), .A2(n_298), .B1(n_255), .B2(n_274), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_350), .A2(n_313), .B(n_120), .Y(n_384) );
CKINVDCx11_ASAP7_75t_R g385 ( .A(n_319), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_317), .B(n_281), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_325), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_354), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_360), .B(n_270), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_316), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_320), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_327), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_356), .B(n_304), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_358), .A2(n_297), .B1(n_299), .B2(n_310), .Y(n_394) );
AOI21xp5_ASAP7_75t_SL g395 ( .A1(n_316), .A2(n_172), .B(n_297), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g396 ( .A1(n_340), .A2(n_285), .B(n_312), .Y(n_396) );
OR2x6_ASAP7_75t_L g397 ( .A(n_316), .B(n_270), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_335), .B(n_304), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_335), .A2(n_298), .B1(n_274), .B2(n_255), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_329), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_330), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_344), .A2(n_285), .B(n_311), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_336), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_339), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_393), .B(n_335), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_377), .A2(n_319), .B1(n_331), .B2(n_323), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_372), .A2(n_333), .B1(n_352), .B2(n_351), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_372), .A2(n_371), .B(n_370), .C(n_323), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_373), .A2(n_351), .B1(n_348), .B2(n_367), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_402), .A2(n_340), .B(n_343), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_393), .A2(n_343), .B1(n_357), .B2(n_364), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_394), .A2(n_331), .B1(n_348), .B2(n_367), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_373), .A2(n_351), .B1(n_318), .B2(n_292), .C(n_311), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_394), .A2(n_367), .B1(n_297), .B2(n_243), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_387), .A2(n_316), .B1(n_368), .B2(n_359), .Y(n_416) );
NOR2x1_ASAP7_75t_SL g417 ( .A(n_388), .B(n_354), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_388), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_386), .A2(n_273), .B1(n_326), .B2(n_346), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_368), .B1(n_250), .B2(n_361), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_398), .A2(n_247), .B1(n_246), .B2(n_349), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_398), .B(n_345), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_374), .B(n_258), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_374), .B(n_354), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_375), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_378), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_382), .B(n_354), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_400), .B1(n_404), .B2(n_403), .C(n_382), .Y(n_428) );
OR2x6_ASAP7_75t_L g429 ( .A(n_388), .B(n_368), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_384), .A2(n_368), .B1(n_354), .B2(n_341), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_380), .A2(n_321), .B1(n_337), .B2(n_353), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_396), .A2(n_368), .B1(n_334), .B2(n_362), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_396), .A2(n_334), .B1(n_338), .B2(n_362), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_433), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_426), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_408), .B(n_405), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_415), .A2(n_405), .B1(n_392), .B2(n_378), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_428), .B(n_378), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_413), .A2(n_399), .B1(n_383), .B2(n_401), .C(n_404), .Y(n_441) );
AOI33xp33_ASAP7_75t_L g442 ( .A1(n_407), .A2(n_410), .A3(n_105), .B1(n_114), .B2(n_118), .B3(n_415), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_409), .A2(n_379), .B1(n_401), .B2(n_403), .Y(n_443) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_412), .A2(n_124), .A3(n_216), .B1(n_217), .B2(n_218), .B3(n_220), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_414), .A2(n_397), .B1(n_376), .B2(n_402), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_429), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_418), .B(n_391), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_391), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_425), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_416), .A2(n_397), .B1(n_376), .B2(n_385), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_430), .A2(n_384), .B1(n_397), .B2(n_392), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_421), .A2(n_397), .B1(n_384), .B2(n_337), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_422), .B(n_326), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_421), .A2(n_294), .B1(n_395), .B2(n_355), .C(n_369), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_419), .B(n_395), .C(n_147), .D(n_148), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_427), .A2(n_392), .B1(n_391), .B2(n_265), .C(n_272), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_417), .B(n_390), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_434), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_431), .A2(n_397), .B1(n_384), .B2(n_321), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_429), .B(n_346), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
OAI211xp5_ASAP7_75t_L g466 ( .A1(n_432), .A2(n_384), .B(n_366), .C(n_337), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_425), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_425), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_432), .B(n_390), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_420), .B(n_390), .Y(n_471) );
OR2x2_ASAP7_75t_SL g472 ( .A(n_424), .B(n_375), .Y(n_472) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_466), .A2(n_381), .B(n_366), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_447), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_435), .B(n_16), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_440), .B(n_375), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_436), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_443), .B(n_136), .C(n_141), .Y(n_479) );
AOI211xp5_ASAP7_75t_SL g480 ( .A1(n_441), .A2(n_390), .B(n_353), .C(n_321), .Y(n_480) );
OAI221xp5_ASAP7_75t_SL g481 ( .A1(n_442), .A2(n_147), .B1(n_148), .B2(n_353), .C(n_338), .Y(n_481) );
OAI211xp5_ASAP7_75t_SL g482 ( .A1(n_441), .A2(n_147), .B(n_148), .C(n_225), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_461), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_451), .B(n_375), .Y(n_484) );
NAND4xp25_ASAP7_75t_SL g485 ( .A(n_450), .B(n_16), .C(n_17), .D(n_18), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_448), .B(n_17), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_472), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_472), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_438), .A2(n_273), .B1(n_341), .B2(n_342), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g491 ( .A1(n_438), .A2(n_18), .B1(n_19), .B2(n_20), .C1(n_21), .C2(n_195), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g492 ( .A1(n_452), .A2(n_375), .B1(n_341), .B2(n_19), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_455), .B(n_375), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_443), .A2(n_381), .B(n_342), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_454), .A2(n_341), .B1(n_265), .B2(n_272), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_445), .A2(n_195), .B1(n_218), .B2(n_220), .C(n_222), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_451), .B(n_141), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_453), .B(n_151), .C(n_141), .Y(n_498) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_439), .A2(n_184), .B(n_192), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
AND4x1_ASAP7_75t_L g501 ( .A(n_464), .B(n_222), .C(n_225), .D(n_31), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_462), .B(n_141), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_462), .B(n_141), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_440), .B(n_195), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_470), .B(n_26), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_465), .B(n_141), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_457), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_457), .B(n_271), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_458), .A2(n_269), .B1(n_213), .B2(n_208), .C(n_184), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_437), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_465), .A2(n_151), .B1(n_226), .B2(n_201), .C(n_192), .Y(n_512) );
AND2x4_ASAP7_75t_SL g513 ( .A(n_461), .B(n_284), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_447), .Y(n_514) );
NAND2xp33_ASAP7_75t_R g515 ( .A(n_452), .B(n_28), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_460), .B(n_271), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_458), .B(n_151), .C(n_188), .Y(n_518) );
AOI211xp5_ASAP7_75t_SL g519 ( .A1(n_439), .A2(n_227), .B(n_194), .C(n_201), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_151), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_446), .B(n_151), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_446), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_463), .A2(n_279), .B(n_194), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_446), .B(n_151), .Y(n_524) );
INVxp33_ASAP7_75t_SL g525 ( .A(n_467), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_471), .B(n_227), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_500), .B(n_467), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_526), .B(n_471), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_478), .Y(n_529) );
NAND4xp25_ASAP7_75t_SL g530 ( .A(n_491), .B(n_456), .C(n_459), .D(n_467), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_485), .B(n_444), .C(n_456), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_526), .B(n_468), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_505), .B(n_469), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
NAND2xp33_ASAP7_75t_L g535 ( .A(n_492), .B(n_468), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_487), .B(n_469), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_476), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_520), .B(n_468), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_520), .B(n_469), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_490), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_508), .B(n_449), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_480), .B(n_188), .C(n_226), .D(n_449), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_516), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_493), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_511), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_511), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_497), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_484), .B(n_437), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_514), .B(n_449), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_484), .B(n_437), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_513), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_515), .B(n_182), .C(n_206), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_475), .B(n_242), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_487), .B(n_242), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_488), .B(n_240), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_518), .A2(n_269), .B(n_271), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_513), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_497), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_502), .B(n_32), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_477), .A2(n_271), .B1(n_263), .B2(n_284), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_486), .Y(n_561) );
NAND3x1_ASAP7_75t_L g562 ( .A(n_515), .B(n_33), .C(n_34), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_502), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_503), .B(n_35), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_474), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_481), .B(n_182), .C(n_206), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_488), .B(n_39), .Y(n_567) );
NAND4xp75_ASAP7_75t_L g568 ( .A(n_483), .B(n_41), .C(n_45), .D(n_50), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_503), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_507), .B(n_53), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_507), .B(n_56), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_483), .B(n_58), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_504), .B(n_60), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_477), .B(n_61), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_525), .B(n_271), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_522), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_506), .B(n_64), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_499), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_525), .B(n_65), .Y(n_579) );
NOR2x1p5_ASAP7_75t_L g580 ( .A(n_506), .B(n_66), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_489), .B(n_67), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_506), .B(n_68), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_499), .Y(n_583) );
AOI31xp33_ASAP7_75t_L g584 ( .A1(n_519), .A2(n_72), .A3(n_74), .B(n_309), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_521), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_524), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_494), .B(n_279), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_509), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_473), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_544), .B(n_473), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_565), .B(n_517), .Y(n_591) );
INVx4_ASAP7_75t_L g592 ( .A(n_551), .Y(n_592) );
NAND2x1_ASAP7_75t_SL g593 ( .A(n_577), .B(n_495), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_537), .Y(n_594) );
NOR2x1p5_ASAP7_75t_L g595 ( .A(n_552), .B(n_479), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_528), .B(n_523), .Y(n_596) );
OAI32xp33_ASAP7_75t_L g597 ( .A1(n_552), .A2(n_498), .A3(n_482), .B1(n_501), .B2(n_496), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_537), .Y(n_598) );
XOR2x2_ASAP7_75t_L g599 ( .A(n_562), .B(n_510), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_528), .B(n_512), .Y(n_600) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_535), .B(n_182), .C(n_206), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_585), .B(n_309), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_557), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_585), .B(n_306), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_586), .B(n_306), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_540), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_544), .B(n_182), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_540), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_567), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_551), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_543), .B(n_182), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_543), .B(n_206), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_580), .A2(n_300), .B1(n_263), .B2(n_284), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_530), .B(n_300), .C(n_211), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_534), .B(n_206), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_576), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_531), .A2(n_263), .B1(n_284), .B2(n_235), .Y(n_618) );
OAI31xp33_ASAP7_75t_L g619 ( .A1(n_580), .A2(n_211), .A3(n_219), .B(n_235), .Y(n_619) );
NAND2x1p5_ASAP7_75t_SL g620 ( .A(n_577), .B(n_211), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_575), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_576), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_534), .Y(n_623) );
NAND2x1_ASAP7_75t_SL g624 ( .A(n_574), .B(n_211), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_572), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_541), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_533), .Y(n_627) );
AOI21xp33_ASAP7_75t_SL g628 ( .A1(n_584), .A2(n_211), .B(n_219), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_561), .B(n_219), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_536), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_567), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_532), .B(n_219), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_527), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_586), .B(n_219), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_588), .B(n_235), .C(n_284), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_569), .B(n_235), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_536), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_569), .B(n_235), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_554), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_554), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_579), .B(n_263), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_563), .B(n_263), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_594), .Y(n_644) );
XNOR2x1_ASAP7_75t_L g645 ( .A(n_599), .B(n_582), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_626), .B(n_633), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_598), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_627), .B(n_546), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_609), .Y(n_650) );
XOR2x2_ASAP7_75t_L g651 ( .A(n_603), .B(n_562), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_617), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_622), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_630), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_638), .B(n_563), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_611), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_634), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_596), .B(n_532), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_592), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_591), .B(n_547), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_615), .B(n_582), .C(n_574), .D(n_542), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_640), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_608), .B(n_641), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_592), .Y(n_665) );
AOI21xp33_ASAP7_75t_SL g666 ( .A1(n_620), .A2(n_566), .B(n_572), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_612), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_610), .A2(n_558), .B1(n_547), .B2(n_553), .C(n_578), .Y(n_668) );
XNOR2x2_ASAP7_75t_L g669 ( .A(n_601), .B(n_566), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_612), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_629), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_613), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_613), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_590), .B(n_545), .Y(n_674) );
XOR2x2_ASAP7_75t_L g675 ( .A(n_593), .B(n_568), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_590), .B(n_545), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_635), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_614), .A2(n_578), .B(n_570), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_631), .B(n_546), .Y(n_679) );
AOI211x1_ASAP7_75t_L g680 ( .A1(n_597), .A2(n_581), .B(n_573), .C(n_564), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_600), .A2(n_558), .B1(n_589), .B2(n_548), .C(n_550), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_607), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g684 ( .A(n_625), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_621), .A2(n_560), .B1(n_568), .B2(n_555), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_607), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_602), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_604), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_605), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_628), .A2(n_555), .B(n_559), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_614), .B(n_564), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_619), .B(n_583), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_632), .B(n_548), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_637), .B(n_550), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_636), .B(n_570), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_637), .B(n_538), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_595), .A2(n_538), .B1(n_539), .B2(n_571), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_642), .A2(n_583), .B(n_559), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_639), .A2(n_571), .B(n_589), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_639), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_643), .B(n_539), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_618), .A2(n_556), .B1(n_587), .B2(n_643), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_624), .A2(n_587), .B(n_616), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_616), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_645), .A2(n_660), .B1(n_665), .B2(n_684), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_646), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_662), .B(n_690), .Y(n_707) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_685), .B(n_692), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_646), .Y(n_709) );
INVxp67_ASAP7_75t_L g710 ( .A(n_651), .Y(n_710) );
NOR2x1_ASAP7_75t_L g711 ( .A(n_692), .B(n_695), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_680), .A2(n_657), .B1(n_681), .B2(n_663), .C(n_668), .Y(n_712) );
AOI31xp33_ASAP7_75t_L g713 ( .A1(n_656), .A2(n_666), .A3(n_695), .B(n_691), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g714 ( .A1(n_675), .A2(n_678), .B(n_691), .Y(n_714) );
OA22x2_ASAP7_75t_L g715 ( .A1(n_697), .A2(n_654), .B1(n_659), .B2(n_687), .Y(n_715) );
AOI322xp5_ASAP7_75t_L g716 ( .A1(n_668), .A2(n_688), .A3(n_689), .B1(n_648), .B2(n_650), .C1(n_652), .C2(n_653), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_698), .B(n_703), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_661), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_706), .Y(n_719) );
NAND4xp75_ASAP7_75t_L g720 ( .A(n_708), .B(n_702), .C(n_677), .D(n_682), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_712), .B(n_671), .Y(n_721) );
OAI211xp5_ASAP7_75t_SL g722 ( .A1(n_710), .A2(n_699), .B(n_679), .C(n_664), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_713), .A2(n_649), .B(n_679), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_707), .A2(n_696), .B1(n_647), .B2(n_644), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_714), .A2(n_700), .B1(n_658), .B2(n_673), .Y(n_725) );
NOR2xp67_ASAP7_75t_L g726 ( .A(n_717), .B(n_674), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_719), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_720), .B(n_705), .C(n_711), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_721), .A2(n_709), .B1(n_718), .B2(n_664), .C(n_672), .Y(n_729) );
NOR3xp33_ASAP7_75t_SL g730 ( .A(n_722), .B(n_715), .C(n_716), .Y(n_730) );
XNOR2x1_ASAP7_75t_L g731 ( .A(n_725), .B(n_669), .Y(n_731) );
OAI211xp5_ASAP7_75t_SL g732 ( .A1(n_728), .A2(n_724), .B(n_716), .C(n_723), .Y(n_732) );
AND3x1_ASAP7_75t_L g733 ( .A(n_730), .B(n_726), .C(n_649), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_731), .A2(n_667), .B1(n_670), .B2(n_683), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_733), .A2(n_729), .B1(n_727), .B2(n_686), .C(n_676), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_732), .A2(n_704), .B1(n_694), .B2(n_701), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_736), .B(n_734), .C(n_674), .Y(n_737) );
AND2x2_ASAP7_75t_SL g738 ( .A(n_735), .B(n_655), .Y(n_738) );
INVx4_ASAP7_75t_L g739 ( .A(n_738), .Y(n_739) );
XNOR2xp5_ASAP7_75t_L g740 ( .A(n_739), .B(n_737), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_740), .A2(n_693), .B1(n_704), .B2(n_676), .Y(n_741) );
endmodule