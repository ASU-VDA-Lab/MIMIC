module fake_netlist_1_2134_n_1306 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1306);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1306;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_92), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_21), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_200), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_14), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_109), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_269), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_194), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_279), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_187), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_215), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_85), .Y(n_291) );
INVxp33_ASAP7_75t_SL g292 ( .A(n_253), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_142), .Y(n_293) );
CKINVDCx16_ASAP7_75t_R g294 ( .A(n_171), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_33), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_129), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_245), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_226), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_143), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_162), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_34), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_155), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_178), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_151), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_248), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_127), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_73), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_251), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_102), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_136), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_227), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_53), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_177), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_6), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_125), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_184), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_72), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_131), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_205), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_130), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_98), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_261), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_272), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_280), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_153), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_15), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_260), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_164), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_74), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_62), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_93), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_38), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_192), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_26), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_148), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_8), .Y(n_339) );
INVxp33_ASAP7_75t_SL g340 ( .A(n_23), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_48), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_161), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_240), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_9), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_146), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_50), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_41), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_198), .Y(n_348) );
CKINVDCx14_ASAP7_75t_R g349 ( .A(n_232), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_81), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_176), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_225), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_111), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_144), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_69), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_54), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_134), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_159), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_264), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_149), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_52), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_33), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_80), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_1), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_145), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_190), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_209), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_189), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_113), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_4), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_141), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_124), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_18), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_40), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_100), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_84), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_197), .Y(n_377) );
INVxp33_ASAP7_75t_L g378 ( .A(n_277), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_163), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_22), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_246), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_15), .Y(n_382) );
INVxp33_ASAP7_75t_SL g383 ( .A(n_167), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_28), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_50), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_135), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_185), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_230), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_28), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_29), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_57), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_181), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_250), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_7), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_249), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_274), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_0), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_154), .Y(n_398) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_75), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_13), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_271), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_101), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_29), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_174), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_235), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_31), .B(n_70), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_115), .Y(n_407) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_114), .B(n_96), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_49), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_9), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_139), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_262), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_199), .Y(n_413) );
BUFx10_ASAP7_75t_L g414 ( .A(n_255), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_132), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_270), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_175), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_51), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_244), .Y(n_419) );
NAND2xp33_ASAP7_75t_L g420 ( .A(n_378), .B(n_66), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_288), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_284), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_288), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_284), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_313), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_375), .B(n_0), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_313), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_288), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_378), .B(n_1), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_297), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_283), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_288), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_289), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_286), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_294), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_349), .B(n_2), .Y(n_436) );
OAI22xp5_ASAP7_75t_SL g437 ( .A1(n_340), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g438 ( .A1(n_340), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_402), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_290), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_414), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_325), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_291), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_293), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_285), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_300), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_314), .Y(n_447) );
BUFx10_ASAP7_75t_L g448 ( .A(n_371), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_371), .B(n_5), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_325), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_325), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_349), .B(n_7), .Y(n_452) );
BUFx10_ASAP7_75t_L g453 ( .A(n_434), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_441), .B(n_309), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_430), .B(n_384), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_430), .B(n_384), .Y(n_459) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_445), .B(n_285), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
AND2x6_ASAP7_75t_L g465 ( .A(n_436), .B(n_314), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_441), .B(n_414), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_423), .Y(n_468) );
AND2x6_ASAP7_75t_L g469 ( .A(n_436), .B(n_411), .Y(n_469) );
INVx6_ASAP7_75t_L g470 ( .A(n_448), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_432), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_441), .Y(n_474) );
INVx8_ASAP7_75t_L g475 ( .A(n_441), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_441), .B(n_414), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_452), .A2(n_282), .B1(n_315), .B2(n_302), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_447), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_450), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_450), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_450), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_451), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_451), .Y(n_484) );
INVx6_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_448), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_452), .A2(n_333), .B1(n_335), .B2(n_329), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_431), .B(n_385), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_448), .Y(n_490) );
AND2x6_ASAP7_75t_L g491 ( .A(n_452), .B(n_411), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_451), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_431), .B(n_385), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_422), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_426), .B(n_356), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_424), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_454), .B(n_467), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_454), .B(n_426), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_458), .B(n_433), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_498), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_496), .B(n_433), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_498), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_475), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_453), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_459), .B(n_440), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_465), .A2(n_443), .B1(n_444), .B2(n_440), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_475), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_489), .B(n_443), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_496), .B(n_444), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_486), .B(n_446), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_486), .B(n_446), .Y(n_513) );
AO22x1_ASAP7_75t_L g514 ( .A1(n_465), .A2(n_439), .B1(n_435), .B2(n_292), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_492), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_494), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_495), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_486), .B(n_449), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_486), .B(n_449), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_487), .B(n_447), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_492), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_474), .A2(n_420), .B(n_413), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_492), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_465), .A2(n_429), .B1(n_383), .B2(n_292), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_492), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_462), .Y(n_527) );
AND3x2_ASAP7_75t_SL g528 ( .A(n_460), .B(n_438), .C(n_437), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_476), .B(n_429), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_487), .B(n_281), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_475), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_453), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_495), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_497), .A2(n_425), .B(n_427), .C(n_424), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_453), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_487), .B(n_301), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_487), .B(n_281), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_474), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_465), .A2(n_383), .B1(n_399), .B2(n_341), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_456), .B(n_342), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_465), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_475), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_475), .A2(n_413), .B(n_305), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_477), .A2(n_311), .B1(n_327), .B2(n_287), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_465), .Y(n_547) );
INVx4_ASAP7_75t_L g548 ( .A(n_470), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_490), .B(n_298), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_469), .A2(n_438), .B1(n_437), .B2(n_311), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_490), .B(n_304), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_469), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_469), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_490), .B(n_306), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_490), .B(n_298), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_466), .Y(n_556) );
NOR2x1p5_ASAP7_75t_L g557 ( .A(n_460), .B(n_397), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_469), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_478), .B(n_308), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_478), .B(n_337), .Y(n_560) );
NOR2x1p5_ASAP7_75t_L g561 ( .A(n_453), .B(n_397), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_488), .A2(n_364), .B(n_382), .C(n_339), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_469), .A2(n_399), .B1(n_347), .B2(n_361), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_457), .A2(n_463), .B(n_461), .Y(n_564) );
BUFx12f_ASAP7_75t_L g565 ( .A(n_469), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_457), .A2(n_305), .B(n_295), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_470), .B(n_299), .Y(n_567) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_469), .B(n_418), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_461), .B(n_310), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_470), .B(n_372), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_491), .B(n_400), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_470), .B(n_299), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_491), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_491), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_491), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_485), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_485), .B(n_303), .Y(n_577) );
OR2x6_ASAP7_75t_L g578 ( .A(n_485), .B(n_344), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_485), .B(n_303), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_491), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_463), .A2(n_317), .B(n_316), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_466), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_491), .A2(n_327), .B1(n_343), .B2(n_287), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_491), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_472), .A2(n_362), .B1(n_374), .B2(n_373), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_502), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_509), .B(n_307), .Y(n_587) );
INVx6_ASAP7_75t_L g588 ( .A(n_561), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_515), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_503), .B(n_409), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g591 ( .A1(n_550), .A2(n_391), .B1(n_403), .B2(n_400), .C(n_296), .Y(n_591) );
BUFx3_ASAP7_75t_L g592 ( .A(n_506), .Y(n_592) );
BUFx10_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_562), .A2(n_389), .B(n_390), .C(n_380), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_511), .B(n_403), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_516), .B(n_500), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_535), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_578), .A2(n_379), .B1(n_419), .B2(n_343), .Y(n_600) );
NOR2xp67_ASAP7_75t_SL g601 ( .A(n_505), .B(n_307), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_505), .Y(n_602) );
INVx4_ASAP7_75t_L g603 ( .A(n_578), .Y(n_603) );
INVx6_ASAP7_75t_L g604 ( .A(n_529), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_578), .A2(n_379), .B1(n_419), .B2(n_388), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_499), .B(n_346), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_532), .B(n_394), .Y(n_607) );
BUFx5_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_518), .A2(n_376), .B(n_358), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_534), .A2(n_410), .B(n_427), .C(n_425), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_501), .B(n_370), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_507), .B(n_324), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_578), .Y(n_613) );
AOI21x1_ASAP7_75t_L g614 ( .A1(n_536), .A2(n_473), .B(n_472), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_529), .B(n_324), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_529), .B(n_510), .Y(n_616) );
OA21x2_ASAP7_75t_L g617 ( .A1(n_581), .A2(n_323), .B(n_295), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_504), .A2(n_319), .B(n_322), .C(n_321), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_585), .A2(n_381), .B1(n_326), .B2(n_328), .C(n_331), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_545), .B(n_388), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_519), .A2(n_479), .B(n_473), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_499), .B(n_318), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_515), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_535), .Y(n_624) );
AO22x1_ASAP7_75t_L g625 ( .A1(n_571), .A2(n_320), .B1(n_334), .B2(n_330), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_517), .Y(n_626) );
INVx4_ASAP7_75t_L g627 ( .A(n_565), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_583), .A2(n_406), .B1(n_332), .B2(n_348), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_499), .B(n_338), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_533), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_571), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_512), .A2(n_484), .B(n_479), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_508), .B(n_367), .Y(n_633) );
CKINVDCx6p67_ASAP7_75t_R g634 ( .A(n_568), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_531), .B(n_377), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_514), .B(n_312), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_531), .A2(n_418), .B1(n_336), .B2(n_351), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_512), .A2(n_493), .B(n_484), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_568), .B(n_407), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_543), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_557), .B(n_418), .Y(n_641) );
BUFx12f_ASAP7_75t_L g642 ( .A(n_560), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_521), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_541), .B(n_416), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_575), .B(n_350), .Y(n_645) );
NAND2x1_ASAP7_75t_SL g646 ( .A(n_528), .B(n_408), .Y(n_646) );
INVx4_ASAP7_75t_L g647 ( .A(n_560), .Y(n_647) );
CKINVDCx11_ASAP7_75t_R g648 ( .A(n_528), .Y(n_648) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_543), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_539), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_573), .B(n_352), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_534), .A2(n_354), .B(n_355), .C(n_353), .Y(n_652) );
INVx4_ASAP7_75t_L g653 ( .A(n_548), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_539), .A2(n_418), .B1(n_359), .B2(n_360), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_559), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_573), .B(n_357), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_521), .Y(n_657) );
INVx3_ASAP7_75t_L g658 ( .A(n_548), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_523), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_524), .B(n_8), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_559), .A2(n_569), .B(n_536), .C(n_554), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_530), .B(n_363), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_566), .A2(n_522), .B(n_570), .C(n_538), .Y(n_663) );
OR2x6_ASAP7_75t_SL g664 ( .A(n_537), .B(n_365), .Y(n_664) );
BUFx4f_ASAP7_75t_SL g665 ( .A(n_569), .Y(n_665) );
O2A1O1Ixp5_ASAP7_75t_SL g666 ( .A1(n_551), .A2(n_368), .B(n_369), .C(n_366), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_549), .B(n_386), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_584), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_523), .Y(n_669) );
INVx5_ASAP7_75t_L g670 ( .A(n_584), .Y(n_670) );
INVx4_ASAP7_75t_L g671 ( .A(n_548), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_546), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_525), .Y(n_673) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_576), .Y(n_674) );
CKINVDCx8_ASAP7_75t_R g675 ( .A(n_540), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_525), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_555), .B(n_392), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_513), .A2(n_493), .B(n_455), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_582), .Y(n_679) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_546), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_563), .A2(n_412), .B1(n_393), .B2(n_395), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_526), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_526), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_513), .A2(n_455), .B(n_404), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_567), .B(n_398), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_572), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_582), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_542), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_547), .Y(n_689) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_577), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_527), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_579), .A2(n_417), .B1(n_415), .B2(n_323), .Y(n_692) );
BUFx2_ASAP7_75t_L g693 ( .A(n_552), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_527), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_553), .B(n_10), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_558), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_544), .A2(n_345), .B(n_401), .C(n_396), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_520), .A2(n_455), .B(n_387), .Y(n_698) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_574), .Y(n_699) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_580), .B(n_345), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_551), .B(n_10), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_564), .A2(n_405), .B(n_401), .C(n_396), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_556), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_554), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_556), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_502), .Y(n_706) );
INVx1_ASAP7_75t_SL g707 ( .A(n_503), .Y(n_707) );
BUFx12f_ASAP7_75t_L g708 ( .A(n_557), .Y(n_708) );
AO21x2_ASAP7_75t_L g709 ( .A1(n_534), .A2(n_405), .B(n_387), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_663), .A2(n_480), .B(n_471), .Y(n_710) );
BUFx3_ASAP7_75t_L g711 ( .A(n_642), .Y(n_711) );
OAI222xp33_ASAP7_75t_L g712 ( .A1(n_600), .A2(n_11), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_16), .Y(n_712) );
OAI21x1_ASAP7_75t_L g713 ( .A1(n_614), .A2(n_480), .B(n_471), .Y(n_713) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_698), .A2(n_482), .B(n_481), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_606), .A2(n_325), .B(n_11), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_624), .Y(n_716) );
OA21x2_ASAP7_75t_L g717 ( .A1(n_702), .A2(n_482), .B(n_481), .Y(n_717) );
NOR2xp33_ASAP7_75t_SL g718 ( .A(n_605), .B(n_483), .Y(n_718) );
OA21x2_ASAP7_75t_L g719 ( .A1(n_697), .A2(n_483), .B(n_442), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_594), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_616), .A2(n_468), .B(n_464), .Y(n_721) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_666), .A2(n_442), .B(n_423), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_593), .Y(n_723) );
OAI21x1_ASAP7_75t_SL g724 ( .A1(n_603), .A2(n_12), .B(n_16), .Y(n_724) );
OAI21x1_ASAP7_75t_L g725 ( .A1(n_678), .A2(n_442), .B(n_423), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_707), .B(n_17), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_664), .A2(n_423), .B1(n_442), .B2(n_19), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_598), .B(n_17), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_604), .B(n_18), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_617), .A2(n_442), .B(n_423), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_603), .Y(n_731) );
AND2x4_ASAP7_75t_L g732 ( .A(n_647), .B(n_19), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_586), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_597), .B(n_20), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_586), .Y(n_735) );
OAI21x1_ASAP7_75t_L g736 ( .A1(n_617), .A2(n_442), .B(n_464), .Y(n_736) );
NOR2x1_ASAP7_75t_SL g737 ( .A(n_613), .B(n_442), .Y(n_737) );
OAI21x1_ASAP7_75t_L g738 ( .A1(n_700), .A2(n_468), .B(n_464), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_595), .Y(n_739) );
AO32x2_ASAP7_75t_L g740 ( .A1(n_692), .A2(n_20), .A3(n_21), .B1(n_22), .B2(n_23), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_620), .B(n_24), .Y(n_741) );
OA21x2_ASAP7_75t_L g742 ( .A1(n_652), .A2(n_468), .B(n_464), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_626), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_626), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_591), .B(n_24), .C(n_25), .Y(n_745) );
INVx1_ASAP7_75t_SL g746 ( .A(n_613), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_703), .Y(n_747) );
OAI21x1_ASAP7_75t_L g748 ( .A1(n_684), .A2(n_468), .B(n_464), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_632), .A2(n_468), .B(n_464), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g750 ( .A(n_613), .B(n_25), .Y(n_750) );
OAI21x1_ASAP7_75t_L g751 ( .A1(n_638), .A2(n_468), .B(n_68), .Y(n_751) );
OA21x2_ASAP7_75t_L g752 ( .A1(n_685), .A2(n_71), .B(n_67), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_630), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_630), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_596), .A2(n_26), .B(n_27), .C(n_30), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_593), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_661), .A2(n_77), .B(n_76), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_590), .B(n_27), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_621), .A2(n_79), .B(n_78), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_590), .B(n_30), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_647), .B(n_31), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_706), .A2(n_705), .B(n_703), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_628), .A2(n_32), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_631), .B(n_32), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_706), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_660), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_604), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_701), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g769 ( .A1(n_705), .A2(n_83), .B(n_82), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_612), .B(n_37), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_690), .A2(n_87), .B(n_86), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_695), .Y(n_772) );
INVx3_ASAP7_75t_L g773 ( .A(n_595), .Y(n_773) );
OAI21x1_ASAP7_75t_L g774 ( .A1(n_673), .A2(n_160), .B(n_276), .Y(n_774) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_691), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_SL g776 ( .A1(n_618), .A2(n_158), .B(n_275), .C(n_273), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_695), .Y(n_777) );
OA21x2_ASAP7_75t_L g778 ( .A1(n_662), .A2(n_157), .B(n_268), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_667), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_592), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_682), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_611), .B(n_38), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_607), .B(n_39), .Y(n_783) );
AO21x2_ASAP7_75t_L g784 ( .A1(n_709), .A2(n_156), .B(n_267), .Y(n_784) );
AOI21xp33_ASAP7_75t_L g785 ( .A1(n_636), .A2(n_39), .B(n_40), .Y(n_785) );
AO31x2_ASAP7_75t_L g786 ( .A1(n_677), .A2(n_41), .A3(n_42), .B(n_43), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_673), .A2(n_166), .B(n_266), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_607), .Y(n_788) );
BUFx2_ASAP7_75t_L g789 ( .A(n_599), .Y(n_789) );
OA21x2_ASAP7_75t_L g790 ( .A1(n_646), .A2(n_165), .B(n_263), .Y(n_790) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_676), .A2(n_152), .B(n_259), .Y(n_791) );
BUFx3_ASAP7_75t_L g792 ( .A(n_595), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_615), .B(n_42), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_708), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_683), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_650), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_694), .Y(n_797) );
OA21x2_ASAP7_75t_L g798 ( .A1(n_676), .A2(n_150), .B(n_258), .Y(n_798) );
INVx3_ASAP7_75t_SL g799 ( .A(n_634), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_641), .Y(n_800) );
BUFx3_ASAP7_75t_L g801 ( .A(n_649), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_679), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_687), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_675), .B(n_43), .Y(n_804) );
INVx2_ASAP7_75t_SL g805 ( .A(n_588), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_704), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_589), .A2(n_168), .B(n_257), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_622), .B(n_44), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_623), .Y(n_809) );
AND2x4_ASAP7_75t_L g810 ( .A(n_627), .B(n_44), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_629), .B(n_45), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_643), .A2(n_147), .B(n_256), .Y(n_812) );
INVx3_ASAP7_75t_L g813 ( .A(n_649), .Y(n_813) );
OAI21x1_ASAP7_75t_L g814 ( .A1(n_657), .A2(n_140), .B(n_252), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_659), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_669), .A2(n_138), .B(n_247), .Y(n_816) );
OA21x2_ASAP7_75t_L g817 ( .A1(n_681), .A2(n_137), .B(n_243), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_688), .Y(n_818) );
AND2x4_ASAP7_75t_L g819 ( .A(n_627), .B(n_45), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_658), .A2(n_169), .B(n_242), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_658), .A2(n_133), .B(n_241), .Y(n_821) );
AO21x2_ASAP7_75t_L g822 ( .A1(n_709), .A2(n_128), .B(n_239), .Y(n_822) );
OR2x2_ASAP7_75t_L g823 ( .A(n_686), .B(n_625), .Y(n_823) );
A2O1A1Ixp33_ASAP7_75t_L g824 ( .A1(n_610), .A2(n_46), .B(n_47), .C(n_48), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_609), .A2(n_126), .B(n_238), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_602), .A2(n_123), .B(n_237), .Y(n_826) );
OAI21x1_ASAP7_75t_L g827 ( .A1(n_602), .A2(n_122), .B(n_236), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_619), .B(n_46), .Y(n_828) );
BUFx3_ASAP7_75t_L g829 ( .A(n_649), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_665), .B(n_47), .Y(n_830) );
AO21x1_ASAP7_75t_L g831 ( .A1(n_639), .A2(n_170), .B(n_234), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_688), .Y(n_832) );
AND2x4_ASAP7_75t_L g833 ( .A(n_670), .B(n_49), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_655), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_588), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_648), .Y(n_836) );
A2O1A1Ixp33_ASAP7_75t_L g837 ( .A1(n_645), .A2(n_51), .B(n_52), .C(n_53), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_668), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_838) );
OAI21x1_ASAP7_75t_L g839 ( .A1(n_637), .A2(n_180), .B(n_233), .Y(n_839) );
AO21x2_ASAP7_75t_L g840 ( .A1(n_651), .A2(n_179), .B(n_231), .Y(n_840) );
AO21x2_ASAP7_75t_L g841 ( .A1(n_651), .A2(n_172), .B(n_229), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_608), .Y(n_842) );
O2A1O1Ixp33_ASAP7_75t_L g843 ( .A1(n_644), .A2(n_55), .B(n_56), .C(n_57), .Y(n_843) );
AOI21x1_ASAP7_75t_L g844 ( .A1(n_736), .A2(n_601), .B(n_656), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_745), .A2(n_727), .B1(n_804), .B2(n_828), .Y(n_845) );
NAND2xp33_ASAP7_75t_L g846 ( .A(n_842), .B(n_608), .Y(n_846) );
OAI21xp33_ASAP7_75t_SL g847 ( .A1(n_762), .A2(n_640), .B(n_674), .Y(n_847) );
BUFx2_ASAP7_75t_L g848 ( .A(n_711), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_711), .B(n_587), .Y(n_849) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_747), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_745), .A2(n_656), .B1(n_672), .B2(n_693), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_747), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g853 ( .A(n_763), .B(n_635), .C(n_633), .Y(n_853) );
AOI22xp5_ASAP7_75t_SL g854 ( .A1(n_716), .A2(n_653), .B1(n_671), .B2(n_680), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_781), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g856 ( .A1(n_721), .A2(n_699), .B(n_696), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_727), .A2(n_654), .B1(n_653), .B2(n_671), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_720), .Y(n_858) );
OAI21xp5_ASAP7_75t_L g859 ( .A1(n_779), .A2(n_670), .B(n_680), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_781), .Y(n_860) );
A2O1A1Ixp33_ASAP7_75t_L g861 ( .A1(n_808), .A2(n_670), .B(n_680), .C(n_689), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_804), .A2(n_699), .B1(n_696), .B2(n_689), .Y(n_862) );
OAI211xp5_ASAP7_75t_L g863 ( .A1(n_838), .A2(n_699), .B(n_696), .C(n_689), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_726), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_730), .A2(n_688), .B(n_608), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_823), .A2(n_608), .B1(n_59), .B2(n_60), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_796), .B(n_608), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g868 ( .A(n_712), .B(n_58), .C(n_59), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_733), .Y(n_869) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_801), .Y(n_870) );
AOI31xp33_ASAP7_75t_L g871 ( .A1(n_838), .A2(n_58), .A3(n_60), .B(n_61), .Y(n_871) );
AOI21xp33_ASAP7_75t_L g872 ( .A1(n_808), .A2(n_61), .B(n_62), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_795), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_741), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_874) );
OAI222xp33_ASAP7_75t_L g875 ( .A1(n_766), .A2(n_63), .B1(n_64), .B2(n_65), .C1(n_88), .C2(n_89), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_795), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_732), .B(n_90), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_735), .B(n_91), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_732), .B(n_94), .Y(n_879) );
NOR2x1_ASAP7_75t_SL g880 ( .A(n_801), .B(n_95), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_743), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_744), .Y(n_882) );
OAI22xp5_ASAP7_75t_SL g883 ( .A1(n_716), .A2(n_97), .B1(n_99), .B2(n_103), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_750), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_772), .A2(n_107), .B1(n_108), .B2(n_110), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_788), .A2(n_112), .B1(n_116), .B2(n_117), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_766), .A2(n_118), .B1(n_119), .B2(n_120), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_753), .B(n_121), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_732), .B(n_182), .Y(n_889) );
AOI222xp33_ASAP7_75t_L g890 ( .A1(n_712), .A2(n_183), .B1(n_186), .B2(n_188), .C1(n_191), .C2(n_193), .Y(n_890) );
INVxp67_ASAP7_75t_L g891 ( .A(n_761), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_768), .B(n_195), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_754), .B(n_196), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_761), .B(n_201), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_796), .B(n_202), .Y(n_895) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_718), .A2(n_203), .B(n_204), .Y(n_896) );
A2O1A1Ixp33_ASAP7_75t_L g897 ( .A1(n_755), .A2(n_206), .B(n_207), .C(n_208), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_765), .B(n_728), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_806), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_797), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_761), .Y(n_901) );
AOI221xp5_ASAP7_75t_L g902 ( .A1(n_715), .A2(n_210), .B1(n_211), .B2(n_212), .C(n_213), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_734), .A2(n_214), .B1(n_216), .B2(n_217), .Y(n_903) );
AOI21xp5_ASAP7_75t_L g904 ( .A1(n_710), .A2(n_218), .B(n_219), .Y(n_904) );
AOI21xp5_ASAP7_75t_SL g905 ( .A1(n_833), .A2(n_220), .B(n_221), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_802), .Y(n_906) );
AOI222xp33_ASAP7_75t_L g907 ( .A1(n_830), .A2(n_222), .B1(n_223), .B2(n_224), .C1(n_228), .C2(n_278), .Y(n_907) );
AOI221xp5_ASAP7_75t_L g908 ( .A1(n_755), .A2(n_758), .B1(n_760), .B2(n_785), .C(n_830), .Y(n_908) );
OA21x2_ASAP7_75t_L g909 ( .A1(n_749), .A2(n_725), .B(n_722), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_748), .A2(n_770), .B(n_757), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_782), .A2(n_729), .B1(n_783), .B2(n_811), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_809), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_729), .A2(n_793), .B1(n_819), .B2(n_810), .Y(n_913) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_775), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_810), .A2(n_819), .B1(n_764), .B2(n_833), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_803), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_833), .A2(n_777), .B1(n_800), .B2(n_724), .Y(n_917) );
AOI222xp33_ASAP7_75t_L g918 ( .A1(n_836), .A2(n_789), .B1(n_799), .B2(n_767), .C1(n_837), .C2(n_780), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_775), .A2(n_834), .B1(n_731), .B2(n_799), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_815), .A2(n_717), .B1(n_840), .B2(n_841), .Y(n_920) );
AND2x4_ASAP7_75t_L g921 ( .A(n_723), .B(n_756), .Y(n_921) );
INVx4_ASAP7_75t_L g922 ( .A(n_842), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_843), .A2(n_824), .B1(n_837), .B2(n_805), .C(n_780), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_815), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_717), .A2(n_840), .B1(n_841), .B2(n_817), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_835), .B(n_746), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_786), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_835), .Y(n_928) );
AOI22xp5_ASAP7_75t_SL g929 ( .A1(n_836), .A2(n_794), .B1(n_790), .B2(n_817), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_794), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_824), .A2(n_829), .B1(n_843), .B2(n_792), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_786), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_717), .A2(n_759), .B(n_719), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_829), .A2(n_792), .B1(n_813), .B2(n_773), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_813), .A2(n_773), .B1(n_739), .B2(n_817), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_739), .B(n_786), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_825), .A2(n_776), .B1(n_771), .B2(n_769), .C(n_831), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_786), .B(n_740), .Y(n_938) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_719), .A2(n_742), .B1(n_776), .B2(n_790), .C(n_752), .Y(n_939) );
AO21x2_ASAP7_75t_L g940 ( .A1(n_784), .A2(n_822), .B(n_751), .Y(n_940) );
OAI21x1_ASAP7_75t_L g941 ( .A1(n_738), .A2(n_807), .B(n_812), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_740), .Y(n_942) );
OAI211xp5_ASAP7_75t_SL g943 ( .A1(n_740), .A2(n_832), .B(n_818), .C(n_790), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_818), .B(n_832), .Y(n_944) );
AND2x4_ASAP7_75t_L g945 ( .A(n_737), .B(n_839), .Y(n_945) );
OR2x2_ASAP7_75t_L g946 ( .A(n_742), .B(n_784), .Y(n_946) );
AND2x4_ASAP7_75t_L g947 ( .A(n_826), .B(n_827), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_742), .B(n_822), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_778), .A2(n_752), .B1(n_798), .B2(n_740), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_778), .B(n_752), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_778), .B(n_714), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_798), .A2(n_821), .B1(n_820), .B2(n_713), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_774), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_798), .B(n_787), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_791), .A2(n_745), .B1(n_727), .B2(n_804), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g956 ( .A1(n_814), .A2(n_596), .B1(n_707), .B2(n_562), .C(n_594), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_816), .A2(n_745), .B1(n_727), .B2(n_804), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_727), .A2(n_600), .B1(n_605), .B2(n_583), .Y(n_958) );
OAI211xp5_ASAP7_75t_L g959 ( .A1(n_745), .A2(n_646), .B(n_550), .C(n_628), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_779), .B(n_598), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_745), .A2(n_727), .B1(n_804), .B2(n_828), .Y(n_961) );
INVx3_ASAP7_75t_L g962 ( .A(n_945), .Y(n_962) );
BUFx3_ASAP7_75t_L g963 ( .A(n_848), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_850), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_852), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_850), .B(n_855), .Y(n_966) );
AND2x4_ASAP7_75t_L g967 ( .A(n_901), .B(n_891), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_927), .Y(n_968) );
OAI321xp33_ASAP7_75t_L g969 ( .A1(n_958), .A2(n_955), .A3(n_957), .B1(n_961), .B2(n_845), .C(n_866), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_932), .Y(n_970) );
INVx3_ASAP7_75t_L g971 ( .A(n_945), .Y(n_971) );
BUFx2_ASAP7_75t_L g972 ( .A(n_891), .Y(n_972) );
INVx4_ASAP7_75t_L g973 ( .A(n_879), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_960), .B(n_959), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_869), .Y(n_975) );
AOI221x1_ASAP7_75t_L g976 ( .A1(n_943), .A2(n_949), .B1(n_933), .B2(n_868), .C(n_935), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_914), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_860), .B(n_873), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_876), .Y(n_979) );
BUFx2_ASAP7_75t_L g980 ( .A(n_847), .Y(n_980) );
HB1xp67_ASAP7_75t_L g981 ( .A(n_914), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_881), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_915), .B(n_942), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_882), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_900), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_912), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g987 ( .A(n_890), .B(n_868), .C(n_955), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_924), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_879), .B(n_906), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_915), .B(n_913), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_865), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_858), .B(n_845), .Y(n_992) );
INVxp67_ASAP7_75t_L g993 ( .A(n_926), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_916), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_877), .B(n_889), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_936), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_938), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_961), .B(n_913), .Y(n_998) );
INVx2_ASAP7_75t_L g999 ( .A(n_865), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_944), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_921), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_894), .B(n_899), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_921), .Y(n_1003) );
INVx3_ASAP7_75t_L g1004 ( .A(n_870), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_923), .B(n_911), .Y(n_1005) );
CKINVDCx16_ASAP7_75t_R g1006 ( .A(n_928), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_898), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_918), .B(n_874), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_874), .B(n_864), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_859), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_854), .B(n_911), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_849), .B(n_908), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_953), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_947), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_947), .Y(n_1015) );
AO21x2_ASAP7_75t_L g1016 ( .A1(n_948), .A2(n_951), .B(n_939), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_919), .B(n_851), .Y(n_1017) );
INVx3_ASAP7_75t_L g1018 ( .A(n_870), .Y(n_1018) );
INVxp67_ASAP7_75t_L g1019 ( .A(n_895), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_878), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_888), .Y(n_1021) );
BUFx3_ASAP7_75t_L g1022 ( .A(n_870), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_922), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_851), .B(n_892), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_893), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_946), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_919), .B(n_956), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_917), .B(n_957), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_867), .B(n_892), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_909), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_917), .B(n_870), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_853), .B(n_872), .Y(n_1032) );
INVx3_ASAP7_75t_L g1033 ( .A(n_922), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_853), .B(n_862), .Y(n_1034) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_934), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_941), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_862), .B(n_929), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_954), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_857), .A2(n_871), .B1(n_887), .B2(n_903), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_880), .Y(n_1040) );
INVx4_ASAP7_75t_L g1041 ( .A(n_950), .Y(n_1041) );
AO31x2_ASAP7_75t_L g1042 ( .A1(n_952), .A2(n_910), .A3(n_931), .B(n_897), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1043 ( .A(n_930), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_940), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_887), .B(n_857), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_940), .Y(n_1046) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_861), .Y(n_1047) );
INVx3_ASAP7_75t_L g1048 ( .A(n_844), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_905), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_920), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_907), .B(n_920), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_925), .B(n_863), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_903), .B(n_846), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_925), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_885), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_886), .B(n_902), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_883), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_997), .B(n_886), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_968), .Y(n_1059) );
AOI33xp33_ASAP7_75t_L g1060 ( .A1(n_1008), .A2(n_884), .A3(n_937), .B1(n_875), .B2(n_896), .B3(n_904), .Y(n_1060) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_963), .Y(n_1061) );
INVx1_ASAP7_75t_SL g1062 ( .A(n_1006), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1007), .B(n_884), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_1008), .A2(n_856), .B1(n_1051), .B2(n_987), .Y(n_1064) );
INVx5_ASAP7_75t_SL g1065 ( .A(n_967), .Y(n_1065) );
INVx2_ASAP7_75t_SL g1066 ( .A(n_963), .Y(n_1066) );
AO21x2_ASAP7_75t_L g1067 ( .A1(n_1044), .A2(n_1046), .B(n_1036), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_997), .B(n_966), .Y(n_1068) );
OAI33xp33_ASAP7_75t_L g1069 ( .A1(n_1012), .A2(n_1057), .A3(n_974), .B1(n_1005), .B2(n_994), .B3(n_1039), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_966), .B(n_1041), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_968), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_1041), .B(n_1031), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_983), .B(n_964), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1041), .B(n_1038), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1041), .B(n_1038), .Y(n_1075) );
NAND4xp25_ASAP7_75t_L g1076 ( .A(n_987), .B(n_1032), .C(n_1017), .D(n_990), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_983), .B(n_964), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_994), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_973), .Y(n_1079) );
INVx3_ASAP7_75t_L g1080 ( .A(n_973), .Y(n_1080) );
INVx3_ASAP7_75t_L g1081 ( .A(n_973), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1007), .B(n_1009), .Y(n_1082) );
OAI21xp33_ASAP7_75t_L g1083 ( .A1(n_1032), .A2(n_1011), .B(n_1028), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_977), .B(n_981), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1026), .B(n_1054), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_1028), .B(n_990), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1009), .B(n_992), .Y(n_1087) );
OR2x6_ASAP7_75t_L g1088 ( .A(n_973), .B(n_1035), .Y(n_1088) );
BUFx3_ASAP7_75t_L g1089 ( .A(n_1033), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1030), .Y(n_1090) );
OAI221xp5_ASAP7_75t_L g1091 ( .A1(n_1019), .A2(n_1027), .B1(n_1029), .B2(n_998), .C(n_993), .Y(n_1091) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1001), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1002), .B(n_975), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_970), .Y(n_1094) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_1034), .B(n_1003), .C(n_1040), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1006), .B(n_1043), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1026), .B(n_1054), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_969), .A2(n_984), .B1(n_982), .B2(n_975), .C(n_1002), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_978), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1100 ( .A(n_996), .B(n_970), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_978), .B(n_982), .Y(n_1101) );
INVx4_ASAP7_75t_L g1102 ( .A(n_1033), .Y(n_1102) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_1033), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_996), .B(n_1050), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_1011), .A2(n_995), .B1(n_1051), .B2(n_1024), .Y(n_1105) );
INVx1_ASAP7_75t_SL g1106 ( .A(n_1043), .Y(n_1106) );
BUFx2_ASAP7_75t_L g1107 ( .A(n_962), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_984), .B(n_965), .Y(n_1108) );
INVx4_ASAP7_75t_L g1109 ( .A(n_1033), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_965), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1013), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1013), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1050), .B(n_988), .Y(n_1113) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_979), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_986), .B(n_988), .Y(n_1115) );
AO21x2_ASAP7_75t_L g1116 ( .A1(n_991), .A2(n_999), .B(n_1016), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1000), .B(n_1010), .Y(n_1117) );
AO21x2_ASAP7_75t_L g1118 ( .A1(n_991), .A2(n_999), .B(n_1016), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1119 ( .A(n_989), .B(n_1023), .Y(n_1119) );
INVx1_ASAP7_75t_SL g1120 ( .A(n_1022), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_985), .B(n_1031), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_1010), .B(n_1015), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_989), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1014), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_962), .Y(n_1125) );
NAND2x1p5_ASAP7_75t_SL g1126 ( .A(n_1049), .B(n_1056), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_1024), .A2(n_1045), .B1(n_1020), .B2(n_1025), .C(n_1021), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1014), .B(n_1015), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1037), .B(n_962), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1101), .B(n_1093), .Y(n_1130) );
NAND2x1_ASAP7_75t_L g1131 ( .A(n_1102), .B(n_962), .Y(n_1131) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1090), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1059), .Y(n_1133) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_1110), .Y(n_1134) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_1061), .Y(n_1135) );
NOR3xp33_ASAP7_75t_L g1136 ( .A(n_1069), .B(n_1025), .C(n_1021), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1121), .B(n_971), .Y(n_1137) );
NOR2x1_ASAP7_75t_L g1138 ( .A(n_1102), .B(n_1047), .Y(n_1138) );
NOR2xp33_ASAP7_75t_SL g1139 ( .A(n_1102), .B(n_995), .Y(n_1139) );
INVx3_ASAP7_75t_L g1140 ( .A(n_1109), .Y(n_1140) );
OAI33xp33_ASAP7_75t_L g1141 ( .A1(n_1105), .A2(n_1020), .A3(n_1052), .B1(n_1053), .B2(n_1055), .B3(n_1049), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1121), .B(n_971), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1086), .B(n_971), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1129), .B(n_971), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1101), .B(n_1045), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1059), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1129), .B(n_980), .Y(n_1147) );
NOR3xp33_ASAP7_75t_L g1148 ( .A(n_1091), .B(n_1047), .C(n_1056), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1074), .B(n_980), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_1076), .A2(n_1037), .B1(n_972), .B2(n_967), .C(n_1035), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1071), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1099), .B(n_967), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_1083), .A2(n_1055), .B1(n_972), .B2(n_1052), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1068), .B(n_1004), .Y(n_1154) );
NOR2xp33_ASAP7_75t_L g1155 ( .A(n_1062), .B(n_1022), .Y(n_1155) );
INVx2_ASAP7_75t_SL g1156 ( .A(n_1109), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1157 ( .A(n_1074), .B(n_1048), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1075), .B(n_1016), .Y(n_1158) );
NAND3xp33_ASAP7_75t_L g1159 ( .A(n_1098), .B(n_976), .C(n_1048), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1075), .B(n_1048), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1070), .B(n_1048), .Y(n_1161) );
NOR3xp33_ASAP7_75t_L g1162 ( .A(n_1095), .B(n_1004), .C(n_1018), .Y(n_1162) );
AND2x4_ASAP7_75t_SL g1163 ( .A(n_1109), .B(n_1004), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_1106), .B(n_1018), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1071), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1070), .B(n_1042), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1068), .B(n_1042), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1094), .Y(n_1168) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1116), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1094), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1066), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1172 ( .A(n_1089), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1085), .B(n_1042), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1111), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1111), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_1096), .Y(n_1176) );
AND2x4_ASAP7_75t_SL g1177 ( .A(n_1088), .B(n_1018), .Y(n_1177) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1067), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1085), .B(n_1042), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1066), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1112), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1086), .B(n_1042), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1082), .B(n_976), .Y(n_1183) );
AOI221xp5_ASAP7_75t_L g1184 ( .A1(n_1127), .A2(n_1064), .B1(n_1123), .B2(n_1119), .C(n_1087), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1097), .B(n_1128), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1073), .B(n_1077), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1185), .B(n_1097), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1166), .B(n_1128), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1133), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1133), .Y(n_1190) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_1140), .Y(n_1191) );
OAI32xp33_ASAP7_75t_L g1192 ( .A1(n_1148), .A2(n_1084), .A3(n_1117), .B1(n_1089), .B2(n_1103), .Y(n_1192) );
INVx1_ASAP7_75t_SL g1193 ( .A(n_1135), .Y(n_1193) );
XOR2xp5_ASAP7_75t_L g1194 ( .A(n_1176), .B(n_1084), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1186), .B(n_1077), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1146), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1166), .B(n_1072), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1185), .B(n_1117), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1167), .B(n_1072), .Y(n_1199) );
INVx3_ASAP7_75t_SL g1200 ( .A(n_1140), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_1134), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1146), .Y(n_1202) );
NOR2xp33_ASAP7_75t_L g1203 ( .A(n_1130), .B(n_1092), .Y(n_1203) );
INVx1_ASAP7_75t_SL g1204 ( .A(n_1171), .Y(n_1204) );
NOR2xp33_ASAP7_75t_L g1205 ( .A(n_1155), .B(n_1078), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1145), .B(n_1113), .Y(n_1206) );
NAND2xp5_ASAP7_75t_SL g1207 ( .A(n_1139), .B(n_1103), .Y(n_1207) );
NOR2x1_ASAP7_75t_L g1208 ( .A(n_1140), .B(n_1081), .Y(n_1208) );
OAI222xp33_ASAP7_75t_L g1209 ( .A1(n_1156), .A2(n_1088), .B1(n_1079), .B2(n_1072), .C1(n_1080), .C2(n_1081), .Y(n_1209) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1132), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1132), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1186), .B(n_1113), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1143), .B(n_1073), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1167), .B(n_1124), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1158), .B(n_1124), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1151), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1132), .Y(n_1217) );
OR2x6_ASAP7_75t_L g1218 ( .A(n_1131), .B(n_1088), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1158), .B(n_1112), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1184), .B(n_1108), .Y(n_1220) );
INVxp67_ASAP7_75t_L g1221 ( .A(n_1180), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1151), .B(n_1108), .Y(n_1222) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_1156), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1137), .B(n_1107), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1137), .B(n_1142), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1142), .B(n_1107), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1165), .Y(n_1227) );
INVx1_ASAP7_75t_SL g1228 ( .A(n_1140), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1165), .B(n_1115), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1143), .B(n_1122), .Y(n_1230) );
AOI222xp33_ASAP7_75t_L g1231 ( .A1(n_1220), .A2(n_1141), .B1(n_1150), .B2(n_1179), .C1(n_1173), .C2(n_1147), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1219), .B(n_1183), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1201), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1234 ( .A1(n_1205), .A2(n_1136), .B1(n_1153), .B2(n_1161), .Y(n_1234) );
INVxp67_ASAP7_75t_SL g1235 ( .A(n_1223), .Y(n_1235) );
OAI322xp33_ASAP7_75t_L g1236 ( .A1(n_1195), .A2(n_1182), .A3(n_1152), .B1(n_1154), .B2(n_1122), .C1(n_1168), .C2(n_1175), .Y(n_1236) );
AOI211xp5_ASAP7_75t_L g1237 ( .A1(n_1192), .A2(n_1159), .B(n_1182), .C(n_1164), .Y(n_1237) );
OAI321xp33_ASAP7_75t_L g1238 ( .A1(n_1218), .A2(n_1159), .A3(n_1088), .B1(n_1179), .B2(n_1173), .C(n_1147), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1195), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1219), .B(n_1181), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_1221), .A2(n_1138), .B1(n_1162), .B2(n_1063), .C(n_1131), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1198), .B(n_1149), .Y(n_1242) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1210), .Y(n_1243) );
AOI322xp5_ASAP7_75t_L g1244 ( .A1(n_1203), .A2(n_1149), .A3(n_1144), .B1(n_1161), .B2(n_1138), .C1(n_1181), .C2(n_1170), .Y(n_1244) );
AOI21xp5_ASAP7_75t_L g1245 ( .A1(n_1192), .A2(n_1163), .B(n_1172), .Y(n_1245) );
INVx3_ASAP7_75t_L g1246 ( .A(n_1200), .Y(n_1246) );
AOI211xp5_ASAP7_75t_L g1247 ( .A1(n_1200), .A2(n_1144), .B(n_1079), .C(n_1172), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1225), .B(n_1160), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1189), .Y(n_1249) );
OAI222xp33_ASAP7_75t_L g1250 ( .A1(n_1218), .A2(n_1125), .B1(n_1100), .B2(n_1160), .C1(n_1157), .C2(n_1174), .Y(n_1250) );
AOI222xp33_ASAP7_75t_L g1251 ( .A1(n_1188), .A2(n_1168), .B1(n_1170), .B2(n_1174), .C1(n_1058), .C2(n_1157), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1225), .B(n_1157), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_1194), .A2(n_1065), .B1(n_1080), .B2(n_1081), .Y(n_1253) );
A2O1A1Ixp33_ASAP7_75t_L g1254 ( .A1(n_1207), .A2(n_1208), .B(n_1191), .C(n_1228), .Y(n_1254) );
INVxp67_ASAP7_75t_L g1255 ( .A(n_1191), .Y(n_1255) );
OAI21xp33_ASAP7_75t_L g1256 ( .A1(n_1193), .A2(n_1060), .B(n_1169), .Y(n_1256) );
INVx1_ASAP7_75t_SL g1257 ( .A(n_1233), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1231), .B(n_1188), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_1247), .A2(n_1194), .B1(n_1200), .B2(n_1218), .Y(n_1259) );
NAND4xp75_ASAP7_75t_L g1260 ( .A(n_1245), .B(n_1208), .C(n_1197), .D(n_1199), .Y(n_1260) );
OAI21xp33_ASAP7_75t_L g1261 ( .A1(n_1244), .A2(n_1204), .B(n_1193), .Y(n_1261) );
AOI221xp5_ASAP7_75t_SL g1262 ( .A1(n_1236), .A2(n_1187), .B1(n_1212), .B2(n_1206), .C(n_1209), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1249), .Y(n_1263) );
XNOR2x1_ASAP7_75t_L g1264 ( .A(n_1234), .B(n_1213), .Y(n_1264) );
INVx1_ASAP7_75t_SL g1265 ( .A(n_1246), .Y(n_1265) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1243), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1251), .B(n_1214), .Y(n_1267) );
INVx1_ASAP7_75t_SL g1268 ( .A(n_1246), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1239), .Y(n_1269) );
AOI222xp33_ASAP7_75t_L g1270 ( .A1(n_1256), .A2(n_1224), .B1(n_1226), .B2(n_1229), .C1(n_1214), .C2(n_1215), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1232), .B(n_1230), .Y(n_1271) );
AOI211xp5_ASAP7_75t_L g1272 ( .A1(n_1254), .A2(n_1228), .B(n_1230), .C(n_1226), .Y(n_1272) );
XOR2x2_ASAP7_75t_L g1273 ( .A(n_1253), .B(n_1215), .Y(n_1273) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1243), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1263), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_1272), .A2(n_1254), .B1(n_1235), .B2(n_1241), .Y(n_1276) );
OAI22xp33_ASAP7_75t_L g1277 ( .A1(n_1259), .A2(n_1238), .B1(n_1218), .B2(n_1255), .Y(n_1277) );
AOI222xp33_ASAP7_75t_L g1278 ( .A1(n_1258), .A2(n_1255), .B1(n_1250), .B2(n_1240), .C1(n_1248), .C2(n_1222), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1262), .B(n_1242), .Y(n_1279) );
AOI21xp33_ASAP7_75t_SL g1280 ( .A1(n_1261), .A2(n_1218), .B(n_1126), .Y(n_1280) );
OAI311xp33_ASAP7_75t_L g1281 ( .A1(n_1270), .A2(n_1237), .A3(n_1104), .B1(n_1169), .C1(n_1250), .Y(n_1281) );
OAI211xp5_ASAP7_75t_SL g1282 ( .A1(n_1267), .A2(n_1268), .B(n_1265), .C(n_1257), .Y(n_1282) );
XOR2xp5_ASAP7_75t_L g1283 ( .A(n_1264), .B(n_1252), .Y(n_1283) );
A2O1A1Ixp33_ASAP7_75t_SL g1284 ( .A1(n_1269), .A2(n_1169), .B(n_1178), .C(n_1080), .Y(n_1284) );
NAND3xp33_ASAP7_75t_SL g1285 ( .A(n_1280), .B(n_1260), .C(n_1271), .Y(n_1285) );
INVx1_ASAP7_75t_SL g1286 ( .A(n_1279), .Y(n_1286) );
AOI21xp33_ASAP7_75t_SL g1287 ( .A1(n_1277), .A2(n_1126), .B(n_1273), .Y(n_1287) );
AOI22xp5_ASAP7_75t_L g1288 ( .A1(n_1282), .A2(n_1274), .B1(n_1266), .B2(n_1227), .Y(n_1288) );
OAI221xp5_ASAP7_75t_L g1289 ( .A1(n_1278), .A2(n_1266), .B1(n_1274), .B2(n_1202), .C(n_1216), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1275), .B(n_1196), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1291 ( .A(n_1286), .B(n_1283), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1288), .B(n_1276), .Y(n_1292) );
NAND2xp5_ASAP7_75t_SL g1293 ( .A(n_1287), .B(n_1277), .Y(n_1293) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_1290), .Y(n_1294) );
OAI221xp5_ASAP7_75t_SL g1295 ( .A1(n_1292), .A2(n_1289), .B1(n_1285), .B2(n_1281), .C(n_1284), .Y(n_1295) );
AOI21xp5_ASAP7_75t_SL g1296 ( .A1(n_1293), .A2(n_1114), .B(n_1115), .Y(n_1296) );
NOR3xp33_ASAP7_75t_L g1297 ( .A(n_1291), .B(n_1120), .C(n_1190), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1297), .B(n_1294), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1296), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1298), .Y(n_1300) );
OR2x6_ASAP7_75t_L g1301 ( .A(n_1299), .B(n_1295), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1300), .Y(n_1302) );
OAI22x1_ASAP7_75t_L g1303 ( .A1(n_1301), .A2(n_1125), .B1(n_1058), .B2(n_1217), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_1302), .A2(n_1177), .B1(n_1217), .B2(n_1211), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_1304), .A2(n_1303), .B1(n_1116), .B2(n_1118), .Y(n_1305) );
AOI22xp5_ASAP7_75t_L g1306 ( .A1(n_1305), .A2(n_1065), .B1(n_1118), .B2(n_1116), .Y(n_1306) );
endmodule