module fake_jpeg_40_n_527 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_57),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_19),
.B(n_8),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_70),
.Y(n_120)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_90),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_29),
.B(n_7),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_50),
.B(n_7),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_97),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_24),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_21),
.B(n_10),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_30),
.B(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_30),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_12),
.Y(n_175)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_18),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_34),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_108),
.B(n_121),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_24),
.B1(n_28),
.B2(n_51),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_112),
.A2(n_147),
.B1(n_35),
.B2(n_41),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_32),
.B1(n_26),
.B2(n_27),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_32),
.B1(n_26),
.B2(n_27),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_39),
.B(n_51),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_22),
.B1(n_24),
.B2(n_48),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_62),
.B(n_52),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_129),
.B(n_175),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_76),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_22),
.B1(n_48),
.B2(n_46),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_32),
.B1(n_34),
.B2(n_28),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_54),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_161),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_105),
.A2(n_60),
.B1(n_65),
.B2(n_96),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_86),
.B1(n_77),
.B2(n_79),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_69),
.A2(n_46),
.B1(n_34),
.B2(n_47),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_74),
.B1(n_82),
.B2(n_107),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_56),
.B(n_46),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_57),
.A2(n_52),
.B1(n_36),
.B2(n_44),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_94),
.B1(n_83),
.B2(n_106),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_58),
.B(n_44),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_63),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_75),
.B(n_36),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_164),
.B(n_1),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_58),
.B(n_47),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_73),
.B(n_34),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_167),
.B(n_1),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_12),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_72),
.Y(n_197)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_123),
.A2(n_67),
.B1(n_71),
.B2(n_87),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_178),
.A2(n_193),
.B1(n_201),
.B2(n_131),
.Y(n_249)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_160),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_189),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_184),
.A2(n_217),
.B1(n_122),
.B2(n_119),
.Y(n_268)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_185),
.Y(n_255)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_187),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_84),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_160),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_120),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_190),
.B(n_192),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_73),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_204),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_194),
.A2(n_219),
.B1(n_230),
.B2(n_139),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_130),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_220),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_197),
.B(n_205),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_13),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_110),
.B(n_0),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_137),
.B(n_14),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_126),
.B(n_0),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_234),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_112),
.A2(n_81),
.B(n_78),
.C(n_35),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_208),
.A2(n_236),
.B(n_2),
.C(n_221),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_136),
.B(n_0),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_227),
.Y(n_275)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_109),
.Y(n_216)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_147),
.A2(n_11),
.B1(n_15),
.B2(n_12),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_113),
.B(n_11),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g221 ( 
.A(n_109),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_221),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_140),
.A2(n_41),
.B(n_25),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_222),
.A2(n_195),
.B(n_236),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_232),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_114),
.B(n_1),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_228),
.Y(n_291)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_229),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_116),
.A2(n_41),
.B1(n_25),
.B2(n_11),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_124),
.B(n_169),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_125),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_239),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_142),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_142),
.B(n_134),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_237),
.Y(n_260)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_128),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_154),
.B(n_15),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_15),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_181),
.A2(n_158),
.B1(n_170),
.B2(n_155),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_242),
.A2(n_243),
.B1(n_279),
.B2(n_284),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_170),
.B1(n_158),
.B2(n_176),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_176),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_246),
.B(n_264),
.C(n_179),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_249),
.A2(n_259),
.B1(n_268),
.B2(n_270),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_198),
.A2(n_145),
.B1(n_131),
.B2(n_125),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_SL g261 ( 
.A(n_191),
.B(n_150),
.C(n_173),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_282),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_190),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_277),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_212),
.B(n_145),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_184),
.A2(n_115),
.B1(n_174),
.B2(n_143),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_180),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_193),
.A2(n_122),
.B1(n_151),
.B2(n_119),
.Y(n_279)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_215),
.A2(n_143),
.A3(n_173),
.B1(n_115),
.B2(n_172),
.Y(n_282)
);

NAND2xp67_ASAP7_75t_L g283 ( 
.A(n_188),
.B(n_128),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_283),
.A2(n_297),
.B(n_274),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_208),
.A2(n_209),
.B1(n_222),
.B2(n_227),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_285),
.B(n_183),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_217),
.A2(n_151),
.B1(n_139),
.B2(n_150),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_219),
.B1(n_185),
.B2(n_189),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_215),
.B(n_172),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_294),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_178),
.A2(n_41),
.B1(n_3),
.B2(n_4),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_195),
.B1(n_196),
.B2(n_185),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_239),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_240),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_234),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_206),
.B(n_186),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

BUFx12_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_300),
.A2(n_321),
.B1(n_255),
.B2(n_243),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_273),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_301),
.B(n_309),
.C(n_318),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_255),
.B1(n_270),
.B2(n_268),
.Y(n_346)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_306),
.Y(n_345)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_207),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_312),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_251),
.Y(n_310)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_246),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_248),
.B(n_188),
.C(n_214),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_317),
.C(n_331),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_314),
.A2(n_315),
.B(n_335),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_236),
.B(n_207),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_248),
.B(n_231),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_241),
.B(n_177),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_269),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_249),
.A2(n_187),
.B1(n_211),
.B2(n_218),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_294),
.B(n_180),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_323),
.B(n_332),
.Y(n_357)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_326),
.B(n_274),
.Y(n_364)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_328),
.A2(n_337),
.B1(n_343),
.B2(n_247),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_264),
.B(n_224),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_330),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_257),
.B(n_226),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_336),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_269),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_342),
.Y(n_382)
);

A2O1A1O1Ixp25_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_200),
.B(n_238),
.C(n_203),
.D(n_229),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_269),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_250),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_257),
.A2(n_225),
.B(n_223),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_341),
.B(n_344),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_276),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_339),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_277),
.A2(n_228),
.B(n_182),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_234),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_280),
.A2(n_202),
.B(n_213),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_342),
.Y(n_347)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_305),
.A2(n_262),
.B1(n_259),
.B2(n_289),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_351),
.A2(n_369),
.B1(n_331),
.B2(n_302),
.Y(n_386)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_340),
.A2(n_262),
.B1(n_286),
.B2(n_282),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_358),
.A2(n_372),
.B1(n_276),
.B2(n_254),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_305),
.A2(n_315),
.B1(n_321),
.B2(n_330),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_360),
.A2(n_371),
.B1(n_322),
.B2(n_313),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_368),
.Y(n_397)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

NAND2xp33_ASAP7_75t_SL g367 ( 
.A(n_324),
.B(n_242),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_367),
.A2(n_265),
.B(n_245),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_312),
.B(n_260),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_305),
.A2(n_260),
.B1(n_274),
.B2(n_295),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_314),
.A2(n_256),
.B(n_283),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_370),
.A2(n_341),
.B(n_344),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_302),
.B1(n_324),
.B2(n_300),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_319),
.A2(n_287),
.B1(n_271),
.B2(n_278),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_266),
.C(n_291),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_379),
.C(n_338),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_306),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_310),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_287),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_322),
.A2(n_336),
.B1(n_334),
.B2(n_310),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_380),
.A2(n_216),
.B1(n_265),
.B2(n_296),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_379),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_386),
.A2(n_390),
.B1(n_399),
.B2(n_402),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_387),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_388),
.A2(n_398),
.B1(n_410),
.B2(n_412),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_329),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_389),
.B(n_396),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_311),
.B1(n_325),
.B2(n_343),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_391),
.A2(n_393),
.B(n_394),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_369),
.A2(n_335),
.B1(n_299),
.B2(n_333),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_355),
.A2(n_298),
.B(n_332),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_404),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_352),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_360),
.A2(n_308),
.B1(n_327),
.B2(n_303),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_328),
.B1(n_316),
.B2(n_307),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_290),
.Y(n_400)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_357),
.B(n_298),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_401),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_361),
.A2(n_339),
.B1(n_278),
.B2(n_337),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_353),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_347),
.B(n_281),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_406),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_378),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_408),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_361),
.B(n_281),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_296),
.C(n_292),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_352),
.C(n_370),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_372),
.A2(n_272),
.B1(n_292),
.B2(n_291),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_414),
.B1(n_354),
.B2(n_356),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_250),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_356),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_210),
.B1(n_254),
.B2(n_252),
.Y(n_414)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_408),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_438),
.C(n_439),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_397),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_368),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_423),
.B(n_425),
.Y(n_450)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_424),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_362),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_359),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_430),
.Y(n_462)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_413),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_382),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_434),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_362),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_389),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_436),
.A2(n_384),
.B1(n_390),
.B2(n_383),
.Y(n_443)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_437),
.A2(n_441),
.B1(n_393),
.B2(n_391),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_382),
.C(n_375),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_348),
.C(n_345),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_371),
.B1(n_355),
.B2(n_348),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_444),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_443),
.A2(n_363),
.B1(n_373),
.B2(n_381),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_432),
.A2(n_410),
.B(n_394),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_447),
.A2(n_429),
.B(n_402),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_423),
.B(n_415),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_453),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_433),
.A2(n_388),
.B1(n_384),
.B2(n_398),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_449),
.A2(n_458),
.B1(n_431),
.B2(n_441),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_418),
.A2(n_395),
.B1(n_392),
.B2(n_386),
.Y(n_451)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_451),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_389),
.C(n_383),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_455),
.C(n_456),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_406),
.C(n_345),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_399),
.C(n_411),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_433),
.A2(n_403),
.B1(n_400),
.B2(n_414),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_367),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_350),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_403),
.C(n_349),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_381),
.C(n_373),
.Y(n_474)
);

A2O1A1O1Ixp25_ASAP7_75t_L g464 ( 
.A1(n_457),
.A2(n_427),
.B(n_434),
.C(n_418),
.D(n_416),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_469),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_465),
.A2(n_478),
.B1(n_374),
.B2(n_350),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_432),
.B(n_438),
.Y(n_467)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_460),
.A2(n_428),
.B1(n_436),
.B2(n_429),
.Y(n_468)
);

AO22x1_ASAP7_75t_L g482 ( 
.A1(n_468),
.A2(n_447),
.B1(n_443),
.B2(n_459),
.Y(n_482)
);

OAI322xp33_ASAP7_75t_L g469 ( 
.A1(n_462),
.A2(n_440),
.A3(n_416),
.B1(n_435),
.B2(n_420),
.C1(n_428),
.C2(n_424),
.Y(n_469)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_454),
.B(n_420),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_472),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_349),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_452),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_475),
.A2(n_464),
.B(n_478),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_480),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_458),
.A2(n_374),
.B1(n_363),
.B2(n_365),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_479),
.B(n_450),
.Y(n_494)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_468),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_484),
.A2(n_465),
.B1(n_468),
.B2(n_475),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_446),
.C(n_456),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_488),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_446),
.C(n_455),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_489),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_463),
.A2(n_449),
.B(n_453),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_490),
.A2(n_491),
.B(n_466),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_463),
.A2(n_450),
.B(n_444),
.Y(n_491)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_492),
.Y(n_499)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_494),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_484),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_500),
.B1(n_482),
.B2(n_490),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_481),
.B(n_474),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_502),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_466),
.C(n_476),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_503),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_476),
.C(n_448),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_483),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_508),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_489),
.C(n_492),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_511),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_485),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_513),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_499),
.A2(n_493),
.B1(n_491),
.B2(n_482),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_507),
.A2(n_496),
.B(n_500),
.C(n_503),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_509),
.Y(n_520)
);

O2A1O1Ixp33_ASAP7_75t_SL g515 ( 
.A1(n_506),
.A2(n_470),
.B(n_480),
.C(n_505),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_515),
.A2(n_508),
.B1(n_498),
.B2(n_513),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_519),
.A2(n_520),
.B(n_521),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_517),
.A2(n_510),
.B(n_502),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_518),
.C(n_516),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_522),
.Y(n_524)
);

O2A1O1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_523),
.B(n_504),
.C(n_365),
.Y(n_525)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_494),
.B(n_252),
.Y(n_526)
);

AOI21x1_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_276),
.B(n_234),
.Y(n_527)
);


endmodule