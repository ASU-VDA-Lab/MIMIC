module real_aes_7209_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_0), .Y(n_452) );
XOR2x2_ASAP7_75t_L g235 ( .A(n_1), .B(n_236), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_2), .A2(n_171), .B1(n_358), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_3), .A2(n_138), .B1(n_266), .B2(n_312), .Y(n_671) );
INVx1_ASAP7_75t_L g665 ( .A(n_4), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g302 ( .A1(n_5), .A2(n_19), .B1(n_179), .B2(n_303), .C1(n_306), .C2(n_311), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_6), .A2(n_191), .B1(n_259), .B2(n_265), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_7), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_8), .A2(n_132), .B1(n_271), .B2(n_297), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_9), .B(n_255), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_10), .A2(n_54), .B1(n_280), .B2(n_283), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_11), .A2(n_318), .B1(n_365), .B2(n_366), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_11), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_12), .A2(n_48), .B1(n_394), .B2(n_396), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_13), .A2(n_574), .B1(n_600), .B2(n_601), .Y(n_573) );
INVx1_ASAP7_75t_L g600 ( .A(n_13), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_14), .A2(n_215), .B1(n_378), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_15), .A2(n_157), .B1(n_386), .B2(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_16), .A2(n_57), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_17), .A2(n_71), .B1(n_311), .B2(n_331), .Y(n_613) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_18), .A2(n_63), .B1(n_244), .B2(n_245), .Y(n_253) );
INVx1_ASAP7_75t_L g656 ( .A(n_18), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_20), .A2(n_115), .B1(n_395), .B2(n_414), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g425 ( .A1(n_21), .A2(n_69), .B1(n_201), .B2(n_308), .C1(n_426), .C2(n_427), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_22), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_23), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_24), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_25), .A2(n_26), .B1(n_239), .B2(n_255), .Y(n_238) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_27), .A2(n_66), .B1(n_244), .B2(n_249), .Y(n_254) );
INVx1_ASAP7_75t_L g657 ( .A(n_27), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_28), .A2(n_187), .B1(n_291), .B2(n_621), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_29), .A2(n_104), .B1(n_470), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_30), .A2(n_53), .B1(n_464), .B2(n_465), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_31), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_32), .A2(n_155), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_33), .A2(n_93), .B1(n_280), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_34), .A2(n_35), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_36), .A2(n_206), .B1(n_306), .B2(n_448), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_37), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_38), .B(n_239), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_39), .Y(n_531) );
INVx1_ASAP7_75t_L g567 ( .A(n_40), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_41), .A2(n_70), .B1(n_472), .B2(n_586), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_42), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_43), .A2(n_154), .B1(n_396), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_44), .A2(n_162), .B1(n_297), .B2(n_364), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_45), .Y(n_532) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_46), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_47), .B(n_420), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_49), .A2(n_205), .B1(n_308), .B2(n_490), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_50), .A2(n_166), .B1(n_297), .B2(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_51), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_52), .B(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_55), .A2(n_144), .B1(n_558), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_56), .A2(n_114), .B1(n_387), .B2(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_58), .A2(n_118), .B1(n_347), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_59), .A2(n_76), .B1(n_362), .B2(n_364), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_60), .A2(n_90), .B1(n_351), .B2(n_390), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_61), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_62), .A2(n_207), .B1(n_256), .B2(n_420), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_64), .A2(n_109), .B1(n_276), .B2(n_299), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_65), .A2(n_131), .B1(n_312), .B2(n_331), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_67), .A2(n_204), .B1(n_351), .B2(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_68), .A2(n_169), .B1(n_289), .B2(n_395), .Y(n_493) );
AND2x2_ASAP7_75t_L g229 ( .A(n_72), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_73), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_74), .A2(n_146), .B1(n_294), .B2(n_364), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_75), .A2(n_159), .B1(n_351), .B2(n_416), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_77), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g226 ( .A(n_78), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_79), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_80), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_81), .A2(n_188), .B1(n_271), .B2(n_276), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_82), .A2(n_110), .B1(n_289), .B2(n_563), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_83), .A2(n_130), .B1(n_291), .B2(n_297), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_84), .A2(n_94), .B1(n_271), .B2(n_364), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_85), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_86), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_87), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_88), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_89), .A2(n_156), .B1(n_358), .B2(n_359), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_91), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_92), .A2(n_124), .B1(n_259), .B2(n_308), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_95), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_96), .A2(n_100), .B1(n_259), .B2(n_265), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_97), .A2(n_172), .B1(n_400), .B2(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_98), .A2(n_435), .B1(n_436), .B2(n_474), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_98), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_99), .B(n_378), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_101), .A2(n_213), .B1(n_289), .B2(n_294), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_102), .A2(n_178), .B1(n_295), .B2(n_696), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_103), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_105), .A2(n_136), .B1(n_618), .B2(n_631), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g641 ( .A1(n_106), .A2(n_137), .B1(n_173), .B2(n_304), .C1(n_342), .C2(n_490), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_107), .A2(n_190), .B1(n_394), .B2(n_467), .Y(n_466) );
AOI22x1_ASAP7_75t_L g501 ( .A1(n_108), .A2(n_502), .B1(n_539), .B2(n_540), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_108), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_111), .A2(n_145), .B1(n_403), .B2(n_404), .Y(n_402) );
INVx2_ASAP7_75t_L g230 ( .A(n_112), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_113), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_116), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_117), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_119), .A2(n_192), .B1(n_331), .B2(n_387), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_120), .B(n_256), .Y(n_705) );
AND2x6_ASAP7_75t_L g225 ( .A(n_121), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_121), .Y(n_650) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_122), .A2(n_184), .B1(n_244), .B2(n_249), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_123), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_125), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_126), .A2(n_185), .B1(n_354), .B2(n_355), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g374 ( .A1(n_127), .A2(n_161), .B1(n_375), .B2(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g498 ( .A(n_128), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_129), .A2(n_183), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_133), .A2(n_219), .B1(n_399), .B2(n_400), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_134), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_135), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_139), .A2(n_212), .B1(n_363), .B2(n_465), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_140), .A2(n_177), .B1(n_260), .B2(n_266), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_141), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_142), .A2(n_175), .B1(n_394), .B2(n_396), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_143), .A2(n_660), .B1(n_661), .B2(n_681), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_143), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_147), .A2(n_180), .B1(n_280), .B2(n_416), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_148), .B(n_255), .Y(n_488) );
AO22x2_ASAP7_75t_L g243 ( .A1(n_149), .A2(n_193), .B1(n_244), .B2(n_245), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_150), .A2(n_199), .B1(n_363), .B2(n_566), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_151), .B(n_381), .Y(n_611) );
XOR2x2_ASAP7_75t_L g625 ( .A(n_152), .B(n_626), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_153), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_158), .A2(n_160), .B1(n_299), .B2(n_416), .Y(n_675) );
INVx1_ASAP7_75t_L g554 ( .A(n_163), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_164), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_165), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_167), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_168), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_170), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_174), .A2(n_217), .B1(n_266), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_176), .A2(n_209), .B1(n_414), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_181), .A2(n_216), .B1(n_394), .B2(n_396), .Y(n_581) );
XOR2x2_ASAP7_75t_L g369 ( .A(n_182), .B(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_184), .B(n_655), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_186), .A2(n_223), .B(n_231), .C(n_658), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_189), .A2(n_196), .B1(n_639), .B2(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g653 ( .A(n_193), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_194), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_195), .A2(n_218), .B1(n_381), .B2(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g373 ( .A(n_197), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_198), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_200), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_202), .Y(n_608) );
INVx1_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
INVx1_ASAP7_75t_L g246 ( .A(n_203), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_208), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_210), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_211), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_214), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_220), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_221), .B(n_420), .Y(n_612) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_226), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_227), .A2(n_648), .B(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_570), .B1(n_571), .B2(n_644), .C(n_645), .Y(n_231) );
INVx1_ASAP7_75t_L g644 ( .A(n_232), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_408), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_314), .B1(n_315), .B2(n_407), .Y(n_233) );
INVx1_ASAP7_75t_L g407 ( .A(n_234), .Y(n_407) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND4xp75_ASAP7_75t_L g236 ( .A(n_237), .B(n_269), .C(n_287), .D(n_302), .Y(n_236) );
AND2x2_ASAP7_75t_SL g237 ( .A(n_238), .B(n_258), .Y(n_237) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g384 ( .A(n_240), .Y(n_384) );
INVx5_ASAP7_75t_L g420 ( .A(n_240), .Y(n_420) );
INVx2_ASAP7_75t_L g670 ( .A(n_240), .Y(n_670) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_250), .Y(n_241) );
AND2x6_ASAP7_75t_L g256 ( .A(n_242), .B(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g282 ( .A(n_242), .B(n_275), .Y(n_282) );
INVx1_ASAP7_75t_L g324 ( .A(n_242), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_242), .B(n_257), .Y(n_328) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVx1_ASAP7_75t_L g262 ( .A(n_243), .Y(n_262) );
INVx1_ASAP7_75t_L g274 ( .A(n_243), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_243), .B(n_248), .Y(n_278) );
INVx1_ASAP7_75t_L g293 ( .A(n_243), .Y(n_293) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g249 ( .A(n_246), .Y(n_249) );
AND2x2_ASAP7_75t_L g292 ( .A(n_247), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g264 ( .A(n_248), .B(n_253), .Y(n_264) );
AND2x2_ASAP7_75t_L g273 ( .A(n_248), .B(n_274), .Y(n_273) );
AND2x6_ASAP7_75t_L g291 ( .A(n_250), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g323 ( .A(n_251), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g257 ( .A(n_252), .B(n_254), .Y(n_257) );
AND2x2_ASAP7_75t_L g275 ( .A(n_252), .B(n_263), .Y(n_275) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g305 ( .A(n_253), .B(n_254), .Y(n_305) );
INVx2_ASAP7_75t_L g263 ( .A(n_254), .Y(n_263) );
INVx1_ASAP7_75t_L g268 ( .A(n_254), .Y(n_268) );
BUFx4f_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_SL g382 ( .A(n_256), .Y(n_382) );
AND2x4_ASAP7_75t_L g295 ( .A(n_257), .B(n_292), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_257), .B(n_273), .Y(n_301) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_259), .Y(n_448) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_260), .Y(n_335) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_260), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g490 ( .A(n_260), .Y(n_490) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g310 ( .A(n_262), .Y(n_310) );
INVx1_ASAP7_75t_L g417 ( .A(n_263), .Y(n_417) );
AND2x4_ASAP7_75t_L g266 ( .A(n_264), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g309 ( .A(n_264), .B(n_310), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_264), .B(n_417), .Y(n_454) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
BUFx2_ASAP7_75t_L g386 ( .A(n_266), .Y(n_386) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x6_ASAP7_75t_L g277 ( .A(n_268), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_279), .Y(n_269) );
INVx1_ASAP7_75t_L g401 ( .A(n_271), .Y(n_401) );
BUFx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx3_ASAP7_75t_L g363 ( .A(n_272), .Y(n_363) );
BUFx3_ASAP7_75t_L g559 ( .A(n_272), .Y(n_559) );
BUFx3_ASAP7_75t_L g621 ( .A(n_272), .Y(n_621) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_273), .B(n_275), .Y(n_519) );
INVx1_ASAP7_75t_L g313 ( .A(n_274), .Y(n_313) );
AND2x4_ASAP7_75t_L g285 ( .A(n_275), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g298 ( .A(n_275), .B(n_292), .Y(n_298) );
BUFx2_ASAP7_75t_L g396 ( .A(n_276), .Y(n_396) );
BUFx2_ASAP7_75t_L g467 ( .A(n_276), .Y(n_467) );
BUFx2_ASAP7_75t_L g631 ( .A(n_276), .Y(n_631) );
INVx6_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_SL g355 ( .A(n_277), .Y(n_355) );
INVx1_ASAP7_75t_L g286 ( .A(n_278), .Y(n_286) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_282), .Y(n_351) );
BUFx3_ASAP7_75t_L g470 ( .A(n_282), .Y(n_470) );
BUFx3_ASAP7_75t_L g509 ( .A(n_282), .Y(n_509) );
BUFx3_ASAP7_75t_L g565 ( .A(n_282), .Y(n_565) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx3_ASAP7_75t_L g364 ( .A(n_285), .Y(n_364) );
BUFx2_ASAP7_75t_SL g404 ( .A(n_285), .Y(n_404) );
BUFx3_ASAP7_75t_L g465 ( .A(n_285), .Y(n_465) );
BUFx2_ASAP7_75t_L g566 ( .A(n_285), .Y(n_566) );
BUFx2_ASAP7_75t_SL g622 ( .A(n_285), .Y(n_622) );
AND2x2_ASAP7_75t_L g416 ( .A(n_286), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_296), .Y(n_287) );
INVx4_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g464 ( .A(n_290), .Y(n_464) );
INVx2_ASAP7_75t_SL g624 ( .A(n_290), .Y(n_624) );
INVx11_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx11_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
AND2x6_ASAP7_75t_L g304 ( .A(n_292), .B(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx6_ASAP7_75t_L g360 ( .A(n_295), .Y(n_360) );
BUFx3_ASAP7_75t_L g414 ( .A(n_295), .Y(n_414) );
BUFx3_ASAP7_75t_L g358 ( .A(n_297), .Y(n_358) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_297), .Y(n_399) );
INVx3_ASAP7_75t_L g505 ( .A(n_297), .Y(n_505) );
BUFx3_ASAP7_75t_L g586 ( .A(n_297), .Y(n_586) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_SL g558 ( .A(n_298), .Y(n_558) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_298), .Y(n_616) );
INVx2_ASAP7_75t_L g680 ( .A(n_298), .Y(n_680) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
INVx5_ASAP7_75t_L g395 ( .A(n_300), .Y(n_395) );
INVx4_ASAP7_75t_L g696 ( .A(n_300), .Y(n_696) );
INVx8_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g530 ( .A(n_303), .Y(n_530) );
INVx2_ASAP7_75t_SL g607 ( .A(n_303), .Y(n_607) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx4_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
BUFx3_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx2_ASAP7_75t_L g482 ( .A(n_304), .Y(n_482) );
AND2x4_ASAP7_75t_L g312 ( .A(n_305), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g459 ( .A(n_305), .Y(n_459) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx4f_ASAP7_75t_SL g342 ( .A(n_308), .Y(n_342) );
BUFx12f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_309), .Y(n_378) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_309), .Y(n_485) );
BUFx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_SL g387 ( .A(n_312), .Y(n_387) );
BUFx3_ASAP7_75t_L g427 ( .A(n_312), .Y(n_427) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_312), .Y(n_702) );
INVx1_ASAP7_75t_L g460 ( .A(n_313), .Y(n_460) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_367), .B1(n_405), .B2(n_406), .Y(n_315) );
INVx1_ASAP7_75t_L g405 ( .A(n_316), .Y(n_405) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_344), .Y(n_318) );
NOR2xp33_ASAP7_75t_SL g319 ( .A(n_320), .B(n_333), .Y(n_319) );
OAI221xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_325), .B1(n_326), .B2(n_329), .C(n_330), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_321), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_321), .A2(n_526), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g440 ( .A(n_322), .Y(n_440) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g546 ( .A(n_323), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_326), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_544) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g526 ( .A(n_327), .Y(n_526) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g444 ( .A(n_328), .Y(n_444) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI222xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B1(n_337), .B2(n_340), .C1(n_341), .C2(n_343), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_337), .A2(n_373), .B(n_374), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g445 ( .A1(n_337), .A2(n_446), .B1(n_447), .B2(n_449), .C(n_450), .Y(n_445) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_339), .A2(n_700), .B(n_701), .Y(n_699) );
OAI222xp33_ASAP7_75t_L g527 ( .A1(n_341), .A2(n_528), .B1(n_529), .B2(n_530), .C1(n_531), .C2(n_532), .Y(n_527) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_356), .Y(n_344) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_349), .B1(n_350), .B2(n_352), .C(n_353), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g582 ( .A1(n_346), .A2(n_507), .B1(n_583), .B2(n_584), .C(n_585), .Y(n_582) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g392 ( .A(n_348), .Y(n_392) );
INVx2_ASAP7_75t_L g512 ( .A(n_348), .Y(n_512) );
INVx1_ASAP7_75t_L g639 ( .A(n_348), .Y(n_639) );
INVx4_ASAP7_75t_L g629 ( .A(n_350), .Y(n_629) );
INVx4_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp33_ASAP7_75t_SL g356 ( .A(n_357), .B(n_361), .Y(n_356) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
INVx3_ASAP7_75t_L g563 ( .A(n_360), .Y(n_563) );
INVx2_ASAP7_75t_L g640 ( .A(n_360), .Y(n_640) );
BUFx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_364), .Y(n_513) );
INVx2_ASAP7_75t_L g579 ( .A(n_364), .Y(n_579) );
INVx1_ASAP7_75t_L g406 ( .A(n_367), .Y(n_406) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND3x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_388), .C(n_397), .Y(n_370) );
NOR2x1_ASAP7_75t_SL g371 ( .A(n_372), .B(n_379), .Y(n_371) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .C(n_385), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_395), .Y(n_618) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g515 ( .A(n_403), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_429), .B2(n_569), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
XOR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_428), .Y(n_410) );
NAND4xp75_ASAP7_75t_L g411 ( .A(n_412), .B(n_418), .C(n_422), .D(n_425), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx3_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_419), .B(n_421), .Y(n_418) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_420), .Y(n_634) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx3_ASAP7_75t_L g550 ( .A(n_426), .Y(n_550) );
INVx1_ASAP7_75t_L g569 ( .A(n_429), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B1(n_541), .B2(n_568), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
XNOR2xp5_ASAP7_75t_SL g431 ( .A(n_432), .B(n_501), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_475), .B2(n_499), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_461), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_445), .C(n_451), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g591 ( .A1(n_447), .A2(n_530), .B1(n_592), .B2(n_593), .C1(n_594), .C2(n_596), .Y(n_591) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_455), .B2(n_456), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_453), .A2(n_458), .B1(n_553), .B2(n_554), .Y(n_552) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g536 ( .A(n_454), .Y(n_536) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g538 ( .A(n_457), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_468), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g500 ( .A(n_478), .Y(n_500) );
XOR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_498), .Y(n_478) );
NAND2x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_491), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_486), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_483), .B(n_484), .Y(n_481) );
BUFx3_ASAP7_75t_L g595 ( .A(n_485), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .C(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g528 ( .A(n_490), .Y(n_528) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g540 ( .A(n_502), .Y(n_540) );
AND2x2_ASAP7_75t_SL g502 ( .A(n_503), .B(n_522), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
OAI221xp5_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_506), .B1(n_507), .B2(n_510), .C(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI221xp5_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_516), .B1(n_517), .B2(n_520), .C(n_521), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g577 ( .A(n_518), .Y(n_577) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .C(n_533), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_537), .B2(n_538), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_535), .A2(n_538), .B1(n_598), .B2(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g568 ( .A(n_541), .Y(n_568) );
XOR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_567), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_555), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .C(n_552), .Y(n_543) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B(n_551), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_550), .A2(n_665), .B(n_666), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_561), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_602), .B1(n_642), .B2(n_643), .Y(n_571) );
INVx1_ASAP7_75t_L g642 ( .A(n_572), .Y(n_642) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_587), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_582), .Y(n_575) );
OAI221xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_578), .B1(n_579), .B2(n_580), .C(n_581), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .C(n_597), .Y(n_587) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g643 ( .A(n_602), .Y(n_643) );
XNOR2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_625), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_614), .C(n_619), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_610), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B(n_609), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .C(n_613), .Y(n_610) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g626 ( .A(n_627), .B(n_632), .C(n_636), .D(n_641), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AND2x2_ASAP7_75t_SL g632 ( .A(n_633), .B(n_635), .Y(n_632) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
OR2x2_ASAP7_75t_SL g712 ( .A(n_647), .B(n_652), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_648), .Y(n_683) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_649), .B(n_687), .Y(n_690) );
CKINVDCx16_ASAP7_75t_R g687 ( .A(n_650), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
OAI322xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_682), .A3(n_684), .B1(n_688), .B2(n_691), .C1(n_692), .C2(n_710), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_672), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .C(n_671), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_689), .Y(n_688) );
XOR2x2_ASAP7_75t_L g692 ( .A(n_691), .B(n_693), .Y(n_692) );
NAND3x1_ASAP7_75t_SL g693 ( .A(n_694), .B(n_698), .C(n_707), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_703), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .C(n_706), .Y(n_703) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
endmodule