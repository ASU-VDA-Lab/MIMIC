module real_jpeg_14805_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_342, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_342;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_3),
.Y(n_340)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_5),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_5),
.A2(n_67),
.B1(n_69),
.B2(n_135),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_135),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_5),
.A2(n_57),
.B1(n_62),
.B2(n_135),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_6),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_184),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_6),
.A2(n_67),
.B1(n_69),
.B2(n_184),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_6),
.A2(n_57),
.B1(n_62),
.B2(n_184),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_39),
.B1(n_57),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_39),
.B1(n_67),
.B2(n_69),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_7),
.A2(n_29),
.B1(n_32),
.B2(n_39),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_8),
.A2(n_29),
.B1(n_32),
.B2(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_9),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_9),
.A2(n_29),
.B1(n_32),
.B2(n_171),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_9),
.A2(n_67),
.B1(n_69),
.B2(n_171),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_9),
.A2(n_57),
.B1(n_62),
.B2(n_171),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_10),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_79),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_67),
.B1(n_69),
.B2(n_79),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_57),
.B1(n_62),
.B2(n_79),
.Y(n_204)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_12),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_29),
.B1(n_32),
.B2(n_81),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_12),
.A2(n_67),
.B1(n_69),
.B2(n_81),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_57),
.B1(n_62),
.B2(n_81),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_16),
.A2(n_42),
.B1(n_67),
.B2(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_16),
.A2(n_29),
.B1(n_32),
.B2(n_42),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_16),
.A2(n_42),
.B1(n_57),
.B2(n_62),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_17),
.A2(n_29),
.B1(n_32),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_17),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_17),
.A2(n_67),
.B1(n_69),
.B2(n_87),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_17),
.A2(n_57),
.B1(n_62),
.B2(n_87),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_18),
.B(n_37),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_18),
.A2(n_34),
.B(n_210),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_18),
.A2(n_67),
.B1(n_69),
.B2(n_201),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_18),
.A2(n_69),
.B(n_72),
.C(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_18),
.B(n_94),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_18),
.B(n_60),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_18),
.B(n_76),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_18),
.A2(n_32),
.B(n_88),
.C(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_339),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_19),
.B(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_37),
.B(n_38),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_26),
.A2(n_37),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_26),
.A2(n_37),
.B1(n_41),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_27),
.A2(n_28),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_27),
.A2(n_28),
.B1(n_80),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_28),
.B1(n_78),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_27),
.A2(n_28),
.B1(n_100),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_27),
.A2(n_28),
.B1(n_134),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_27),
.A2(n_28),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_29),
.A2(n_32),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_29),
.B(n_201),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_29),
.A2(n_31),
.A3(n_34),
.B1(n_211),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_30),
.B(n_32),
.Y(n_225)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_32),
.A2(n_67),
.A3(n_90),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_35),
.B(n_201),
.Y(n_211)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_40),
.B(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_44),
.B(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_334),
.B(n_336),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_322),
.B(n_333),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_149),
.B(n_319),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_136),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_111),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_50),
.B(n_111),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_82),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_51),
.B(n_97),
.C(n_109),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B(n_77),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_53),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_55),
.B1(n_77),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_61),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_56),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_56),
.A2(n_60),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_56),
.A2(n_60),
.B1(n_190),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_56),
.A2(n_60),
.B1(n_162),
.B2(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_56),
.A2(n_60),
.B1(n_204),
.B2(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_56),
.A2(n_60),
.B1(n_201),
.B2(n_257),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_56),
.A2(n_60),
.B1(n_250),
.B2(n_257),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_57),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_62),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_57),
.B(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_125),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_59),
.A2(n_160),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_62),
.A2(n_73),
.B(n_201),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_70),
.B1(n_76),
.B2(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_69),
.B1(n_90),
.B2(n_91),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_69),
.B(n_91),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_75),
.B1(n_76),
.B2(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_76),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_70),
.A2(n_76),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_70),
.A2(n_76),
.B1(n_165),
.B2(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_70),
.A2(n_76),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_70),
.A2(n_76),
.B1(n_236),
.B2(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_74),
.A2(n_129),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_74),
.A2(n_166),
.B1(n_194),
.B2(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_77),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_97),
.B1(n_109),
.B2(n_110),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_84),
.B(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_92),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_88),
.A2(n_94),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_88),
.A2(n_94),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_88),
.A2(n_94),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_92),
.A2(n_107),
.B1(n_131),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_92),
.A2(n_131),
.B1(n_132),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_92),
.A2(n_131),
.B1(n_186),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_92),
.A2(n_183),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_99),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_103),
.C(n_105),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_99),
.B(n_139),
.C(n_142),
.Y(n_323)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_108),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_103),
.B(n_145),
.C(n_147),
.Y(n_332)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_119),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.C(n_133),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_121),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_304)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_136),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_137),
.B(n_138),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_146),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_148),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_174),
.B(n_318),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_172),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_172),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_152),
.B(n_155),
.Y(n_316)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_156),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.C(n_169),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_157),
.A2(n_158),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_159),
.B(n_163),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_167),
.B(n_169),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_168),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_170),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_313),
.B(n_317),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_300),
.B1(n_311),
.B2(n_312),
.C(n_342),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_285),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_228),
.B(n_284),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_205),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_179),
.B(n_205),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_192),
.C(n_196),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_180),
.B(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_188),
.C(n_189),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_192),
.A2(n_196),
.B1(n_197),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_198),
.A2(n_199),
.B1(n_203),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_219),
.B2(n_227),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_206),
.B(n_220),
.C(n_226),
.Y(n_286)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_208),
.B(n_214),
.C(n_218),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_215),
.Y(n_294)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_221),
.B(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_278),
.B(n_283),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_266),
.B(n_277),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_246),
.B(n_265),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_232),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_242),
.C(n_244),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_254),
.B(n_264),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_252),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_260),
.B(n_263),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_268),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_287),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_296),
.C(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_302),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_308),
.B2(n_309),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_309),
.C(n_310),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_330),
.C(n_332),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_335),
.Y(n_338)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule