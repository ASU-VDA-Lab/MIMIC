module real_jpeg_19536_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_77),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_3),
.A2(n_66),
.B1(n_67),
.B2(n_84),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_84),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_84),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_82),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_4),
.A2(n_14),
.B(n_29),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_78),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_4),
.A2(n_26),
.B1(n_116),
.B2(n_151),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_4),
.B(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_66),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_4),
.A2(n_66),
.B(n_177),
.Y(n_181)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_5),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_58),
.B1(n_66),
.B2(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_72),
.B1(n_77),
.B2(n_85),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_72),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_74),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_91)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_80),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_39),
.B(n_42),
.C(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_106),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_52),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_26),
.A2(n_32),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_26),
.A2(n_31),
.B1(n_135),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_26),
.A2(n_138),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_27),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_27),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_27),
.A2(n_35),
.B(n_169),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_28),
.B(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_30),
.B(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_39),
.A2(n_50),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_39),
.B(n_78),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_39),
.A2(n_50),
.B1(n_146),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_39),
.A2(n_50),
.B1(n_166),
.B2(n_184),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_40),
.A2(n_43),
.B(n_78),
.C(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_43),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_42),
.A2(n_67),
.A3(n_70),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_43),
.B(n_64),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_50),
.A2(n_184),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.C(n_75),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_57),
.B(n_60),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_63),
.A2(n_69),
.B1(n_122),
.B2(n_181),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_66),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_80),
.Y(n_89)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_76),
.B1(n_81),
.B2(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_71),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.CON(n_76),
.SN(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_80),
.Y(n_81)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_78),
.B(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_112),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_108),
.B(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_120),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_120),
.B(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_202),
.B(n_206),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_189),
.B(n_201),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_171),
.B(n_188),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_158),
.B(n_170),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_147),
.B(n_157),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_143),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_152),
.B(n_156),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_160),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_173),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_179),
.B1(n_186),
.B2(n_187),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_185),
.C(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_191),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_198),
.C(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);


endmodule