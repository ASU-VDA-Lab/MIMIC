module fake_netlist_1_12396_n_695 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_695);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_695;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_584;
wire n_121;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_29), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_85), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_25), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_36), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_61), .Y(n_98) );
OR2x2_ASAP7_75t_L g99 ( .A(n_43), .B(n_75), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_19), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_68), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_26), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_16), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_7), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_84), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_20), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_22), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_83), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_69), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_10), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_49), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_62), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_77), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_47), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_10), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_51), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_55), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_30), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_48), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_67), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_9), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_17), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_72), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_9), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_11), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_81), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_54), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_34), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_122), .B(n_0), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_102), .B(n_0), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_102), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_93), .B(n_1), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_105), .B(n_1), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_95), .B(n_2), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_137), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_103), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_106), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_97), .B(n_2), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_101), .Y(n_156) );
AO22x2_ASAP7_75t_L g157 ( .A1(n_139), .A2(n_146), .B1(n_155), .B2(n_148), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
INVx5_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_148), .B(n_118), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
INVx5_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_149), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_150), .B(n_125), .C(n_128), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_145), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_150), .B(n_96), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_146), .B(n_151), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_156), .B(n_98), .Y(n_181) );
INVx5_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_175), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g185 ( .A(n_177), .B(n_94), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_175), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_157), .A2(n_155), .B1(n_151), .B2(n_145), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_177), .B(n_138), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_169), .B(n_152), .Y(n_189) );
NOR2x2_ASAP7_75t_L g190 ( .A(n_169), .B(n_153), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_181), .B(n_153), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_174), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
NOR2x2_ASAP7_75t_L g194 ( .A(n_174), .B(n_154), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_147), .B(n_133), .C(n_129), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_177), .B(n_154), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_157), .A2(n_113), .B1(n_107), .B2(n_134), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_177), .B(n_98), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_175), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_160), .B(n_101), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_176), .B(n_110), .Y(n_201) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_182), .B(n_124), .Y(n_202) );
AOI221xp5_ASAP7_75t_L g203 ( .A1(n_157), .A2(n_104), .B1(n_108), .B2(n_130), .C(n_116), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_164), .B(n_104), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_182), .B(n_110), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_182), .B(n_119), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_164), .B(n_144), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_182), .B(n_119), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_159), .A2(n_108), .B1(n_116), .B2(n_130), .Y(n_210) );
NOR2xp67_ASAP7_75t_L g211 ( .A(n_182), .B(n_99), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_159), .A2(n_123), .B1(n_131), .B2(n_127), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_167), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_159), .A2(n_123), .B1(n_135), .B2(n_126), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_159), .B(n_120), .Y(n_215) );
AND2x6_ASAP7_75t_SL g216 ( .A(n_168), .B(n_3), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_200), .A2(n_168), .B(n_178), .C(n_171), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_202), .B(n_182), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_203), .A2(n_182), .B1(n_173), .B2(n_163), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_188), .A2(n_163), .B(n_159), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_213), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_213), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_187), .A2(n_163), .B1(n_159), .B2(n_173), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_200), .B(n_159), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_193), .B(n_163), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_184), .A2(n_163), .B1(n_178), .B2(n_172), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_202), .B(n_163), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
AO21x1_ASAP7_75t_L g229 ( .A1(n_184), .A2(n_158), .B(n_165), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_185), .B(n_120), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_204), .B(n_163), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_204), .B(n_171), .Y(n_232) );
NOR2x1p5_ASAP7_75t_SL g233 ( .A(n_183), .B(n_161), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_193), .B(n_189), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_192), .Y(n_235) );
NAND3xp33_ASAP7_75t_L g236 ( .A(n_203), .B(n_172), .C(n_175), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_189), .B(n_180), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_196), .A2(n_158), .B(n_165), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_196), .B(n_180), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g240 ( .A1(n_209), .A2(n_167), .B(n_179), .C(n_170), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_208), .A2(n_179), .B(n_170), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_198), .B(n_180), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_185), .B(n_180), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_212), .B(n_167), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_197), .A2(n_179), .B1(n_170), .B2(n_175), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_208), .A2(n_162), .B(n_161), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_235), .B(n_201), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_241), .A2(n_215), .B(n_211), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_218), .A2(n_161), .B(n_162), .Y(n_250) );
AOI21xp5_ASAP7_75t_SL g251 ( .A1(n_221), .A2(n_211), .B(n_215), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_238), .A2(n_207), .B(n_206), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_222), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_236), .A2(n_207), .B(n_191), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_240), .A2(n_205), .B(n_186), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_234), .B(n_210), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_229), .A2(n_183), .B(n_186), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_228), .A2(n_186), .B(n_199), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_199), .B(n_162), .Y(n_260) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_222), .A2(n_199), .A3(n_175), .B(n_194), .Y(n_261) );
AO31x2_ASAP7_75t_L g262 ( .A1(n_223), .A2(n_195), .A3(n_216), .B(n_190), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_225), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_234), .B(n_195), .Y(n_264) );
NOR4xp25_ASAP7_75t_L g265 ( .A(n_217), .B(n_216), .C(n_214), .D(n_114), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_232), .A2(n_136), .B(n_135), .C(n_126), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_227), .A2(n_50), .B(n_92), .C(n_91), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_225), .Y(n_268) );
AO22x2_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_239), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_253), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_270), .B(n_224), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_258), .B(n_226), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_269), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_249), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_250), .A2(n_246), .B(n_242), .Y(n_278) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_250), .A2(n_231), .A3(n_228), .B(n_220), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_257), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_248), .A2(n_245), .B(n_226), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_269), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_268), .B(n_243), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_249), .Y(n_284) );
INVx8_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_260), .A2(n_245), .B(n_244), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_255), .A2(n_230), .B(n_244), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_268), .B(n_219), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_265), .B(n_235), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
AO31x2_ASAP7_75t_L g291 ( .A1(n_264), .A2(n_233), .A3(n_5), .B(n_6), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_275), .B(n_261), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_289), .A2(n_256), .B1(n_268), .B2(n_263), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_291), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_291), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_287), .A2(n_254), .B(n_252), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_285), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_291), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_275), .B(n_261), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_286), .A2(n_256), .B(n_266), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_274), .B(n_263), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_291), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_271), .Y(n_307) );
AO21x1_ASAP7_75t_L g308 ( .A1(n_282), .A2(n_260), .B(n_259), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_291), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_272), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_291), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_282), .B(n_261), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_274), .B(n_263), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_272), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_272), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_272), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_294), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_292), .B(n_290), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_290), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_280), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_316), .B(n_272), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_301), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_296), .B(n_280), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_300), .B(n_291), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_317), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_300), .B(n_286), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_301), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_305), .B(n_286), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_305), .B(n_281), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_302), .A2(n_289), .B1(n_288), .B2(n_283), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_299), .B(n_247), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_309), .B(n_281), .Y(n_339) );
INVx5_ASAP7_75t_L g340 ( .A(n_317), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_295), .Y(n_341) );
AND2x4_ASAP7_75t_SL g342 ( .A(n_310), .B(n_283), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_309), .B(n_281), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_312), .B(n_281), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_312), .B(n_284), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_306), .B(n_279), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_311), .B(n_281), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_311), .B(n_279), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_316), .B(n_279), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_297), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_298), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_297), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_310), .B(n_279), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_302), .B(n_279), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_297), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_298), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_324), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_325), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_322), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_319), .B(n_307), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_358), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_321), .B(n_307), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_319), .B(n_315), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_361), .A2(n_288), .B1(n_283), .B2(n_293), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_358), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_360), .B(n_297), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_319), .B(n_315), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_320), .B(n_318), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_321), .B(n_318), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_321), .B(n_308), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_361), .B(n_308), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_361), .B(n_304), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_334), .B(n_304), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_338), .B(n_317), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_334), .B(n_314), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_333), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_360), .B(n_314), .Y(n_393) );
AND2x4_ASAP7_75t_SL g394 ( .A(n_360), .B(n_276), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_346), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_326), .B(n_261), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_326), .B(n_276), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_338), .B(n_4), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_334), .B(n_279), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_331), .B(n_279), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_340), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_331), .B(n_262), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_351), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_336), .B(n_284), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_339), .B(n_288), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_339), .B(n_287), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_336), .B(n_284), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_339), .B(n_278), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_329), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_345), .B(n_278), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_337), .B(n_262), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_340), .B(n_284), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_329), .Y(n_414) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_360), .B(n_284), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_337), .B(n_262), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_333), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_345), .B(n_262), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_352), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_345), .B(n_6), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_360), .B(n_233), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_347), .B(n_7), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_347), .B(n_273), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_347), .B(n_352), .Y(n_424) );
AND2x2_ASAP7_75t_SL g425 ( .A(n_342), .B(n_273), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_333), .Y(n_426) );
AOI21xp5_ASAP7_75t_SL g427 ( .A1(n_348), .A2(n_266), .B(n_136), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_328), .B(n_8), .Y(n_428) );
AND2x4_ASAP7_75t_SL g429 ( .A(n_355), .B(n_285), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_370), .B(n_355), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_371), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_379), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_420), .B(n_328), .Y(n_433) );
AND2x4_ASAP7_75t_SL g434 ( .A(n_370), .B(n_355), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_371), .B(n_341), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_379), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_376), .B(n_342), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_374), .B(n_341), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_420), .B(n_328), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_376), .B(n_342), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_381), .B(n_355), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_381), .B(n_341), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_425), .A2(n_335), .B1(n_355), .B2(n_340), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_389), .B(n_354), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_400), .B(n_354), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_422), .B(n_335), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_400), .B(n_354), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_414), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_424), .B(n_344), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_373), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_385), .B(n_353), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_425), .B(n_340), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_365), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_389), .B(n_330), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_365), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_424), .B(n_344), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_368), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_370), .B(n_349), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_368), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_391), .B(n_330), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_391), .B(n_330), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_422), .B(n_332), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_384), .B(n_344), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_428), .B(n_332), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_384), .B(n_350), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_399), .B(n_340), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_370), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_409), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_387), .B(n_332), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_428), .B(n_353), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_377), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_369), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_387), .B(n_353), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_369), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_406), .B(n_323), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_406), .B(n_323), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_372), .B(n_350), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_372), .B(n_350), .Y(n_479) );
OR2x2_ASAP7_75t_SL g480 ( .A(n_418), .B(n_340), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_375), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_375), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_382), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_382), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_403), .B(n_349), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_364), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_388), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_429), .B(n_323), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_412), .B(n_349), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_423), .B(n_327), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_364), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_388), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_364), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_429), .B(n_327), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_429), .B(n_327), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_385), .B(n_349), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_377), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_398), .B(n_349), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_395), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_395), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_386), .B(n_359), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_398), .B(n_325), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_416), .B(n_356), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_366), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_386), .B(n_359), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_390), .B(n_340), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_367), .B(n_359), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_377), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_409), .B(n_359), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_383), .B(n_356), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_383), .B(n_359), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_425), .B(n_348), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_451), .B(n_402), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_434), .B(n_394), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_446), .B(n_394), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_452), .B(n_411), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_452), .B(n_411), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_446), .B(n_401), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_453), .A2(n_378), .B1(n_402), .B2(n_394), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_448), .B(n_401), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_448), .B(n_393), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_485), .B(n_393), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_473), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_454), .B(n_407), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_442), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_445), .B(n_393), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_442), .B(n_427), .C(n_362), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_489), .B(n_393), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_501), .B(n_407), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_474), .B(n_415), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_481), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_482), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_501), .B(n_396), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_443), .B(n_397), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_464), .B(n_405), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_472), .B(n_413), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_456), .B(n_396), .Y(n_540) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_453), .A2(n_367), .B1(n_408), .B2(n_405), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_496), .B(n_415), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_466), .B(n_408), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_468), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_435), .B(n_404), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_483), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_496), .B(n_415), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_431), .B(n_404), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_449), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_432), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_468), .B(n_367), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_508), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_449), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_492), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_441), .B(n_380), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_438), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_467), .B(n_427), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_434), .B(n_367), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_505), .B(n_419), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_455), .B(n_380), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_450), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_493), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_505), .B(n_419), .Y(n_569) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_506), .B(n_421), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_457), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_478), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_486), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_506), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_479), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_430), .B(n_421), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_498), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_469), .B(n_421), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_469), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_444), .A2(n_421), .B1(n_426), .B2(n_366), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_380), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_436), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_436), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_511), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_461), .B(n_380), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_503), .B(n_357), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_582), .B(n_470), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_562), .A2(n_574), .B1(n_521), .B2(n_570), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_566), .B(n_509), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_530), .A2(n_430), .B(n_467), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_551), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_572), .B(n_462), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_586), .B(n_509), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_564), .B(n_497), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_554), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g597 ( .A1(n_521), .A2(n_447), .B1(n_512), .B2(n_433), .C1(n_439), .C2(n_463), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_530), .A2(n_430), .B(n_459), .Y(n_598) );
NAND3xp33_ASAP7_75t_SL g599 ( .A(n_554), .B(n_512), .C(n_502), .Y(n_599) );
AOI32xp33_ASAP7_75t_L g600 ( .A1(n_516), .A2(n_495), .A3(n_494), .B1(n_488), .B2(n_440), .Y(n_600) );
AO221x1_ASAP7_75t_L g601 ( .A1(n_541), .A2(n_480), .B1(n_472), .B2(n_497), .C(n_459), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_579), .B(n_477), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_583), .B(n_471), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_550), .A2(n_465), .B1(n_459), .B2(n_507), .C1(n_437), .C2(n_504), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_556), .B(n_507), .C(n_362), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_513), .A2(n_507), .B1(n_504), .B2(n_491), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_527), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_573), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_575), .B(n_491), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_536), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_584), .B(n_357), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_559), .B(n_357), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_528), .B(n_362), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_580), .B(n_267), .C(n_121), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_362), .Y(n_617) );
AOI32xp33_ASAP7_75t_L g618 ( .A1(n_515), .A2(n_426), .A3(n_366), .B1(n_392), .B2(n_417), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
AOI322xp5_ASAP7_75t_L g620 ( .A1(n_517), .A2(n_426), .A3(n_417), .B1(n_392), .B2(n_363), .C1(n_362), .C2(n_285), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_544), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_576), .A2(n_362), .B1(n_363), .B2(n_267), .C(n_121), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_515), .A2(n_362), .B1(n_285), .B2(n_112), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_578), .A2(n_285), .B1(n_166), .B2(n_12), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_519), .B(n_8), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_563), .B(n_11), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_523), .A2(n_251), .B1(n_13), .B2(n_14), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_563), .A2(n_14), .B1(n_15), .B2(n_17), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_569), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_553), .A2(n_166), .B(n_18), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_544), .B(n_15), .C(n_18), .D(n_20), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_514), .Y(n_632) );
AOI21xp33_ASAP7_75t_SL g633 ( .A1(n_539), .A2(n_21), .B(n_22), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_533), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_589), .A2(n_552), .B1(n_539), .B2(n_540), .C(n_532), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_631), .A2(n_561), .B(n_532), .C(n_518), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_596), .B(n_517), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_603), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_601), .A2(n_587), .B(n_548), .Y(n_639) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_599), .A2(n_518), .A3(n_577), .B1(n_526), .B2(n_585), .C1(n_571), .C2(n_567), .Y(n_640) );
AOI222xp33_ASAP7_75t_L g641 ( .A1(n_628), .A2(n_587), .B1(n_560), .B2(n_558), .C1(n_557), .C2(n_555), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_628), .A2(n_535), .B(n_549), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_597), .B(n_520), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_597), .A2(n_547), .B1(n_524), .B2(n_531), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_605), .A2(n_525), .B1(n_529), .B2(n_546), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_626), .A2(n_522), .B1(n_581), .B2(n_534), .C(n_545), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_605), .B(n_537), .C(n_538), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_626), .A2(n_543), .B1(n_23), .B2(n_21), .C(n_166), .Y(n_648) );
CKINVDCx6p67_ASAP7_75t_R g649 ( .A(n_625), .Y(n_649) );
AOI322xp5_ASAP7_75t_L g650 ( .A1(n_593), .A2(n_23), .A3(n_166), .B1(n_27), .B2(n_28), .C1(n_32), .C2(n_33), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_590), .B(n_24), .Y(n_651) );
AOI31xp33_ASAP7_75t_L g652 ( .A1(n_623), .A2(n_35), .A3(n_37), .B(n_38), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_618), .A2(n_166), .B1(n_41), .B2(n_42), .C(n_44), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_612), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_610), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g656 ( .A1(n_600), .A2(n_40), .B(n_45), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_598), .A2(n_46), .B1(n_52), .B2(n_53), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_591), .A2(n_56), .B(n_57), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_619), .A2(n_59), .B1(n_60), .B2(n_64), .C(n_65), .Y(n_659) );
AOI221x1_ASAP7_75t_L g660 ( .A1(n_631), .A2(n_66), .B1(n_70), .B2(n_71), .C(n_73), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_633), .A2(n_76), .B(n_78), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_620), .A2(n_80), .B(n_86), .C(n_87), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_629), .B(n_88), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g664 ( .A(n_627), .B(n_89), .C(n_632), .D(n_624), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_630), .A2(n_595), .B(n_634), .C(n_616), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_627), .A2(n_604), .B1(n_602), .B2(n_588), .C1(n_611), .C2(n_613), .Y(n_666) );
OAI21xp33_ASAP7_75t_SL g667 ( .A1(n_607), .A2(n_594), .B(n_621), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_622), .A2(n_606), .B(n_611), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_609), .B(n_592), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_614), .A2(n_601), .B1(n_599), .B2(n_628), .C(n_589), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_608), .A2(n_615), .B(n_617), .C(n_631), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_643), .B(n_649), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_670), .B(n_665), .C(n_648), .D(n_636), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g674 ( .A1(n_664), .A2(n_656), .B(n_642), .C(n_671), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_654), .Y(n_675) );
AOI21xp33_ASAP7_75t_SL g676 ( .A1(n_652), .A2(n_641), .B(n_666), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_645), .A2(n_647), .B1(n_644), .B2(n_646), .Y(n_677) );
NAND4xp25_ASAP7_75t_SL g678 ( .A(n_641), .B(n_667), .C(n_640), .D(n_639), .Y(n_678) );
NAND4xp75_ASAP7_75t_L g679 ( .A(n_672), .B(n_660), .C(n_658), .D(n_668), .Y(n_679) );
NOR3xp33_ASAP7_75t_SL g680 ( .A(n_678), .B(n_657), .C(n_653), .Y(n_680) );
XOR2xp5_ASAP7_75t_L g681 ( .A(n_673), .B(n_651), .Y(n_681) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_674), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_679), .Y(n_683) );
NAND4xp75_ASAP7_75t_L g684 ( .A(n_680), .B(n_676), .C(n_661), .D(n_659), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_682), .B(n_677), .C(n_650), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_683), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_685), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_686), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_687), .Y(n_689) );
INVxp33_ASAP7_75t_L g690 ( .A(n_688), .Y(n_690) );
XNOR2x1_ASAP7_75t_L g691 ( .A(n_689), .B(n_684), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_690), .A2(n_689), .B1(n_691), .B2(n_675), .C1(n_681), .C2(n_635), .Y(n_692) );
AOI21xp33_ASAP7_75t_SL g693 ( .A1(n_692), .A2(n_652), .B(n_637), .Y(n_693) );
AO21x2_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_663), .B(n_638), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_669), .B1(n_662), .B2(n_655), .Y(n_695) );
endmodule