module fake_ibex_847_n_6460 (n_151, n_1084, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1104, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_1090, n_177, n_1110, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_1097, n_9, n_1079, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_1080, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_1106, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_1098, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_1096, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_1109, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_1112, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_1099, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_1103, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_1081, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_1117, n_30, n_1101, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_1083, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_1116, n_623, n_585, n_1030, n_1094, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_1082, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_1120, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_1089, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_1092, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_1115, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1100, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1078, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_1086, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_1118, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_1087, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_1114, n_409, n_1093, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_1107, n_223, n_381, n_1073, n_1108, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_1111, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_1113, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_1119, n_903, n_519, n_345, n_408, n_119, n_1085, n_361, n_1095, n_455, n_419, n_774, n_72, n_1048, n_319, n_1091, n_195, n_885, n_513, n_212, n_588, n_877, n_1121, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_1088, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_1102, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_1105, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_6460);

input n_151;
input n_1084;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1104;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_1090;
input n_177;
input n_1110;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_1097;
input n_9;
input n_1079;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_1080;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_1106;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_1098;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_1096;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_1109;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_1112;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_1099;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_1103;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_1081;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_1117;
input n_30;
input n_1101;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_1083;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_1116;
input n_623;
input n_585;
input n_1030;
input n_1094;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_1082;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_1120;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_1089;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_1092;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_1115;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1100;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1078;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_1086;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_1118;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_1087;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_1114;
input n_409;
input n_1093;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_1107;
input n_223;
input n_381;
input n_1073;
input n_1108;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_1111;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_1113;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_1119;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_1085;
input n_361;
input n_1095;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_1091;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_1121;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_1088;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_1102;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_1105;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_6460;

wire n_4557;
wire n_6210;
wire n_5285;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_3147;
wire n_3983;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3529;
wire n_3222;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4625;
wire n_4151;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_5566;
wire n_6185;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_1878;
wire n_4803;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_2982;
wire n_2634;
wire n_3124;
wire n_5384;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2682;
wire n_1666;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6117;
wire n_1312;
wire n_5844;
wire n_6448;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6361;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_2463;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5755;
wire n_5098;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5862;
wire n_5869;
wire n_1238;
wire n_3959;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_5489;
wire n_2316;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_3223;
wire n_2005;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_5940;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_3261;
wire n_5324;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5510;
wire n_5329;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_5618;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6420;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_2565;
wire n_4201;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_5359;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4681;
wire n_4253;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_5985;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_2300;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_2833;
wire n_1750;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5595;
wire n_5334;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_2684;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_6356;
wire n_5313;
wire n_2108;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6364;
wire n_5715;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_1770;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_5853;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2855;
wire n_2653;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_5377;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6175;
wire n_5279;
wire n_4650;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5523;
wire n_5456;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_5214;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6214;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5855;
wire n_5819;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_3449;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5992;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_3940;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_6075;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_1161;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_1193;
wire n_3557;
wire n_3380;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5594;
wire n_5335;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_5393;
wire n_4782;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

INVx1_ASAP7_75t_L g1122 ( 
.A(n_767),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_9),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_86),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1096),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_897),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_482),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_556),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_672),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_398),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_990),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_866),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_571),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1110),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_614),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_238),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_200),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1042),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_907),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1064),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_62),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_407),
.Y(n_1142)
);

BUFx10_ASAP7_75t_L g1143 ( 
.A(n_795),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_153),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_492),
.Y(n_1145)
);

BUFx5_ASAP7_75t_L g1146 ( 
.A(n_970),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_300),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1029),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_642),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_7),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1081),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_482),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1058),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_1064),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_875),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_875),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_312),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_402),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_547),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1043),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_435),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_487),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_543),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_526),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_178),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1110),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_597),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_713),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_678),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_284),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_697),
.Y(n_1171)
);

BUFx10_ASAP7_75t_L g1172 ( 
.A(n_1056),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_349),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_338),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_789),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_485),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_931),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_1046),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_412),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_91),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_559),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_720),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1019),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1055),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_806),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_240),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_485),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_967),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_192),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_821),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1053),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_481),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_681),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_948),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_409),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_530),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_360),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_900),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_978),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_52),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_748),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_10),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_27),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_623),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_290),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_991),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_384),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_449),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_475),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_320),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_499),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_708),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_38),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1068),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1079),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_890),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1063),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_107),
.Y(n_1218)
);

CKINVDCx16_ASAP7_75t_R g1219 ( 
.A(n_350),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_347),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_140),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_444),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_90),
.Y(n_1223)
);

BUFx8_ASAP7_75t_SL g1224 ( 
.A(n_410),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_709),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1093),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_695),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_738),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_610),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_749),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1062),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_559),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_152),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_785),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_308),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_820),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_419),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_908),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_355),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_317),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_159),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_644),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_111),
.Y(n_1243)
);

BUFx5_ASAP7_75t_L g1244 ( 
.A(n_941),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_164),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_791),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_460),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_976),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_355),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1070),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_769),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_378),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_771),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_599),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_966),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1023),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_9),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_677),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_889),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_786),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1069),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1039),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1077),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_622),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_757),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_129),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_233),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_978),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_416),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_210),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_114),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_57),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_84),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_602),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_510),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1013),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_407),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1073),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_615),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_908),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1083),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1015),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_786),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_726),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_604),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_399),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_933),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_386),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_823),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_455),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_244),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_750),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1106),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_587),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_518),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1069),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_711),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1025),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_320),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_718),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_536),
.Y(n_1301)
);

BUFx10_ASAP7_75t_L g1302 ( 
.A(n_725),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_442),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_571),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_754),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_768),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_194),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_847),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_104),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_759),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_573),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_697),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_306),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_281),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1108),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_20),
.Y(n_1316)
);

CKINVDCx16_ASAP7_75t_R g1317 ( 
.A(n_426),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_146),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_25),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_744),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_48),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_433),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_955),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_583),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_329),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_477),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_386),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_320),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_333),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_493),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_451),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1012),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_719),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_836),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_992),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_387),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_544),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_57),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_155),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_417),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_50),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_498),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1082),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_398),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_899),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_782),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_659),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_493),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_151),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_152),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_118),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1092),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1047),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1027),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_538),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_952),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_892),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_420),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_579),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_974),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_805),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_344),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_991),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1078),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_615),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_718),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1097),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_237),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_739),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_135),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_293),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_205),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_532),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_185),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_404),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_612),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_348),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_88),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_993),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_953),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1008),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_514),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_961),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_673),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_445),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_652),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_128),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_530),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_527),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_59),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1054),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_246),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_740),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_588),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_953),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_843),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_524),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_68),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_561),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_472),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1067),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_796),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1042),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_903),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_352),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_732),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_394),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_968),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1078),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_401),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_869),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_353),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_98),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_598),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_881),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_710),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_727),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_504),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_484),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_788),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_970),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_108),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_731),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_735),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_39),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_294),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1074),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1114),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1079),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_959),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_159),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_628),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_610),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_4),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_165),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_993),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1019),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_40),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_909),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_752),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_811),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1041),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_695),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_732),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_242),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1048),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_270),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_19),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_467),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_799),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_74),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_388),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1115),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_43),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_131),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_664),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_479),
.Y(n_1457)
);

BUFx5_ASAP7_75t_L g1458 ( 
.A(n_400),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_285),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_425),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_809),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_352),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_532),
.Y(n_1463)
);

BUFx10_ASAP7_75t_L g1464 ( 
.A(n_831),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_995),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_995),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_513),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_236),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_822),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_325),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_644),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_687),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_598),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_363),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_961),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_64),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_992),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_10),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_742),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_41),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_85),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1060),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_391),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1080),
.Y(n_1484)
);

BUFx10_ASAP7_75t_L g1485 ( 
.A(n_740),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_78),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_496),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1095),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1044),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_516),
.Y(n_1490)
);

BUFx5_ASAP7_75t_L g1491 ( 
.A(n_478),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_755),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_495),
.Y(n_1493)
);

BUFx10_ASAP7_75t_L g1494 ( 
.A(n_421),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_485),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1116),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_957),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_539),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_733),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_876),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_152),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_534),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1029),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_458),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_332),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_127),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_403),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_75),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_15),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_417),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_866),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_228),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_79),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1087),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_70),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1094),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_951),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_483),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_976),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1061),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_861),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_73),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1018),
.Y(n_1523)
);

CKINVDCx14_ASAP7_75t_R g1524 ( 
.A(n_104),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_131),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_211),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1090),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_661),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_282),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_91),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_580),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_276),
.Y(n_1532)
);

CKINVDCx16_ASAP7_75t_R g1533 ( 
.A(n_342),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_408),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_244),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_548),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1050),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_90),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_798),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_678),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_785),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1084),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_967),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_946),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_565),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_510),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_430),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1068),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_411),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1046),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_469),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_119),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_939),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1049),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_850),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_85),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_570),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_801),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_58),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_688),
.Y(n_1560)
);

BUFx10_ASAP7_75t_L g1561 ( 
.A(n_923),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_265),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_348),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_635),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_113),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_960),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_273),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_197),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_188),
.Y(n_1569)
);

BUFx5_ASAP7_75t_L g1570 ( 
.A(n_871),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_578),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_391),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1118),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1032),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1089),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_948),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_644),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_420),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_737),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_112),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_100),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_243),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_674),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_137),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_855),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_361),
.Y(n_1586)
);

CKINVDCx16_ASAP7_75t_R g1587 ( 
.A(n_1009),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1071),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_996),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_672),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1024),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_951),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_387),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_751),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_538),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1011),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_490),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_563),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_102),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_932),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_489),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_138),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_264),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_694),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_929),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_734),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1076),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1086),
.Y(n_1608)
);

CKINVDCx14_ASAP7_75t_R g1609 ( 
.A(n_201),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_511),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_874),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_938),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_951),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_151),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_47),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_278),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_965),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_351),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_235),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1023),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1065),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_294),
.Y(n_1622)
);

CKINVDCx14_ASAP7_75t_R g1623 ( 
.A(n_1081),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_303),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_241),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_422),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_852),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_821),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_901),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_204),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_137),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_915),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_355),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_751),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_113),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_171),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_755),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_761),
.Y(n_1638)
);

BUFx5_ASAP7_75t_L g1639 ( 
.A(n_390),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1066),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_483),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_325),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1040),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1109),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_952),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_155),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_289),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_65),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_891),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_870),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_563),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1075),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1085),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_367),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1111),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1032),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_268),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_872),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_765),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_859),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1072),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_631),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_851),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1091),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_857),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_909),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_152),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_539),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_779),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_621),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_660),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1045),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_701),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_477),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_735),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_155),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_656),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_358),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_227),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_615),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_261),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_811),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_459),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_933),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_980),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_254),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_397),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_906),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_890),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_654),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_849),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1053),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_846),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_302),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_672),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1022),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_958),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_548),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1085),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1098),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_750),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1100),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_875),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1099),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_593),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_188),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1059),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_86),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_456),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1095),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_420),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_535),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_198),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1005),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_680),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_882),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1103),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_983),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_646),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_614),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_117),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_157),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_834),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_786),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1028),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_516),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_629),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_443),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_66),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_920),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_388),
.Y(n_1731)
);

BUFx10_ASAP7_75t_L g1732 ( 
.A(n_294),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_86),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1052),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_324),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_715),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_353),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_585),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_566),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_296),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_12),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_154),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_671),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_872),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_169),
.Y(n_1745)
);

CKINVDCx14_ASAP7_75t_R g1746 ( 
.A(n_146),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_575),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_871),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_831),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_883),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_611),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_948),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_998),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_25),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_59),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_335),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_247),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1057),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_911),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_239),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_356),
.Y(n_1761)
);

CKINVDCx14_ASAP7_75t_R g1762 ( 
.A(n_1000),
.Y(n_1762)
);

BUFx5_ASAP7_75t_L g1763 ( 
.A(n_1096),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1038),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_251),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_867),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1114),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_535),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_154),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1042),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1040),
.Y(n_1771)
);

BUFx10_ASAP7_75t_L g1772 ( 
.A(n_203),
.Y(n_1772)
);

BUFx8_ASAP7_75t_SL g1773 ( 
.A(n_1068),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_586),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1057),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_86),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_338),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_843),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_126),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1051),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_234),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1103),
.Y(n_1782)
);

BUFx10_ASAP7_75t_L g1783 ( 
.A(n_789),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_759),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1075),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_217),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_141),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_304),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1045),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_607),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_302),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1088),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_907),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_977),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_518),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_5),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_343),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_860),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_222),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_854),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_491),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_2),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1772),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1203),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1772),
.Y(n_1805)
);

INVxp33_ASAP7_75t_L g1806 ( 
.A(n_1481),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1146),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1772),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1552),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1321),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1137),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1146),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1273),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1273),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1150),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_1524),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1165),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1526),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1524),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1180),
.Y(n_1820)
);

INVxp33_ASAP7_75t_SL g1821 ( 
.A(n_1347),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1609),
.Y(n_1822)
);

CKINVDCx16_ASAP7_75t_R g1823 ( 
.A(n_1351),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1200),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1218),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1241),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1307),
.Y(n_1827)
);

INVxp67_ASAP7_75t_SL g1828 ( 
.A(n_1526),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1350),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1609),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1746),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1413),
.Y(n_1832)
);

BUFx2_ASAP7_75t_SL g1833 ( 
.A(n_1569),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1146),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1146),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1422),
.Y(n_1836)
);

CKINVDCx20_ASAP7_75t_R g1837 ( 
.A(n_1746),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1431),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1569),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1582),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1434),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1435),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1454),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1582),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1509),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1235),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1525),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1623),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1556),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1584),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1599),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1623),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1602),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1636),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1667),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1729),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1741),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1762),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1760),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1776),
.Y(n_1860)
);

CKINVDCx20_ASAP7_75t_R g1861 ( 
.A(n_1370),
.Y(n_1861)
);

INVxp33_ASAP7_75t_L g1862 ( 
.A(n_1527),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1786),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1762),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1523),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1799),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1515),
.Y(n_1867)
);

INVxp33_ASAP7_75t_L g1868 ( 
.A(n_1540),
.Y(n_1868)
);

INVxp33_ASAP7_75t_L g1869 ( 
.A(n_1564),
.Y(n_1869)
);

CKINVDCx16_ASAP7_75t_R g1870 ( 
.A(n_1219),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1706),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1159),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1263),
.Y(n_1873)
);

CKINVDCx14_ASAP7_75t_R g1874 ( 
.A(n_1133),
.Y(n_1874)
);

INVxp33_ASAP7_75t_L g1875 ( 
.A(n_1681),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1337),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1650),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1790),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1538),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1557),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1737),
.Y(n_1881)
);

BUFx10_ASAP7_75t_L g1882 ( 
.A(n_1796),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1370),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1224),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1598),
.Y(n_1885)
);

CKINVDCx16_ASAP7_75t_R g1886 ( 
.A(n_1317),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1613),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1785),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1785),
.Y(n_1889)
);

INVxp33_ASAP7_75t_L g1890 ( 
.A(n_1747),
.Y(n_1890)
);

CKINVDCx16_ASAP7_75t_R g1891 ( 
.A(n_1459),
.Y(n_1891)
);

INVxp67_ASAP7_75t_SL g1892 ( 
.A(n_1339),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1271),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1271),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1372),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1146),
.Y(n_1896)
);

INVxp67_ASAP7_75t_SL g1897 ( 
.A(n_1318),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1224),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1259),
.Y(n_1899)
);

INVxp67_ASAP7_75t_SL g1900 ( 
.A(n_1318),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1259),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1122),
.Y(n_1902)
);

INVxp67_ASAP7_75t_SL g1903 ( 
.A(n_1387),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1125),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1135),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1139),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1773),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1147),
.Y(n_1908)
);

CKINVDCx20_ASAP7_75t_R g1909 ( 
.A(n_1372),
.Y(n_1909)
);

INVxp33_ASAP7_75t_L g1910 ( 
.A(n_1773),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1149),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1123),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1802),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1781),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1124),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1156),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1158),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1160),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1162),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1167),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1174),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1787),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1188),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1191),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_1438),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1136),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1194),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1195),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1438),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1197),
.Y(n_1930)
);

CKINVDCx14_ASAP7_75t_R g1931 ( 
.A(n_1133),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1199),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1141),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1206),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1210),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1211),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1533),
.B(n_0),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1212),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1146),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1288),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1144),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1214),
.Y(n_1942)
);

CKINVDCx20_ASAP7_75t_R g1943 ( 
.A(n_1580),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1146),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1133),
.Y(n_1945)
);

INVxp33_ASAP7_75t_SL g1946 ( 
.A(n_1189),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1805),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1804),
.B(n_1288),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1813),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1805),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1882),
.Y(n_1951)
);

CKINVDCx8_ASAP7_75t_R g1952 ( 
.A(n_1823),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1833),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1893),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1804),
.A2(n_1202),
.B1(n_1213),
.B2(n_1186),
.Y(n_1955)
);

XNOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1884),
.B(n_1126),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1811),
.A2(n_1476),
.B(n_1387),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1807),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1892),
.B(n_1221),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1944),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1874),
.Y(n_1961)
);

INVx2_ASAP7_75t_SL g1962 ( 
.A(n_1882),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1815),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1817),
.A2(n_1508),
.B(n_1476),
.Y(n_1964)
);

INVx3_ASAP7_75t_L g1965 ( 
.A(n_1945),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1812),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1821),
.A2(n_1646),
.B1(n_1580),
.B2(n_1621),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1820),
.Y(n_1968)
);

CKINVDCx6p67_ASAP7_75t_R g1969 ( 
.A(n_1870),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1824),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1879),
.B(n_1353),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1825),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1806),
.A2(n_1233),
.B1(n_1245),
.B2(n_1243),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1893),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1945),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1862),
.B(n_1143),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1826),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1894),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1834),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1858),
.B(n_1353),
.Y(n_1980)
);

AND2x6_ASAP7_75t_L g1981 ( 
.A(n_1803),
.B(n_1367),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1808),
.B(n_1587),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1835),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1814),
.B(n_1839),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1868),
.B(n_1143),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1894),
.Y(n_1986)
);

CKINVDCx6p67_ASAP7_75t_R g1987 ( 
.A(n_1886),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1814),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1896),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1939),
.Y(n_1990)
);

BUFx8_ASAP7_75t_L g1991 ( 
.A(n_1865),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1888),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1819),
.B(n_1266),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1839),
.Y(n_1994)
);

AND2x6_ASAP7_75t_L g1995 ( 
.A(n_1937),
.B(n_1367),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1827),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1889),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_SL g1998 ( 
.A1(n_1861),
.A2(n_1168),
.B1(n_1277),
.B2(n_1153),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1899),
.Y(n_1999)
);

XNOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1898),
.B(n_1127),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1901),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1840),
.B(n_1272),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1867),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1840),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_SL g2005 ( 
.A1(n_1883),
.A2(n_1168),
.B1(n_1277),
.B2(n_1153),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1869),
.B(n_1143),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1829),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1844),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1844),
.B(n_1291),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1846),
.B(n_1432),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1931),
.B(n_1309),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1832),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1871),
.Y(n_2013)
);

INVx5_ASAP7_75t_L g2014 ( 
.A(n_1891),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1836),
.Y(n_2015)
);

AND2x6_ASAP7_75t_L g2016 ( 
.A(n_1809),
.B(n_1432),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1818),
.Y(n_2017)
);

AND2x6_ASAP7_75t_L g2018 ( 
.A(n_1914),
.B(n_1505),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1872),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1822),
.B(n_1319),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1828),
.Y(n_2021)
);

AND2x2_ASAP7_75t_SL g2022 ( 
.A(n_1912),
.B(n_1128),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1946),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1873),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1876),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1940),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1877),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1940),
.B(n_1338),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1830),
.B(n_1341),
.Y(n_2029)
);

BUFx3_ASAP7_75t_L g2030 ( 
.A(n_1913),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1897),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1838),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1902),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1915),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1841),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1900),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1846),
.B(n_1349),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1904),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1905),
.Y(n_2039)
);

BUFx3_ASAP7_75t_L g2040 ( 
.A(n_1922),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1816),
.A2(n_1368),
.B1(n_1378),
.B2(n_1374),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1837),
.A2(n_1890),
.B1(n_1875),
.B2(n_1831),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1878),
.B(n_1505),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_1926),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1842),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1903),
.B(n_1390),
.Y(n_2046)
);

INVx4_ASAP7_75t_L g2047 ( 
.A(n_1933),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1906),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1843),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1908),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1881),
.B(n_1810),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1880),
.B(n_1685),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1885),
.B(n_1685),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1911),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1941),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1916),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1845),
.B(n_1398),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1887),
.B(n_1178),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1847),
.B(n_1425),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1849),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1850),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1917),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1918),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1851),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1848),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1919),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1852),
.A2(n_1445),
.B1(n_1451),
.B2(n_1448),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1853),
.B(n_1455),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1854),
.B(n_1468),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1920),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1855),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1921),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1864),
.Y(n_2073)
);

AND2x2_ASAP7_75t_SL g2074 ( 
.A(n_1910),
.B(n_1128),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1856),
.Y(n_2075)
);

OAI22xp5_ASAP7_75t_SL g2076 ( 
.A1(n_1895),
.A2(n_1310),
.B1(n_1325),
.B2(n_1282),
.Y(n_2076)
);

BUFx8_ASAP7_75t_L g2077 ( 
.A(n_1907),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1909),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1857),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1859),
.Y(n_2080)
);

OA21x2_ASAP7_75t_L g2081 ( 
.A1(n_1860),
.A2(n_1559),
.B(n_1508),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1863),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1923),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1924),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1866),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1927),
.Y(n_2086)
);

INVx4_ASAP7_75t_L g2087 ( 
.A(n_1928),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1930),
.Y(n_2088)
);

INVx3_ASAP7_75t_L g2089 ( 
.A(n_1932),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1934),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_SL g2091 ( 
.A(n_1935),
.B(n_1478),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1936),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1938),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_1942),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_1925),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1929),
.A2(n_1480),
.B1(n_1501),
.B2(n_1486),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1943),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_1813),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_1804),
.B(n_1700),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_SL g2100 ( 
.A(n_1879),
.B(n_1506),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1807),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1805),
.B(n_1512),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1813),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1833),
.Y(n_2104)
);

BUFx12f_ASAP7_75t_L g2105 ( 
.A(n_1882),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1813),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1823),
.A2(n_1513),
.B1(n_1530),
.B2(n_1522),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1813),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1833),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1833),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1813),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1813),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1805),
.B(n_1535),
.Y(n_2113)
);

BUFx6f_ASAP7_75t_L g2114 ( 
.A(n_1813),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1833),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1813),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1821),
.A2(n_1646),
.B1(n_1568),
.B2(n_1615),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1833),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1813),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_1813),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1821),
.A2(n_1614),
.B1(n_1625),
.B2(n_1619),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1806),
.B(n_1152),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1833),
.Y(n_2123)
);

OAI21x1_ASAP7_75t_L g2124 ( 
.A1(n_1805),
.A2(n_1565),
.B(n_1559),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1813),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_1813),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1805),
.B(n_1630),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_SL g2128 ( 
.A1(n_1861),
.A2(n_1310),
.B1(n_1325),
.B2(n_1282),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1833),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1823),
.A2(n_1631),
.B1(n_1676),
.B2(n_1648),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1805),
.B(n_1679),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1805),
.B(n_1708),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1813),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1813),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1813),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1805),
.B(n_1721),
.Y(n_2136)
);

INVxp67_ASAP7_75t_SL g2137 ( 
.A(n_1806),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_1805),
.A2(n_1581),
.B(n_1565),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_1879),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_1805),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1833),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1813),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1813),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1805),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1813),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1806),
.B(n_1152),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_1813),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1806),
.B(n_1152),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1805),
.B(n_1722),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1813),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1813),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1821),
.A2(n_1745),
.B1(n_1754),
.B2(n_1742),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1833),
.Y(n_2153)
);

CKINVDCx6p67_ASAP7_75t_R g2154 ( 
.A(n_1823),
.Y(n_2154)
);

OA21x2_ASAP7_75t_L g2155 ( 
.A1(n_1807),
.A2(n_1635),
.B(n_1581),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_1821),
.A2(n_1769),
.B1(n_1779),
.B2(n_1755),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1813),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1833),
.Y(n_2158)
);

OAI22x1_ASAP7_75t_L g2159 ( 
.A1(n_1937),
.A2(n_1130),
.B1(n_1132),
.B2(n_1129),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1813),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1805),
.B(n_1134),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_1805),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1813),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1807),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1813),
.Y(n_2165)
);

INVx5_ASAP7_75t_L g2166 ( 
.A(n_1805),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1805),
.B(n_1138),
.Y(n_2167)
);

INVxp33_ASAP7_75t_SL g2168 ( 
.A(n_1879),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1805),
.B(n_1140),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1813),
.Y(n_2170)
);

NAND2xp33_ASAP7_75t_L g2171 ( 
.A(n_1819),
.B(n_1244),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1804),
.B(n_1700),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1813),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1805),
.B(n_1142),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1806),
.B(n_1154),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1833),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1945),
.B(n_1514),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1813),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1945),
.B(n_1148),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1954),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_2168),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_2139),
.Y(n_2182)
);

CKINVDCx16_ASAP7_75t_R g2183 ( 
.A(n_2105),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_2154),
.Y(n_2184)
);

CKINVDCx16_ASAP7_75t_R g2185 ( 
.A(n_2100),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_R g2186 ( 
.A(n_1961),
.B(n_1223),
.Y(n_2186)
);

BUFx2_ASAP7_75t_L g2187 ( 
.A(n_2137),
.Y(n_2187)
);

CKINVDCx20_ASAP7_75t_R g2188 ( 
.A(n_2078),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_2023),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1974),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1969),
.Y(n_2191)
);

BUFx10_ASAP7_75t_L g2192 ( 
.A(n_1951),
.Y(n_2192)
);

AOI21x1_ASAP7_75t_L g2193 ( 
.A1(n_1957),
.A2(n_1964),
.B(n_2124),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1978),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1987),
.Y(n_2195)
);

CKINVDCx20_ASAP7_75t_R g2196 ( 
.A(n_1991),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_2034),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1952),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_2122),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1986),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_2081),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_2042),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_2077),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2003),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2013),
.Y(n_2205)
);

CKINVDCx20_ASAP7_75t_R g2206 ( 
.A(n_1998),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2019),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2025),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2138),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1947),
.B(n_1151),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2081),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_2096),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_2122),
.Y(n_2213)
);

CKINVDCx16_ASAP7_75t_R g2214 ( 
.A(n_2030),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_2040),
.Y(n_2215)
);

NOR2xp67_ASAP7_75t_L g2216 ( 
.A(n_2014),
.B(n_0),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_R g2217 ( 
.A(n_2091),
.B(n_1713),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_2044),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2146),
.B(n_1154),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2027),
.Y(n_2220)
);

NOR2x1p5_ASAP7_75t_L g2221 ( 
.A(n_1951),
.B(n_1155),
.Y(n_2221)
);

CKINVDCx20_ASAP7_75t_R g2222 ( 
.A(n_2005),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_2055),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2155),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2146),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_R g2226 ( 
.A(n_1962),
.B(n_2014),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_2098),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_2076),
.Y(n_2228)
);

HB1xp67_ASAP7_75t_L g2229 ( 
.A(n_2148),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2128),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_R g2231 ( 
.A(n_2014),
.B(n_1346),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2107),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1984),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_2130),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1973),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_R g2236 ( 
.A(n_2095),
.B(n_2065),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_2117),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_2041),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2148),
.B(n_1562),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_R g2240 ( 
.A(n_2073),
.B(n_1346),
.Y(n_2240)
);

CKINVDCx20_ASAP7_75t_R g2241 ( 
.A(n_1967),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_1955),
.Y(n_2242)
);

CKINVDCx20_ASAP7_75t_R g2243 ( 
.A(n_2047),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2155),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2032),
.Y(n_2245)
);

CKINVDCx20_ASAP7_75t_R g2246 ( 
.A(n_2121),
.Y(n_2246)
);

NAND2xp33_ASAP7_75t_SL g2247 ( 
.A(n_2175),
.B(n_1161),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_R g2248 ( 
.A(n_2175),
.B(n_1379),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1976),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_1976),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2035),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2080),
.Y(n_2252)
);

CKINVDCx20_ASAP7_75t_R g2253 ( 
.A(n_2152),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1963),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1985),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_2166),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1985),
.Y(n_2257)
);

CKINVDCx20_ASAP7_75t_R g2258 ( 
.A(n_2156),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_2006),
.Y(n_2259)
);

BUFx10_ASAP7_75t_L g2260 ( 
.A(n_2018),
.Y(n_2260)
);

CKINVDCx16_ASAP7_75t_R g2261 ( 
.A(n_2006),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_2067),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2022),
.A2(n_1982),
.B1(n_2037),
.B2(n_2051),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2011),
.B(n_1154),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_1971),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2024),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2031),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1963),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2036),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1968),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_2098),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2097),
.Y(n_2272)
);

CKINVDCx20_ASAP7_75t_R g2273 ( 
.A(n_2051),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_2018),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_2018),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2002),
.B(n_1244),
.Y(n_2276)
);

CKINVDCx5p33_ASAP7_75t_R g2277 ( 
.A(n_2074),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_1959),
.B(n_1131),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_2159),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_2159),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_2016),
.Y(n_2281)
);

BUFx3_ASAP7_75t_L g2282 ( 
.A(n_2112),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_2016),
.Y(n_2283)
);

CKINVDCx16_ASAP7_75t_R g2284 ( 
.A(n_1995),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1968),
.Y(n_2285)
);

CKINVDCx20_ASAP7_75t_R g2286 ( 
.A(n_2111),
.Y(n_2286)
);

INVx2_ASAP7_75t_SL g2287 ( 
.A(n_1948),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2009),
.B(n_1244),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2089),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_2016),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1995),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1970),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_2112),
.Y(n_2293)
);

INVxp67_ASAP7_75t_SL g2294 ( 
.A(n_2028),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1950),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_R g2296 ( 
.A(n_1995),
.B(n_1379),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1992),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1997),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1999),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2001),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_R g2301 ( 
.A(n_2171),
.B(n_1424),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_2134),
.Y(n_2302)
);

BUFx2_ASAP7_75t_L g2303 ( 
.A(n_1956),
.Y(n_2303)
);

NOR2xp67_ASAP7_75t_L g2304 ( 
.A(n_2140),
.B(n_0),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1970),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2021),
.Y(n_2306)
);

NOR2xp67_ASAP7_75t_L g2307 ( 
.A(n_2144),
.B(n_0),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_2099),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_2114),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_2172),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1972),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_R g2312 ( 
.A(n_1953),
.B(n_1424),
.Y(n_2312)
);

INVxp67_ASAP7_75t_L g2313 ( 
.A(n_2046),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2010),
.B(n_1176),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1972),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_2114),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_L g2317 ( 
.A(n_2162),
.B(n_1965),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_1993),
.Y(n_2318)
);

BUFx10_ASAP7_75t_L g2319 ( 
.A(n_2058),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_2020),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2021),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2094),
.Y(n_2322)
);

CKINVDCx20_ASAP7_75t_R g2323 ( 
.A(n_1975),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_2029),
.Y(n_2324)
);

CKINVDCx20_ASAP7_75t_R g2325 ( 
.A(n_2102),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_2104),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1977),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2094),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_R g2329 ( 
.A(n_2109),
.B(n_1446),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_2110),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1977),
.Y(n_2331)
);

BUFx10_ASAP7_75t_L g2332 ( 
.A(n_2179),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1996),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_2115),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2118),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_2120),
.Y(n_2336)
);

INVxp67_ASAP7_75t_L g2337 ( 
.A(n_2113),
.Y(n_2337)
);

XNOR2xp5_ASAP7_75t_L g2338 ( 
.A(n_2000),
.B(n_1446),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2123),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1996),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_2129),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2057),
.B(n_1244),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2007),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2007),
.Y(n_2344)
);

BUFx10_ASAP7_75t_L g2345 ( 
.A(n_2177),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_1981),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_1980),
.B(n_1172),
.Y(n_2347)
);

CKINVDCx20_ASAP7_75t_R g2348 ( 
.A(n_2127),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_2141),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2012),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_R g2351 ( 
.A(n_2153),
.B(n_1471),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2012),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_2158),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2043),
.B(n_1663),
.Y(n_2354)
);

CKINVDCx20_ASAP7_75t_R g2355 ( 
.A(n_2131),
.Y(n_2355)
);

AO21x2_ASAP7_75t_L g2356 ( 
.A1(n_2075),
.A2(n_1217),
.B(n_1216),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2015),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2015),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2045),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_2176),
.Y(n_2360)
);

CKINVDCx20_ASAP7_75t_R g2361 ( 
.A(n_2132),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2045),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2049),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2049),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_2120),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_2125),
.Y(n_2366)
);

INVx3_ASAP7_75t_L g2367 ( 
.A(n_2166),
.Y(n_2367)
);

CKINVDCx16_ASAP7_75t_R g2368 ( 
.A(n_1981),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2125),
.Y(n_2369)
);

NAND2xp33_ASAP7_75t_R g2370 ( 
.A(n_2052),
.B(n_1163),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2126),
.Y(n_2371)
);

CKINVDCx5p33_ASAP7_75t_R g2372 ( 
.A(n_2126),
.Y(n_2372)
);

BUFx3_ASAP7_75t_L g2373 ( 
.A(n_2133),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1949),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2133),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_2143),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2143),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_2147),
.Y(n_2378)
);

NOR2xp67_ASAP7_75t_L g2379 ( 
.A(n_2166),
.B(n_1),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2103),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_2147),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2053),
.B(n_1727),
.Y(n_2382)
);

INVx3_ASAP7_75t_L g2383 ( 
.A(n_2150),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_1981),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_R g2385 ( 
.A(n_1988),
.B(n_1471),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2106),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2108),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2150),
.Y(n_2388)
);

NOR2xp67_ASAP7_75t_L g2389 ( 
.A(n_2161),
.B(n_1),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_2170),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2017),
.Y(n_2391)
);

OA21x2_ASAP7_75t_L g2392 ( 
.A1(n_1958),
.A2(n_1733),
.B(n_1635),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_R g2393 ( 
.A(n_1994),
.B(n_1511),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2075),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_R g2395 ( 
.A(n_2004),
.B(n_1511),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2170),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2033),
.Y(n_2397)
);

CKINVDCx20_ASAP7_75t_R g2398 ( 
.A(n_2149),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2038),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2178),
.Y(n_2400)
);

CKINVDCx20_ASAP7_75t_R g2401 ( 
.A(n_2178),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2116),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_2059),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_R g2404 ( 
.A(n_2008),
.B(n_1607),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2119),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_2167),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2169),
.Y(n_2407)
);

CKINVDCx5p33_ASAP7_75t_R g2408 ( 
.A(n_2068),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_2069),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_2136),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2039),
.Y(n_2411)
);

CKINVDCx20_ASAP7_75t_R g2412 ( 
.A(n_2174),
.Y(n_2412)
);

INVx1_ASAP7_75t_SL g2413 ( 
.A(n_2026),
.Y(n_2413)
);

CKINVDCx16_ASAP7_75t_R g2414 ( 
.A(n_2087),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2048),
.Y(n_2415)
);

NAND2xp33_ASAP7_75t_R g2416 ( 
.A(n_2135),
.B(n_1164),
.Y(n_2416)
);

CKINVDCx5p33_ASAP7_75t_R g2417 ( 
.A(n_2142),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2145),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2151),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_2157),
.Y(n_2420)
);

NOR2xp67_ASAP7_75t_L g2421 ( 
.A(n_2160),
.B(n_1),
.Y(n_2421)
);

AO21x2_ASAP7_75t_L g2422 ( 
.A1(n_1958),
.A2(n_1234),
.B(n_1220),
.Y(n_2422)
);

XOR2xp5_ASAP7_75t_L g2423 ( 
.A(n_2086),
.B(n_1607),
.Y(n_2423)
);

CKINVDCx20_ASAP7_75t_R g2424 ( 
.A(n_2090),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2050),
.Y(n_2425)
);

BUFx10_ASAP7_75t_L g2426 ( 
.A(n_2060),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_2054),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2163),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_2165),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_2173),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_L g2431 ( 
.A(n_2092),
.B(n_1166),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2056),
.Y(n_2432)
);

CKINVDCx20_ASAP7_75t_R g2433 ( 
.A(n_2093),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2062),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2063),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2066),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_2070),
.Y(n_2437)
);

CKINVDCx20_ASAP7_75t_R g2438 ( 
.A(n_2072),
.Y(n_2438)
);

NAND2xp33_ASAP7_75t_R g2439 ( 
.A(n_2061),
.B(n_1169),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2083),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2084),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2088),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2064),
.Y(n_2443)
);

INVx3_ASAP7_75t_L g2444 ( 
.A(n_2071),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2079),
.Y(n_2445)
);

AOI21x1_ASAP7_75t_L g2446 ( 
.A1(n_2101),
.A2(n_1733),
.B(n_1248),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2082),
.Y(n_2447)
);

INVx3_ASAP7_75t_L g2448 ( 
.A(n_2085),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2101),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_2164),
.Y(n_2450)
);

CKINVDCx20_ASAP7_75t_R g2451 ( 
.A(n_2164),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_1966),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_1979),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_1983),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_1989),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_1990),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_1960),
.Y(n_2457)
);

NOR2xp67_ASAP7_75t_L g2458 ( 
.A(n_2139),
.B(n_1),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1954),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2124),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2139),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1954),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_2168),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_R g2464 ( 
.A(n_1961),
.B(n_1626),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_2139),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_R g2466 ( 
.A(n_1961),
.B(n_1626),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_2168),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2168),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1954),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_1954),
.Y(n_2470)
);

CKINVDCx20_ASAP7_75t_R g2471 ( 
.A(n_2139),
.Y(n_2471)
);

CKINVDCx20_ASAP7_75t_R g2472 ( 
.A(n_2139),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2139),
.B(n_1181),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2168),
.Y(n_2474)
);

INVx3_ASAP7_75t_L g2475 ( 
.A(n_2081),
.Y(n_2475)
);

CKINVDCx20_ASAP7_75t_R g2476 ( 
.A(n_2139),
.Y(n_2476)
);

OAI22xp5_ASAP7_75t_SL g2477 ( 
.A1(n_2078),
.A2(n_1637),
.B1(n_1658),
.B2(n_1629),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2168),
.Y(n_2478)
);

BUFx10_ASAP7_75t_L g2479 ( 
.A(n_2139),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2168),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1954),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_1954),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2168),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_2168),
.Y(n_2484)
);

NAND2xp33_ASAP7_75t_R g2485 ( 
.A(n_2168),
.B(n_1171),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_1947),
.B(n_1173),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2124),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2168),
.Y(n_2488)
);

INVxp67_ASAP7_75t_L g2489 ( 
.A(n_2139),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2168),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2449),
.Y(n_2491)
);

INVx4_ASAP7_75t_L g2492 ( 
.A(n_2183),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2443),
.Y(n_2493)
);

OR2x2_ASAP7_75t_L g2494 ( 
.A(n_2473),
.B(n_1198),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2465),
.B(n_1629),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2471),
.Y(n_2496)
);

INVx3_ASAP7_75t_L g2497 ( 
.A(n_2479),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2426),
.B(n_1177),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2261),
.B(n_1175),
.Y(n_2499)
);

AOI22xp33_ASAP7_75t_L g2500 ( 
.A1(n_2233),
.A2(n_1797),
.B1(n_1658),
.B2(n_1680),
.Y(n_2500)
);

BUFx3_ASAP7_75t_L g2501 ( 
.A(n_2472),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2443),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2444),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2444),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_2199),
.B(n_1179),
.Y(n_2505)
);

AND2x4_ASAP7_75t_L g2506 ( 
.A(n_2476),
.B(n_1637),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2403),
.B(n_1185),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2313),
.B(n_1182),
.Y(n_2508)
);

AND2x4_ASAP7_75t_L g2509 ( 
.A(n_2243),
.B(n_1680),
.Y(n_2509)
);

OR2x6_ASAP7_75t_L g2510 ( 
.A(n_2477),
.B(n_2489),
.Y(n_2510)
);

INVx2_ASAP7_75t_SL g2511 ( 
.A(n_2479),
.Y(n_2511)
);

INVx1_ASAP7_75t_SL g2512 ( 
.A(n_2182),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2337),
.B(n_2294),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2461),
.B(n_1770),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2448),
.Y(n_2515)
);

OR2x2_ASAP7_75t_SL g2516 ( 
.A(n_2185),
.B(n_1770),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2192),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2448),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2201),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2408),
.B(n_1226),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2239),
.A2(n_1797),
.B1(n_1788),
.B2(n_1172),
.Y(n_2521)
);

INVx1_ASAP7_75t_SL g2522 ( 
.A(n_2451),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2426),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2306),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2321),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2267),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2192),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2271),
.Y(n_2528)
);

INVxp67_ASAP7_75t_SL g2529 ( 
.A(n_2438),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2269),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2409),
.B(n_1229),
.Y(n_2531)
);

AND2x4_ASAP7_75t_SL g2532 ( 
.A(n_2286),
.B(n_1788),
.Y(n_2532)
);

BUFx2_ASAP7_75t_L g2533 ( 
.A(n_2217),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2271),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2180),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2414),
.B(n_1183),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_2181),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2213),
.B(n_1231),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2201),
.Y(n_2539)
);

INVx4_ASAP7_75t_SL g2540 ( 
.A(n_2239),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2475),
.Y(n_2541)
);

BUFx3_ASAP7_75t_L g2542 ( 
.A(n_2401),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2190),
.Y(n_2543)
);

INVx1_ASAP7_75t_SL g2544 ( 
.A(n_2463),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2194),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2467),
.B(n_1236),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2468),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2406),
.B(n_1184),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2200),
.Y(n_2549)
);

OAI221xp5_ASAP7_75t_L g2550 ( 
.A1(n_2263),
.A2(n_1793),
.B1(n_1320),
.B2(n_1360),
.C(n_1314),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2459),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2474),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2227),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2445),
.B(n_1187),
.Y(n_2554)
);

INVx4_ASAP7_75t_L g2555 ( 
.A(n_2478),
.Y(n_2555)
);

INVx4_ASAP7_75t_L g2556 ( 
.A(n_2480),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2282),
.Y(n_2557)
);

INVx3_ASAP7_75t_L g2558 ( 
.A(n_2293),
.Y(n_2558)
);

INVx2_ASAP7_75t_SL g2559 ( 
.A(n_2483),
.Y(n_2559)
);

INVxp67_ASAP7_75t_L g2560 ( 
.A(n_2485),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2475),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2462),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2484),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2278),
.B(n_1190),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2211),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2271),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2469),
.Y(n_2567)
);

AND2x6_ASAP7_75t_L g2568 ( 
.A(n_2394),
.B(n_1145),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2488),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_2229),
.B(n_1240),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2470),
.Y(n_2571)
);

INVxp67_ASAP7_75t_L g2572 ( 
.A(n_2187),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2368),
.B(n_1192),
.Y(n_2573)
);

INVx3_ASAP7_75t_L g2574 ( 
.A(n_2373),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2407),
.B(n_1193),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2481),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_SL g2577 ( 
.A(n_2490),
.B(n_1255),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2323),
.B(n_1260),
.Y(n_2578)
);

INVx6_ASAP7_75t_L g2579 ( 
.A(n_2214),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2482),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2450),
.B(n_1196),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2250),
.B(n_1393),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2219),
.B(n_1201),
.Y(n_2583)
);

INVx5_ASAP7_75t_L g2584 ( 
.A(n_2284),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2427),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2193),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2447),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2326),
.B(n_1204),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2347),
.B(n_1402),
.Y(n_2589)
);

BUFx6f_ASAP7_75t_L g2590 ( 
.A(n_2309),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2391),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2204),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2225),
.B(n_1414),
.Y(n_2593)
);

AND2x4_ASAP7_75t_L g2594 ( 
.A(n_2221),
.B(n_2184),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2205),
.Y(n_2595)
);

BUFx3_ASAP7_75t_L g2596 ( 
.A(n_2196),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2413),
.B(n_1205),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2249),
.B(n_1519),
.Y(n_2598)
);

AND3x2_ASAP7_75t_L g2599 ( 
.A(n_2303),
.B(n_2423),
.C(n_2240),
.Y(n_2599)
);

NOR2xp33_ASAP7_75t_L g2600 ( 
.A(n_2255),
.B(n_1537),
.Y(n_2600)
);

BUFx6f_ASAP7_75t_L g2601 ( 
.A(n_2309),
.Y(n_2601)
);

BUFx3_ASAP7_75t_L g2602 ( 
.A(n_2365),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2191),
.B(n_2195),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2207),
.Y(n_2604)
);

BUFx4f_ASAP7_75t_L g2605 ( 
.A(n_2354),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2437),
.B(n_1207),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2208),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2330),
.B(n_2334),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_SL g2609 ( 
.A1(n_2338),
.A2(n_1705),
.B1(n_1697),
.B2(n_1209),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2314),
.B(n_1308),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2220),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2424),
.B(n_1391),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2441),
.B(n_1208),
.Y(n_2613)
);

NOR2xp33_ASAP7_75t_L g2614 ( 
.A(n_2257),
.B(n_1215),
.Y(n_2614)
);

BUFx6f_ASAP7_75t_L g2615 ( 
.A(n_2309),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2335),
.B(n_2339),
.Y(n_2616)
);

BUFx10_ASAP7_75t_L g2617 ( 
.A(n_2203),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2316),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2431),
.B(n_1222),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2397),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2248),
.B(n_1172),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2385),
.B(n_1232),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_2259),
.B(n_1227),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2296),
.Y(n_2624)
);

BUFx6f_ASAP7_75t_L g2625 ( 
.A(n_2316),
.Y(n_2625)
);

AND2x6_ASAP7_75t_L g2626 ( 
.A(n_2224),
.B(n_1145),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2452),
.B(n_1228),
.Y(n_2627)
);

OAI21xp33_ASAP7_75t_L g2628 ( 
.A1(n_2393),
.A2(n_1238),
.B(n_1230),
.Y(n_2628)
);

AND2x6_ASAP7_75t_L g2629 ( 
.A(n_2244),
.B(n_1145),
.Y(n_2629)
);

AND2x6_ASAP7_75t_L g2630 ( 
.A(n_2245),
.B(n_2251),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2399),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2374),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2380),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2341),
.B(n_1239),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2411),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2453),
.B(n_1242),
.Y(n_2636)
);

BUFx3_ASAP7_75t_L g2637 ( 
.A(n_2366),
.Y(n_2637)
);

BUFx10_ASAP7_75t_L g2638 ( 
.A(n_2198),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2395),
.B(n_1232),
.Y(n_2639)
);

CKINVDCx20_ASAP7_75t_R g2640 ( 
.A(n_2231),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2404),
.B(n_1232),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2386),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2433),
.B(n_1482),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2387),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2454),
.B(n_1252),
.Y(n_2645)
);

INVxp33_ASAP7_75t_L g2646 ( 
.A(n_2186),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2415),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2312),
.B(n_1287),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2455),
.B(n_1253),
.Y(n_2649)
);

INVx4_ASAP7_75t_L g2650 ( 
.A(n_2215),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2316),
.Y(n_2651)
);

AND2x6_ASAP7_75t_L g2652 ( 
.A(n_2252),
.B(n_1145),
.Y(n_2652)
);

AND2x6_ASAP7_75t_L g2653 ( 
.A(n_2289),
.B(n_1292),
.Y(n_2653)
);

OR2x2_ASAP7_75t_L g2654 ( 
.A(n_2189),
.B(n_1499),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2319),
.B(n_1254),
.Y(n_2655)
);

AND2x6_ASAP7_75t_L g2656 ( 
.A(n_2266),
.B(n_1292),
.Y(n_2656)
);

INVxp67_ASAP7_75t_SL g2657 ( 
.A(n_2273),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2336),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2425),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2432),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2336),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2349),
.B(n_1264),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2434),
.Y(n_2663)
);

AND2x2_ASAP7_75t_SL g2664 ( 
.A(n_2346),
.B(n_1157),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2329),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2456),
.B(n_1268),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2336),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2405),
.Y(n_2668)
);

NAND3x1_ASAP7_75t_L g2669 ( 
.A(n_2188),
.B(n_1249),
.C(n_1247),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2435),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2436),
.Y(n_2671)
);

AOI22xp33_ASAP7_75t_L g2672 ( 
.A1(n_2235),
.A2(n_1302),
.B1(n_1327),
.B2(n_1287),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2440),
.B(n_1274),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_2464),
.Y(n_2674)
);

INVxp67_ASAP7_75t_SL g2675 ( 
.A(n_2439),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2442),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2353),
.B(n_1275),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2297),
.Y(n_2678)
);

INVx2_ASAP7_75t_SL g2679 ( 
.A(n_2226),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2319),
.B(n_1284),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2360),
.B(n_1290),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2298),
.Y(n_2682)
);

BUFx6f_ASAP7_75t_L g2683 ( 
.A(n_2376),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2351),
.B(n_1287),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2299),
.Y(n_2685)
);

INVx1_ASAP7_75t_SL g2686 ( 
.A(n_2466),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2458),
.B(n_1294),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2218),
.B(n_2223),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2300),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2389),
.B(n_1297),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2295),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2304),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2325),
.B(n_1298),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2210),
.B(n_1299),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2376),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2307),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2209),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2197),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2354),
.B(n_1302),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2236),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2421),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2342),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2276),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2460),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2288),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2237),
.B(n_1576),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2376),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2379),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2369),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2348),
.B(n_1300),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2486),
.B(n_1301),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2216),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2355),
.B(n_1303),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2317),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2383),
.Y(n_2715)
);

AND2x6_ASAP7_75t_L g2716 ( 
.A(n_2256),
.B(n_1292),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2382),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2382),
.B(n_1302),
.Y(n_2718)
);

AOI22xp5_ASAP7_75t_L g2719 ( 
.A1(n_2247),
.A2(n_1306),
.B1(n_1312),
.B2(n_1305),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2384),
.B(n_1313),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2332),
.B(n_1322),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2212),
.B(n_2238),
.Y(n_2722)
);

AND2x6_ASAP7_75t_L g2723 ( 
.A(n_2256),
.B(n_1292),
.Y(n_2723)
);

BUFx3_ASAP7_75t_L g2724 ( 
.A(n_2371),
.Y(n_2724)
);

AND2x6_ASAP7_75t_L g2725 ( 
.A(n_2367),
.B(n_1369),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2416),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2383),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2356),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2265),
.B(n_1620),
.Y(n_2729)
);

CKINVDCx20_ASAP7_75t_R g2730 ( 
.A(n_2361),
.Y(n_2730)
);

NAND2xp33_ASAP7_75t_L g2731 ( 
.A(n_2281),
.B(n_1244),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_L g2732 ( 
.A(n_2398),
.B(n_1324),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2487),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2446),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2356),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2422),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2402),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2402),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2332),
.B(n_1333),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2422),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_R g2741 ( 
.A(n_2202),
.B(n_2370),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2367),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2412),
.B(n_1334),
.Y(n_2743)
);

AND2x2_ASAP7_75t_SL g2744 ( 
.A(n_2301),
.B(n_2246),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2283),
.B(n_2290),
.Y(n_2745)
);

BUFx6f_ASAP7_75t_L g2746 ( 
.A(n_2392),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2402),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2345),
.B(n_1336),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2457),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2372),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2392),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2287),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2345),
.B(n_1342),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2417),
.B(n_1343),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2254),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2418),
.B(n_1345),
.Y(n_2756)
);

INVx4_ASAP7_75t_L g2757 ( 
.A(n_2375),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_SL g2758 ( 
.A(n_2291),
.B(n_1352),
.Y(n_2758)
);

BUFx2_ASAP7_75t_L g2759 ( 
.A(n_2308),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2377),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2419),
.B(n_1356),
.Y(n_2761)
);

NAND2xp33_ASAP7_75t_SL g2762 ( 
.A(n_2274),
.B(n_1359),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2302),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2420),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2428),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2268),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_L g2767 ( 
.A(n_2310),
.B(n_1361),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2272),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2429),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2275),
.B(n_1362),
.Y(n_2770)
);

OR2x2_ASAP7_75t_L g2771 ( 
.A(n_2242),
.B(n_1641),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2270),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2430),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2264),
.B(n_1364),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2285),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_R g2776 ( 
.A(n_2262),
.B(n_2232),
.Y(n_2776)
);

OR2x2_ASAP7_75t_L g2777 ( 
.A(n_2234),
.B(n_1643),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2322),
.Y(n_2778)
);

INVx3_ASAP7_75t_L g2779 ( 
.A(n_2378),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2410),
.B(n_1365),
.Y(n_2780)
);

INVx1_ASAP7_75t_SL g2781 ( 
.A(n_2381),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2328),
.Y(n_2782)
);

NAND2x1p5_ASAP7_75t_L g2783 ( 
.A(n_2388),
.B(n_1714),
.Y(n_2783)
);

OAI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2253),
.A2(n_1373),
.B1(n_1375),
.B2(n_1371),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2228),
.B(n_1376),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2258),
.B(n_1327),
.Y(n_2786)
);

INVxp67_ASAP7_75t_SL g2787 ( 
.A(n_2241),
.Y(n_2787)
);

AO21x2_ASAP7_75t_L g2788 ( 
.A1(n_2331),
.A2(n_1251),
.B(n_1250),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2333),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2318),
.B(n_1377),
.Y(n_2790)
);

CKINVDCx20_ASAP7_75t_R g2791 ( 
.A(n_2390),
.Y(n_2791)
);

INVx2_ASAP7_75t_SL g2792 ( 
.A(n_2396),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2320),
.B(n_1382),
.Y(n_2793)
);

BUFx4f_ASAP7_75t_L g2794 ( 
.A(n_2340),
.Y(n_2794)
);

INVx2_ASAP7_75t_SL g2795 ( 
.A(n_2400),
.Y(n_2795)
);

BUFx2_ASAP7_75t_L g2796 ( 
.A(n_2279),
.Y(n_2796)
);

INVx3_ASAP7_75t_L g2797 ( 
.A(n_2260),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2343),
.Y(n_2798)
);

INVx4_ASAP7_75t_SL g2799 ( 
.A(n_2350),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2324),
.B(n_1327),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2277),
.B(n_1385),
.Y(n_2801)
);

BUFx10_ASAP7_75t_L g2802 ( 
.A(n_2280),
.Y(n_2802)
);

INVxp33_ASAP7_75t_L g2803 ( 
.A(n_2292),
.Y(n_2803)
);

OR2x6_ASAP7_75t_L g2804 ( 
.A(n_2206),
.B(n_1157),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2352),
.B(n_1386),
.Y(n_2805)
);

NAND2x1p5_ASAP7_75t_L g2806 ( 
.A(n_2357),
.B(n_1256),
.Y(n_2806)
);

AND2x4_ASAP7_75t_L g2807 ( 
.A(n_2222),
.B(n_1389),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2362),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2230),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2363),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2305),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2364),
.B(n_1394),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2311),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2315),
.B(n_1399),
.Y(n_2814)
);

AND2x2_ASAP7_75t_SL g2815 ( 
.A(n_2260),
.B(n_1170),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_SL g2816 ( 
.A(n_2327),
.B(n_1400),
.Y(n_2816)
);

AOI22xp33_ASAP7_75t_L g2817 ( 
.A1(n_2359),
.A2(n_1406),
.B1(n_1464),
.B2(n_1335),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2344),
.B(n_1403),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2358),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2313),
.B(n_1405),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2449),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2313),
.B(n_1407),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2443),
.Y(n_2823)
);

BUFx2_ASAP7_75t_L g2824 ( 
.A(n_2465),
.Y(n_2824)
);

BUFx10_ASAP7_75t_L g2825 ( 
.A(n_2203),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2261),
.B(n_1408),
.Y(n_2826)
);

BUFx6f_ASAP7_75t_L g2827 ( 
.A(n_2192),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2461),
.B(n_1335),
.Y(n_2828)
);

INVx2_ASAP7_75t_SL g2829 ( 
.A(n_2479),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2443),
.Y(n_2830)
);

NAND2xp33_ASAP7_75t_L g2831 ( 
.A(n_2281),
.B(n_1244),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2443),
.Y(n_2832)
);

INVx4_ASAP7_75t_L g2833 ( 
.A(n_2183),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2261),
.B(n_1409),
.Y(n_2834)
);

INVxp33_ASAP7_75t_L g2835 ( 
.A(n_2461),
.Y(n_2835)
);

NAND2xp33_ASAP7_75t_L g2836 ( 
.A(n_2281),
.B(n_1244),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_2465),
.Y(n_2837)
);

BUFx10_ASAP7_75t_L g2838 ( 
.A(n_2203),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2449),
.Y(n_2839)
);

AND2x6_ASAP7_75t_L g2840 ( 
.A(n_2443),
.B(n_1369),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2473),
.B(n_1410),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2449),
.Y(n_2842)
);

AND2x6_ASAP7_75t_L g2843 ( 
.A(n_2443),
.B(n_1369),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2449),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2479),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_SL g2846 ( 
.A(n_2426),
.B(n_1411),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2443),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2449),
.Y(n_2848)
);

AND2x4_ASAP7_75t_L g2849 ( 
.A(n_2465),
.B(n_1412),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_2192),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2449),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2313),
.B(n_1415),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2443),
.Y(n_2853)
);

CKINVDCx16_ASAP7_75t_R g2854 ( 
.A(n_2217),
.Y(n_2854)
);

BUFx2_ASAP7_75t_L g2855 ( 
.A(n_2465),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2313),
.B(n_1418),
.Y(n_2856)
);

NAND2x1p5_ASAP7_75t_L g2857 ( 
.A(n_2473),
.B(n_1258),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2313),
.A2(n_1433),
.B1(n_1436),
.B2(n_1427),
.Y(n_2858)
);

OR2x2_ASAP7_75t_L g2859 ( 
.A(n_2473),
.B(n_1437),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2261),
.B(n_1440),
.Y(n_2860)
);

AND2x4_ASAP7_75t_L g2861 ( 
.A(n_2465),
.B(n_1441),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2465),
.Y(n_2862)
);

BUFx2_ASAP7_75t_L g2863 ( 
.A(n_2465),
.Y(n_2863)
);

INVxp67_ASAP7_75t_L g2864 ( 
.A(n_2461),
.Y(n_2864)
);

INVx4_ASAP7_75t_L g2865 ( 
.A(n_2183),
.Y(n_2865)
);

AND2x4_ASAP7_75t_L g2866 ( 
.A(n_2465),
.B(n_1442),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2313),
.B(n_1443),
.Y(n_2867)
);

INVx1_ASAP7_75t_SL g2868 ( 
.A(n_2465),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2465),
.Y(n_2869)
);

INVx1_ASAP7_75t_SL g2870 ( 
.A(n_2465),
.Y(n_2870)
);

AOI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2233),
.A2(n_1406),
.B1(n_1464),
.B2(n_1335),
.Y(n_2871)
);

INVxp67_ASAP7_75t_SL g2872 ( 
.A(n_2461),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2465),
.B(n_1449),
.Y(n_2873)
);

INVxp33_ASAP7_75t_L g2874 ( 
.A(n_2461),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2465),
.Y(n_2875)
);

AOI22xp33_ASAP7_75t_L g2876 ( 
.A1(n_2233),
.A2(n_1464),
.B1(n_1485),
.B2(n_1406),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2461),
.B(n_1485),
.Y(n_2877)
);

INVx1_ASAP7_75t_SL g2878 ( 
.A(n_2465),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2443),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2449),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2313),
.B(n_1452),
.Y(n_2881)
);

BUFx6f_ASAP7_75t_L g2882 ( 
.A(n_2192),
.Y(n_2882)
);

INVx3_ASAP7_75t_L g2883 ( 
.A(n_2479),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2443),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2513),
.B(n_1453),
.Y(n_2885)
);

INVx2_ASAP7_75t_SL g2886 ( 
.A(n_2517),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2585),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2857),
.B(n_1456),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2576),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2526),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2530),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2522),
.B(n_1457),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_SL g2893 ( 
.A(n_2523),
.B(n_1463),
.Y(n_2893)
);

OAI22xp5_ASAP7_75t_L g2894 ( 
.A1(n_2565),
.A2(n_1225),
.B1(n_1237),
.B2(n_1170),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_SL g2895 ( 
.A(n_2864),
.B(n_2512),
.Y(n_2895)
);

INVx4_ASAP7_75t_L g2896 ( 
.A(n_2517),
.Y(n_2896)
);

INVx1_ASAP7_75t_SL g2897 ( 
.A(n_2868),
.Y(n_2897)
);

NOR2x1_ASAP7_75t_L g2898 ( 
.A(n_2492),
.B(n_1262),
.Y(n_2898)
);

NOR3xp33_ASAP7_75t_L g2899 ( 
.A(n_2507),
.B(n_1269),
.C(n_1265),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2524),
.B(n_1465),
.Y(n_2900)
);

OR2x6_ASAP7_75t_L g2901 ( 
.A(n_2833),
.B(n_1225),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2525),
.B(n_1466),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2535),
.B(n_2543),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2520),
.A2(n_2531),
.B1(n_2593),
.B2(n_2570),
.Y(n_2904)
);

NAND2xp33_ASAP7_75t_L g2905 ( 
.A(n_2840),
.B(n_1469),
.Y(n_2905)
);

OAI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2728),
.A2(n_1246),
.B1(n_1261),
.B2(n_1237),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2545),
.B(n_1470),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2591),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2549),
.B(n_1473),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2551),
.B(n_1477),
.Y(n_2910)
);

BUFx6f_ASAP7_75t_L g2911 ( 
.A(n_2528),
.Y(n_2911)
);

BUFx3_ASAP7_75t_L g2912 ( 
.A(n_2527),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_SL g2913 ( 
.A(n_2511),
.B(n_1483),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_2829),
.B(n_1484),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2572),
.B(n_1489),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2589),
.B(n_1490),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2562),
.B(n_1492),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2527),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2567),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2571),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2827),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2580),
.B(n_1493),
.Y(n_2922)
);

HB1xp67_ASAP7_75t_L g2923 ( 
.A(n_2496),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_SL g2924 ( 
.A(n_2497),
.B(n_1495),
.Y(n_2924)
);

AND2x6_ASAP7_75t_SL g2925 ( 
.A(n_2495),
.B(n_1276),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2845),
.B(n_1496),
.Y(n_2926)
);

INVxp67_ASAP7_75t_L g2927 ( 
.A(n_2824),
.Y(n_2927)
);

BUFx8_ASAP7_75t_L g2928 ( 
.A(n_2824),
.Y(n_2928)
);

NOR2xp67_ASAP7_75t_L g2929 ( 
.A(n_2865),
.B(n_245),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2491),
.Y(n_2930)
);

A2O1A1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2702),
.A2(n_1261),
.B(n_1332),
.C(n_1246),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_SL g2932 ( 
.A(n_2883),
.B(n_1500),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2835),
.B(n_1502),
.Y(n_2933)
);

NAND2xp33_ASAP7_75t_L g2934 ( 
.A(n_2840),
.B(n_1503),
.Y(n_2934)
);

OR2x6_ASAP7_75t_L g2935 ( 
.A(n_2579),
.B(n_1332),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2538),
.A2(n_1520),
.B1(n_1532),
.B2(n_1504),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2821),
.Y(n_2937)
);

HB1xp67_ASAP7_75t_L g2938 ( 
.A(n_2837),
.Y(n_2938)
);

INVx1_ASAP7_75t_SL g2939 ( 
.A(n_2870),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2582),
.A2(n_1485),
.B1(n_1561),
.B2(n_1494),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_2874),
.B(n_1534),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2494),
.B(n_1494),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2839),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2842),
.B(n_2844),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2848),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2598),
.B(n_1541),
.Y(n_2946)
);

INVx2_ASAP7_75t_SL g2947 ( 
.A(n_2827),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2851),
.B(n_1542),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2850),
.B(n_1543),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2600),
.B(n_1545),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2880),
.B(n_1546),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2564),
.B(n_1548),
.Y(n_2952)
);

INVxp67_ASAP7_75t_L g2953 ( 
.A(n_2855),
.Y(n_2953)
);

OAI221xp5_ASAP7_75t_L g2954 ( 
.A1(n_2521),
.A2(n_2550),
.B1(n_2500),
.B2(n_2505),
.C(n_2771),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2872),
.B(n_1551),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2841),
.B(n_1553),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2777),
.B(n_1554),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2859),
.B(n_2610),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2706),
.B(n_1555),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2508),
.B(n_2820),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_L g2961 ( 
.A(n_2499),
.B(n_2605),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2587),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2592),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2786),
.B(n_1494),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2822),
.B(n_1558),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2850),
.B(n_1560),
.Y(n_2966)
);

A2O1A1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2703),
.A2(n_1363),
.B(n_1383),
.C(n_1358),
.Y(n_2967)
);

NOR2xp67_ASAP7_75t_L g2968 ( 
.A(n_2552),
.B(n_245),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2852),
.B(n_1563),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2856),
.B(n_1566),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2697),
.Y(n_2971)
);

NOR2x1p5_ASAP7_75t_L g2972 ( 
.A(n_2862),
.B(n_1571),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2867),
.B(n_1572),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2881),
.B(n_2548),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2858),
.B(n_1574),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_2514),
.B(n_1577),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2595),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2575),
.B(n_1586),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2704),
.Y(n_2979)
);

HB1xp67_ASAP7_75t_L g2980 ( 
.A(n_2869),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2597),
.B(n_1588),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2604),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2540),
.B(n_1278),
.Y(n_2983)
);

BUFx6f_ASAP7_75t_L g2984 ( 
.A(n_2528),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2534),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2828),
.B(n_1590),
.Y(n_2986)
);

NAND3xp33_ASAP7_75t_L g2987 ( 
.A(n_2655),
.B(n_1595),
.C(n_1591),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2733),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2882),
.B(n_1597),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2607),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2611),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2670),
.Y(n_2992)
);

INVx2_ASAP7_75t_SL g2993 ( 
.A(n_2882),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2877),
.B(n_1601),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2622),
.B(n_1603),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2612),
.A2(n_1604),
.B1(n_1606),
.B2(n_1605),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2826),
.B(n_1608),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2639),
.B(n_1610),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2641),
.B(n_1611),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2621),
.B(n_1616),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2620),
.Y(n_3001)
);

O2A1O1Ixp33_ASAP7_75t_L g3002 ( 
.A1(n_2583),
.A2(n_1280),
.B(n_1281),
.C(n_1279),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2834),
.B(n_1617),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2648),
.B(n_2684),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2768),
.B(n_1618),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2717),
.B(n_1622),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_2510),
.A2(n_1732),
.B1(n_1783),
.B2(n_1561),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2685),
.Y(n_3008)
);

A2O1A1Ixp33_ASAP7_75t_L g3009 ( 
.A1(n_2705),
.A2(n_1363),
.B(n_1383),
.C(n_1358),
.Y(n_3009)
);

NOR2xp33_ASAP7_75t_L g3010 ( 
.A(n_2860),
.B(n_1624),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2631),
.Y(n_3011)
);

AOI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2643),
.A2(n_1627),
.B1(n_1632),
.B2(n_1628),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2729),
.B(n_1633),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_SL g3014 ( 
.A(n_2665),
.B(n_1634),
.Y(n_3014)
);

INVx8_ASAP7_75t_L g3015 ( 
.A(n_2840),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_SL g3016 ( 
.A(n_2665),
.B(n_1638),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2657),
.B(n_1640),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2699),
.B(n_1645),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2718),
.B(n_1649),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2635),
.Y(n_3020)
);

AOI22x1_ASAP7_75t_SL g3021 ( 
.A1(n_2730),
.A2(n_1652),
.B1(n_1653),
.B2(n_1651),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_2529),
.B(n_1655),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2647),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2659),
.Y(n_3024)
);

OAI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2735),
.A2(n_1285),
.B(n_1283),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2619),
.B(n_1656),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2660),
.Y(n_3027)
);

INVx2_ASAP7_75t_SL g3028 ( 
.A(n_2579),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2804),
.B(n_1561),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2663),
.B(n_1657),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2785),
.B(n_1659),
.Y(n_3031)
);

OR2x6_ASAP7_75t_L g3032 ( 
.A(n_2783),
.B(n_1417),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2671),
.Y(n_3033)
);

AND2x4_ASAP7_75t_SL g3034 ( 
.A(n_2791),
.B(n_1732),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2676),
.B(n_2678),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2682),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2689),
.Y(n_3037)
);

INVxp67_ASAP7_75t_L g3038 ( 
.A(n_2855),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_SL g3039 ( 
.A(n_2626),
.B(n_1732),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2784),
.B(n_1660),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2664),
.B(n_1665),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2753),
.B(n_1666),
.Y(n_3042)
);

OAI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_2736),
.A2(n_2740),
.B1(n_2751),
.B2(n_2746),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2614),
.B(n_1668),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2680),
.B(n_1670),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2691),
.Y(n_3046)
);

CKINVDCx5p33_ASAP7_75t_R g3047 ( 
.A(n_2596),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_L g3048 ( 
.A1(n_2510),
.A2(n_1783),
.B1(n_1672),
.B2(n_1673),
.Y(n_3048)
);

OR2x2_ASAP7_75t_L g3049 ( 
.A(n_2878),
.B(n_2506),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2714),
.B(n_1671),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_2623),
.B(n_1674),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2693),
.B(n_1678),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2710),
.B(n_1683),
.Y(n_3053)
);

AOI22xp33_ASAP7_75t_L g3054 ( 
.A1(n_2744),
.A2(n_1783),
.B1(n_1688),
.B2(n_1691),
.Y(n_3054)
);

INVxp67_ASAP7_75t_L g3055 ( 
.A(n_2863),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2713),
.B(n_1686),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2673),
.B(n_1692),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2732),
.B(n_1693),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2519),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2743),
.B(n_1694),
.Y(n_3060)
);

HB1xp67_ASAP7_75t_L g3061 ( 
.A(n_2501),
.Y(n_3061)
);

NOR2xp33_ASAP7_75t_L g3062 ( 
.A(n_2749),
.B(n_1695),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2533),
.B(n_2815),
.Y(n_3063)
);

NOR2xp33_ASAP7_75t_L g3064 ( 
.A(n_2764),
.B(n_1696),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2539),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2814),
.B(n_1698),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2632),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2533),
.B(n_1701),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2654),
.B(n_1703),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2606),
.B(n_1704),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2613),
.B(n_2694),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2711),
.B(n_1710),
.Y(n_3072)
);

AOI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_2577),
.A2(n_1712),
.B1(n_1715),
.B2(n_1711),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2765),
.B(n_1717),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2633),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2642),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2644),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2541),
.Y(n_3078)
);

A2O1A1Ixp33_ASAP7_75t_L g3079 ( 
.A1(n_2493),
.A2(n_1461),
.B(n_1479),
.C(n_1417),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2668),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2806),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2503),
.B(n_1719),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2504),
.B(n_1720),
.Y(n_3083)
);

CKINVDCx11_ASAP7_75t_R g3084 ( 
.A(n_2617),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2586),
.A2(n_1289),
.B(n_1286),
.Y(n_3085)
);

NAND2xp33_ASAP7_75t_SL g3086 ( 
.A(n_2741),
.B(n_2776),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2769),
.B(n_1723),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2804),
.B(n_1725),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2773),
.B(n_1735),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2561),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2515),
.B(n_2518),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2818),
.Y(n_3092)
);

OAI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2854),
.A2(n_1743),
.B1(n_1744),
.B2(n_1736),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2800),
.B(n_1748),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2540),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2719),
.B(n_1749),
.Y(n_3096)
);

BUFx8_ASAP7_75t_L g3097 ( 
.A(n_2863),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2627),
.B(n_1750),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2746),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2805),
.Y(n_3100)
);

NAND2xp33_ASAP7_75t_L g3101 ( 
.A(n_2843),
.B(n_1751),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_SL g3102 ( 
.A(n_2584),
.B(n_1753),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2875),
.B(n_1758),
.Y(n_3103)
);

AND2x4_ASAP7_75t_L g3104 ( 
.A(n_2584),
.B(n_1293),
.Y(n_3104)
);

INVx2_ASAP7_75t_SL g3105 ( 
.A(n_2542),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2609),
.B(n_1759),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2812),
.Y(n_3107)
);

CKINVDCx5p33_ASAP7_75t_R g3108 ( 
.A(n_2825),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2751),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2752),
.Y(n_3110)
);

INVxp67_ASAP7_75t_L g3111 ( 
.A(n_2875),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2722),
.A2(n_1766),
.B1(n_1767),
.B2(n_1765),
.Y(n_3112)
);

INVx2_ASAP7_75t_SL g3113 ( 
.A(n_2838),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2712),
.Y(n_3114)
);

INVx4_ASAP7_75t_L g3115 ( 
.A(n_2584),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2849),
.B(n_1771),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2701),
.Y(n_3117)
);

NAND2xp33_ASAP7_75t_L g3118 ( 
.A(n_2843),
.B(n_1774),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2602),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2581),
.B(n_1775),
.Y(n_3120)
);

INVxp67_ASAP7_75t_L g3121 ( 
.A(n_2861),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2554),
.B(n_1784),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2866),
.B(n_1789),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_2873),
.A2(n_1795),
.B1(n_1791),
.B2(n_1491),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2636),
.B(n_1295),
.Y(n_3125)
);

AOI221xp5_ASAP7_75t_L g3126 ( 
.A1(n_2560),
.A2(n_1311),
.B1(n_1315),
.B2(n_1304),
.C(n_1296),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2645),
.B(n_1323),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2649),
.B(n_1326),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2666),
.B(n_1328),
.Y(n_3129)
);

AOI22xp33_ASAP7_75t_L g3130 ( 
.A1(n_2809),
.A2(n_1491),
.B1(n_1570),
.B2(n_1458),
.Y(n_3130)
);

BUFx3_ASAP7_75t_L g3131 ( 
.A(n_2637),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2502),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2628),
.B(n_1329),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2498),
.B(n_1330),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2846),
.B(n_1331),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2708),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2871),
.B(n_2876),
.Y(n_3137)
);

BUFx3_ASAP7_75t_L g3138 ( 
.A(n_2724),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2690),
.B(n_1340),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2754),
.B(n_1344),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2726),
.B(n_1257),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2756),
.B(n_1348),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_SL g3143 ( 
.A(n_2763),
.B(n_1257),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2767),
.B(n_1354),
.Y(n_3144)
);

NAND3xp33_ASAP7_75t_L g3145 ( 
.A(n_2721),
.B(n_1380),
.C(n_1369),
.Y(n_3145)
);

INVxp67_ASAP7_75t_R g3146 ( 
.A(n_2688),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2761),
.B(n_1355),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_L g3148 ( 
.A(n_2608),
.B(n_1357),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2672),
.B(n_1366),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2650),
.B(n_1257),
.Y(n_3150)
);

NAND2x1p5_ASAP7_75t_L g3151 ( 
.A(n_2534),
.B(n_1380),
.Y(n_3151)
);

INVx2_ASAP7_75t_SL g3152 ( 
.A(n_2750),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2739),
.B(n_1381),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2675),
.B(n_1388),
.Y(n_3154)
);

OR2x6_ASAP7_75t_L g3155 ( 
.A(n_2555),
.B(n_1461),
.Y(n_3155)
);

AOI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2537),
.A2(n_1395),
.B1(n_1396),
.B2(n_1392),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2630),
.B(n_2780),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2630),
.B(n_1397),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2630),
.B(n_1401),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2823),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2809),
.A2(n_1491),
.B1(n_1570),
.B2(n_1458),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2790),
.B(n_1404),
.Y(n_3162)
);

INVx4_ASAP7_75t_L g3163 ( 
.A(n_2700),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2793),
.B(n_1416),
.Y(n_3164)
);

INVx4_ASAP7_75t_L g3165 ( 
.A(n_2843),
.Y(n_3165)
);

INVx8_ASAP7_75t_L g3166 ( 
.A(n_2716),
.Y(n_3166)
);

AOI22xp33_ASAP7_75t_L g3167 ( 
.A1(n_2807),
.A2(n_1491),
.B1(n_1570),
.B2(n_1458),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2801),
.B(n_1419),
.Y(n_3168)
);

INVx5_ASAP7_75t_L g3169 ( 
.A(n_2716),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2692),
.Y(n_3170)
);

INVx8_ASAP7_75t_L g3171 ( 
.A(n_2716),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2696),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2884),
.B(n_2830),
.Y(n_3173)
);

HB1xp67_ASAP7_75t_L g3174 ( 
.A(n_2532),
.Y(n_3174)
);

INVx3_ASAP7_75t_L g3175 ( 
.A(n_2566),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2832),
.B(n_1420),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2879),
.B(n_1421),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2847),
.B(n_1426),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_SL g3179 ( 
.A(n_2544),
.B(n_1257),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2679),
.B(n_1428),
.Y(n_3180)
);

OR2x2_ASAP7_75t_L g3181 ( 
.A(n_2509),
.B(n_1429),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_2546),
.B(n_1430),
.Y(n_3182)
);

NOR3xp33_ASAP7_75t_L g3183 ( 
.A(n_2616),
.B(n_1801),
.C(n_1800),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2638),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2778),
.Y(n_3185)
);

NOR2x1p5_ASAP7_75t_L g3186 ( 
.A(n_2698),
.B(n_1439),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_2787),
.B(n_1447),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2687),
.B(n_1450),
.Y(n_3188)
);

BUFx6f_ASAP7_75t_L g3189 ( 
.A(n_2566),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2782),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2853),
.Y(n_3191)
);

NOR2x2_ASAP7_75t_L g3192 ( 
.A(n_2599),
.B(n_1479),
.Y(n_3192)
);

AOI22xp33_ASAP7_75t_L g3193 ( 
.A1(n_2796),
.A2(n_2559),
.B1(n_2624),
.B2(n_2569),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2817),
.B(n_1460),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_2734),
.A2(n_1467),
.B(n_1462),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2788),
.B(n_2742),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2590),
.Y(n_3197)
);

INVx8_ASAP7_75t_L g3198 ( 
.A(n_2723),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2789),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_SL g3200 ( 
.A(n_2686),
.B(n_1267),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2798),
.A2(n_1474),
.B(n_1472),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2624),
.B(n_1267),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2590),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2774),
.B(n_1487),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2588),
.B(n_1488),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2634),
.B(n_1498),
.Y(n_3206)
);

OR2x2_ASAP7_75t_L g3207 ( 
.A(n_2578),
.B(n_1507),
.Y(n_3207)
);

NOR2xp67_ASAP7_75t_SL g3208 ( 
.A(n_2556),
.B(n_2674),
.Y(n_3208)
);

INVx2_ASAP7_75t_SL g3209 ( 
.A(n_2709),
.Y(n_3209)
);

OR2x2_ASAP7_75t_L g3210 ( 
.A(n_2547),
.B(n_1510),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2563),
.B(n_1267),
.Y(n_3211)
);

AOI22xp5_ASAP7_75t_L g3212 ( 
.A1(n_2640),
.A2(n_1521),
.B1(n_1528),
.B2(n_1517),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2808),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2662),
.B(n_1529),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2794),
.B(n_1267),
.Y(n_3215)
);

NAND2x1_ASAP7_75t_L g3216 ( 
.A(n_2723),
.B(n_1380),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2810),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_SL g3218 ( 
.A(n_2601),
.B(n_1270),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2677),
.B(n_1531),
.Y(n_3219)
);

AOI22xp33_ASAP7_75t_L g3220 ( 
.A1(n_2796),
.A2(n_1491),
.B1(n_1570),
.B2(n_1458),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2681),
.B(n_1544),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_2601),
.B(n_1270),
.Y(n_3222)
);

AND2x6_ASAP7_75t_SL g3223 ( 
.A(n_2603),
.B(n_1547),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2615),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2748),
.B(n_1549),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_2615),
.B(n_1270),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2625),
.B(n_1270),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2625),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_2651),
.B(n_1316),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2816),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2720),
.B(n_2536),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_L g3232 ( 
.A1(n_2759),
.A2(n_2762),
.B1(n_2795),
.B2(n_2792),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_SL g3233 ( 
.A(n_2651),
.B(n_1316),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2813),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_SL g3235 ( 
.A(n_2658),
.B(n_1316),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_2658),
.B(n_2661),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2661),
.Y(n_3237)
);

OAI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_2646),
.A2(n_1573),
.B1(n_1575),
.B2(n_1550),
.Y(n_3238)
);

AND2x4_ASAP7_75t_L g3239 ( 
.A(n_2799),
.B(n_1578),
.Y(n_3239)
);

BUFx6f_ASAP7_75t_L g3240 ( 
.A(n_2683),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2573),
.B(n_1583),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2683),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2758),
.B(n_1585),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2770),
.B(n_1589),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2759),
.A2(n_1593),
.B1(n_1594),
.B2(n_1592),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_2695),
.B(n_1316),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2760),
.B(n_1596),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2819),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_2695),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2779),
.B(n_1600),
.Y(n_3250)
);

NAND3xp33_ASAP7_75t_L g3251 ( 
.A(n_2731),
.B(n_1384),
.C(n_1380),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2781),
.B(n_1763),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_2516),
.B(n_1612),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2553),
.B(n_2557),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_2755),
.Y(n_3255)
);

OAI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_2516),
.A2(n_1516),
.B1(n_1518),
.B2(n_1497),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_2594),
.B(n_1642),
.Y(n_3257)
);

A2O1A1Ixp33_ASAP7_75t_L g3258 ( 
.A1(n_2766),
.A2(n_1516),
.B(n_1518),
.C(n_1497),
.Y(n_3258)
);

AOI22xp5_ASAP7_75t_L g3259 ( 
.A1(n_2669),
.A2(n_1647),
.B1(n_1654),
.B2(n_1644),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_SL g3260 ( 
.A(n_2757),
.B(n_1458),
.Y(n_3260)
);

NAND2xp33_ASAP7_75t_L g3261 ( 
.A(n_2626),
.B(n_1763),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2558),
.B(n_1661),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2715),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2727),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_2574),
.B(n_1664),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2797),
.B(n_2745),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2772),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2723),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2725),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_2802),
.Y(n_3270)
);

NAND2xp33_ASAP7_75t_L g3271 ( 
.A(n_2626),
.B(n_1458),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2803),
.B(n_1669),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2725),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2725),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2629),
.B(n_1675),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_SL g3276 ( 
.A1(n_2618),
.A2(n_1684),
.B1(n_1687),
.B2(n_1677),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2629),
.B(n_1689),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2629),
.B(n_1690),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_SL g3279 ( 
.A(n_2667),
.B(n_1458),
.Y(n_3279)
);

INVx2_ASAP7_75t_SL g3280 ( 
.A(n_2799),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2775),
.Y(n_3281)
);

INVx2_ASAP7_75t_SL g3282 ( 
.A(n_2707),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2737),
.B(n_1699),
.Y(n_3283)
);

O2A1O1Ixp5_ASAP7_75t_L g3284 ( 
.A1(n_2738),
.A2(n_1536),
.B(n_1567),
.C(n_1539),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_SL g3285 ( 
.A(n_2747),
.B(n_1491),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_2811),
.B(n_1491),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2568),
.B(n_1702),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2831),
.B(n_1707),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2652),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2568),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2568),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_2652),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2652),
.B(n_1709),
.Y(n_3293)
);

OR2x2_ASAP7_75t_L g3294 ( 
.A(n_2653),
.B(n_1716),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_2653),
.B(n_1570),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_SL g3296 ( 
.A(n_2653),
.B(n_1570),
.Y(n_3296)
);

NOR2xp33_ASAP7_75t_SL g3297 ( 
.A(n_2656),
.B(n_1570),
.Y(n_3297)
);

NAND2x1p5_ASAP7_75t_L g3298 ( 
.A(n_2656),
.B(n_1384),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2656),
.B(n_1718),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2836),
.B(n_1724),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2513),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_2576),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_2522),
.B(n_1726),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_2513),
.B(n_1763),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_2513),
.B(n_1728),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2513),
.B(n_1730),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_2513),
.B(n_1763),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2513),
.B(n_1763),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2513),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_2576),
.Y(n_3310)
);

AOI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_2507),
.A2(n_1734),
.B1(n_1739),
.B2(n_1738),
.Y(n_3311)
);

AOI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_2507),
.A2(n_1740),
.B1(n_1756),
.B2(n_1752),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_2576),
.Y(n_3313)
);

NOR2xp67_ASAP7_75t_L g3314 ( 
.A(n_2492),
.B(n_245),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_2522),
.B(n_1757),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_2513),
.B(n_1768),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_2522),
.B(n_1777),
.Y(n_3317)
);

INVx2_ASAP7_75t_SL g3318 ( 
.A(n_2517),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_2513),
.Y(n_3319)
);

NAND2xp33_ASAP7_75t_L g3320 ( 
.A(n_2840),
.B(n_1639),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_L g3321 ( 
.A(n_2522),
.B(n_1778),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2576),
.Y(n_3322)
);

BUFx6f_ASAP7_75t_L g3323 ( 
.A(n_2528),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_L g3324 ( 
.A(n_2522),
.B(n_1780),
.Y(n_3324)
);

NOR3xp33_ASAP7_75t_L g3325 ( 
.A(n_2507),
.B(n_1792),
.C(n_1782),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2524),
.B(n_1794),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2513),
.Y(n_3327)
);

NOR3xp33_ASAP7_75t_L g3328 ( 
.A(n_2507),
.B(n_1798),
.C(n_1539),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2524),
.B(n_1639),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2513),
.Y(n_3330)
);

NOR2xp33_ASAP7_75t_L g3331 ( 
.A(n_2522),
.B(n_1536),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_2538),
.A2(n_1763),
.B1(n_1639),
.B2(n_1423),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2513),
.B(n_1639),
.Y(n_3333)
);

AO221x1_ASAP7_75t_L g3334 ( 
.A1(n_2533),
.A2(n_1444),
.B1(n_1423),
.B2(n_1384),
.C(n_1475),
.Y(n_3334)
);

OR2x6_ASAP7_75t_L g3335 ( 
.A(n_2492),
.B(n_1567),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_2517),
.Y(n_3336)
);

BUFx2_ASAP7_75t_L g3337 ( 
.A(n_2496),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_2576),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_2576),
.Y(n_3339)
);

INVx3_ASAP7_75t_L g3340 ( 
.A(n_2517),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_2522),
.B(n_1579),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2513),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_2513),
.B(n_1639),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2513),
.B(n_1639),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_SL g3345 ( 
.A(n_2626),
.B(n_1639),
.Y(n_3345)
);

AND2x2_ASAP7_75t_SL g3346 ( 
.A(n_2532),
.B(n_1579),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2513),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_2513),
.B(n_1763),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_2507),
.A2(n_1761),
.B1(n_1764),
.B2(n_1662),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2513),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_2576),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2513),
.B(n_1662),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2513),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2513),
.B(n_1761),
.Y(n_3354)
);

AOI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_2507),
.A2(n_1764),
.B1(n_1423),
.B2(n_1444),
.Y(n_3355)
);

OR2x2_ASAP7_75t_L g3356 ( 
.A(n_2868),
.B(n_246),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_2513),
.B(n_2),
.Y(n_3357)
);

O2A1O1Ixp5_ASAP7_75t_L g3358 ( 
.A1(n_2687),
.A2(n_1423),
.B(n_1444),
.C(n_1384),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2513),
.B(n_2),
.Y(n_3359)
);

INVx2_ASAP7_75t_SL g3360 ( 
.A(n_2517),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_2522),
.B(n_246),
.Y(n_3361)
);

OR2x6_ASAP7_75t_L g3362 ( 
.A(n_2492),
.B(n_1444),
.Y(n_3362)
);

BUFx6f_ASAP7_75t_L g3363 ( 
.A(n_2528),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2513),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_2522),
.B(n_247),
.Y(n_3365)
);

AND2x6_ASAP7_75t_SL g3366 ( 
.A(n_2495),
.B(n_2),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_2522),
.B(n_247),
.Y(n_3367)
);

OAI221xp5_ASAP7_75t_L g3368 ( 
.A1(n_2521),
.A2(n_1731),
.B1(n_1682),
.B2(n_1475),
.C(n_250),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2513),
.B(n_3),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_2513),
.B(n_1475),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2522),
.B(n_248),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_2538),
.A2(n_1682),
.B1(n_1731),
.B2(n_1475),
.Y(n_3372)
);

INVx2_ASAP7_75t_SL g3373 ( 
.A(n_2517),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2513),
.B(n_3),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_2513),
.B(n_1682),
.Y(n_3375)
);

INVxp67_ASAP7_75t_L g3376 ( 
.A(n_2824),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_2576),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2513),
.B(n_3),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_2513),
.B(n_3),
.Y(n_3379)
);

INVxp67_ASAP7_75t_SL g3380 ( 
.A(n_2513),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_2517),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_2513),
.B(n_1682),
.Y(n_3382)
);

OAI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_2728),
.A2(n_4),
.B(n_5),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_2513),
.B(n_1731),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2513),
.B(n_4),
.Y(n_3385)
);

NOR2xp67_ASAP7_75t_SL g3386 ( 
.A(n_2700),
.B(n_1731),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_2538),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_2513),
.B(n_248),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_2576),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_2522),
.B(n_248),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2513),
.B(n_5),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_L g3392 ( 
.A(n_2522),
.B(n_249),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2576),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_SL g3394 ( 
.A(n_2513),
.B(n_249),
.Y(n_3394)
);

OAI221xp5_ASAP7_75t_L g3395 ( 
.A1(n_2521),
.A2(n_251),
.B1(n_252),
.B2(n_250),
.C(n_249),
.Y(n_3395)
);

O2A1O1Ixp33_ASAP7_75t_L g3396 ( 
.A1(n_2550),
.A2(n_251),
.B(n_252),
.C(n_250),
.Y(n_3396)
);

INVx2_ASAP7_75t_SL g3397 ( 
.A(n_2517),
.Y(n_3397)
);

BUFx3_ASAP7_75t_L g3398 ( 
.A(n_2517),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_2513),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2513),
.B(n_6),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2513),
.B(n_6),
.Y(n_3401)
);

BUFx8_ASAP7_75t_L g3402 ( 
.A(n_2824),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2513),
.B(n_6),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_2522),
.B(n_252),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_SL g3405 ( 
.A(n_2513),
.B(n_253),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_L g3406 ( 
.A(n_2840),
.B(n_7),
.Y(n_3406)
);

INVxp67_ASAP7_75t_L g3407 ( 
.A(n_2824),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2513),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2513),
.B(n_7),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2522),
.B(n_253),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_SL g3411 ( 
.A1(n_2577),
.A2(n_254),
.B1(n_255),
.B2(n_253),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2513),
.B(n_7),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_2576),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2513),
.B(n_8),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_2576),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_SL g3416 ( 
.A(n_2513),
.B(n_254),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_2513),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_2513),
.B(n_255),
.Y(n_3418)
);

OR2x2_ASAP7_75t_L g3419 ( 
.A(n_2868),
.B(n_255),
.Y(n_3419)
);

AOI221xp5_ASAP7_75t_L g3420 ( 
.A1(n_2550),
.A2(n_258),
.B1(n_259),
.B2(n_257),
.C(n_256),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2513),
.B(n_8),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2513),
.Y(n_3422)
);

BUFx2_ASAP7_75t_L g3423 ( 
.A(n_2496),
.Y(n_3423)
);

O2A1O1Ixp33_ASAP7_75t_L g3424 ( 
.A1(n_2550),
.A2(n_257),
.B(n_258),
.C(n_256),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2513),
.B(n_8),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2576),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2513),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2513),
.Y(n_3428)
);

OR2x2_ASAP7_75t_L g3429 ( 
.A(n_2868),
.B(n_256),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_2522),
.B(n_257),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_2522),
.B(n_258),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_2522),
.B(n_259),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_2513),
.B(n_8),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_2522),
.B(n_259),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2513),
.Y(n_3435)
);

NOR2x1p5_ASAP7_75t_L g3436 ( 
.A(n_2496),
.B(n_260),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_2513),
.B(n_260),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2576),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_2513),
.B(n_260),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2513),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2513),
.B(n_9),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2513),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2513),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2513),
.B(n_9),
.Y(n_3444)
);

BUFx6f_ASAP7_75t_L g3445 ( 
.A(n_2528),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_2513),
.B(n_262),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_2513),
.Y(n_3447)
);

OR2x2_ASAP7_75t_L g3448 ( 
.A(n_2868),
.B(n_261),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_2513),
.B(n_10),
.Y(n_3449)
);

NOR3xp33_ASAP7_75t_L g3450 ( 
.A(n_2507),
.B(n_263),
.C(n_262),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2565),
.A2(n_262),
.B1(n_263),
.B2(n_261),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_2513),
.B(n_10),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_L g3453 ( 
.A(n_2522),
.B(n_263),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_2513),
.B(n_264),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_2513),
.B(n_11),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_2513),
.B(n_11),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_2513),
.B(n_264),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_2513),
.B(n_11),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_2507),
.A2(n_266),
.B1(n_267),
.B2(n_265),
.Y(n_3459)
);

NAND2xp33_ASAP7_75t_L g3460 ( 
.A(n_2840),
.B(n_11),
.Y(n_3460)
);

AOI22xp33_ASAP7_75t_L g3461 ( 
.A1(n_2538),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2513),
.B(n_12),
.Y(n_3462)
);

AOI22xp5_ASAP7_75t_L g3463 ( 
.A1(n_2507),
.A2(n_266),
.B1(n_267),
.B2(n_265),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_L g3464 ( 
.A(n_2522),
.B(n_266),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_2513),
.B(n_12),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2513),
.Y(n_3466)
);

AND2x4_ASAP7_75t_L g3467 ( 
.A(n_2523),
.B(n_267),
.Y(n_3467)
);

NOR3xp33_ASAP7_75t_L g3468 ( 
.A(n_2507),
.B(n_269),
.C(n_268),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2513),
.Y(n_3469)
);

AOI22xp33_ASAP7_75t_L g3470 ( 
.A1(n_2538),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_2522),
.B(n_268),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2513),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_2576),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_2513),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_2524),
.B(n_13),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_2576),
.Y(n_3476)
);

AOI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_2507),
.A2(n_270),
.B1(n_271),
.B2(n_269),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_2524),
.B(n_13),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_2524),
.B(n_14),
.Y(n_3479)
);

INVx2_ASAP7_75t_SL g3480 ( 
.A(n_2517),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2513),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_2513),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_2524),
.B(n_14),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_2524),
.B(n_15),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_2524),
.B(n_15),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_2522),
.B(n_269),
.Y(n_3486)
);

NOR2xp33_ASAP7_75t_L g3487 ( 
.A(n_2522),
.B(n_270),
.Y(n_3487)
);

AOI22xp5_ASAP7_75t_L g3488 ( 
.A1(n_2507),
.A2(n_272),
.B1(n_273),
.B2(n_271),
.Y(n_3488)
);

AOI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_2507),
.A2(n_272),
.B1(n_273),
.B2(n_271),
.Y(n_3489)
);

NOR2xp33_ASAP7_75t_L g3490 ( 
.A(n_2522),
.B(n_272),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_2524),
.B(n_16),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_2524),
.B(n_16),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_2576),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_2513),
.B(n_274),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_2524),
.B(n_16),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_2513),
.B(n_274),
.Y(n_3496)
);

XNOR2xp5_ASAP7_75t_L g3497 ( 
.A(n_2609),
.B(n_16),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_SL g3498 ( 
.A(n_2513),
.B(n_274),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_2524),
.B(n_17),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_2513),
.Y(n_3500)
);

BUFx3_ASAP7_75t_L g3501 ( 
.A(n_2517),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2524),
.B(n_17),
.Y(n_3502)
);

NAND2xp33_ASAP7_75t_L g3503 ( 
.A(n_2840),
.B(n_17),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_2513),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_2576),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_2857),
.B(n_1121),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_2576),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_2524),
.B(n_17),
.Y(n_3508)
);

O2A1O1Ixp5_ASAP7_75t_L g3509 ( 
.A1(n_2687),
.A2(n_276),
.B(n_277),
.C(n_275),
.Y(n_3509)
);

INVx2_ASAP7_75t_SL g3510 ( 
.A(n_2517),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_2513),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_2524),
.B(n_18),
.Y(n_3512)
);

INVxp67_ASAP7_75t_L g3513 ( 
.A(n_2824),
.Y(n_3513)
);

INVx8_ASAP7_75t_L g3514 ( 
.A(n_2517),
.Y(n_3514)
);

CKINVDCx20_ASAP7_75t_R g3515 ( 
.A(n_2496),
.Y(n_3515)
);

INVx2_ASAP7_75t_SL g3516 ( 
.A(n_2517),
.Y(n_3516)
);

NOR2xp33_ASAP7_75t_L g3517 ( 
.A(n_2522),
.B(n_275),
.Y(n_3517)
);

INVx3_ASAP7_75t_L g3518 ( 
.A(n_2517),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_2524),
.B(n_18),
.Y(n_3519)
);

INVx4_ASAP7_75t_L g3520 ( 
.A(n_2517),
.Y(n_3520)
);

OAI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_2565),
.A2(n_276),
.B1(n_277),
.B2(n_275),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2524),
.B(n_18),
.Y(n_3522)
);

NAND3xp33_ASAP7_75t_L g3523 ( 
.A(n_2655),
.B(n_278),
.C(n_277),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_SL g3524 ( 
.A(n_2626),
.B(n_278),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2524),
.B(n_18),
.Y(n_3525)
);

INVx1_ASAP7_75t_SL g3526 ( 
.A(n_2513),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_2513),
.B(n_19),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_2576),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_2576),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_2576),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_2522),
.B(n_279),
.Y(n_3531)
);

BUFx6f_ASAP7_75t_L g3532 ( 
.A(n_2528),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_2513),
.B(n_279),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_2513),
.B(n_19),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_2576),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2513),
.B(n_19),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_2513),
.B(n_20),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_2576),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_2513),
.B(n_20),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2513),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_SL g3541 ( 
.A(n_2513),
.B(n_279),
.Y(n_3541)
);

NOR2x1p5_ASAP7_75t_L g3542 ( 
.A(n_2496),
.B(n_280),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_2513),
.B(n_20),
.Y(n_3543)
);

AO22x1_ASAP7_75t_L g3544 ( 
.A1(n_2533),
.A2(n_281),
.B1(n_282),
.B2(n_280),
.Y(n_3544)
);

A2O1A1Ixp33_ASAP7_75t_L g3545 ( 
.A1(n_3380),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3545)
);

BUFx6f_ASAP7_75t_L g3546 ( 
.A(n_2911),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3301),
.Y(n_3547)
);

INVxp67_ASAP7_75t_L g3548 ( 
.A(n_3032),
.Y(n_3548)
);

INVxp67_ASAP7_75t_L g3549 ( 
.A(n_3032),
.Y(n_3549)
);

BUFx5_ASAP7_75t_L g3550 ( 
.A(n_3342),
.Y(n_3550)
);

O2A1O1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_2954),
.A2(n_281),
.B(n_282),
.C(n_280),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3039),
.A2(n_284),
.B(n_283),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_SL g3553 ( 
.A(n_3346),
.B(n_3526),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3526),
.B(n_283),
.Y(n_3554)
);

O2A1O1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_2960),
.A2(n_3396),
.B(n_3424),
.C(n_2974),
.Y(n_3555)
);

OAI22xp5_ASAP7_75t_L g3556 ( 
.A1(n_3309),
.A2(n_284),
.B1(n_285),
.B2(n_283),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3319),
.B(n_3327),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_2944),
.Y(n_3558)
);

BUFx6f_ASAP7_75t_L g3559 ( 
.A(n_2911),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3330),
.B(n_285),
.Y(n_3560)
);

OAI21xp33_ASAP7_75t_L g3561 ( 
.A1(n_3144),
.A2(n_21),
.B(n_22),
.Y(n_3561)
);

A2O1A1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_3071),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3562)
);

AOI21xp5_ASAP7_75t_L g3563 ( 
.A1(n_3039),
.A2(n_287),
.B(n_286),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3347),
.B(n_286),
.Y(n_3564)
);

CKINVDCx5p33_ASAP7_75t_R g3565 ( 
.A(n_3084),
.Y(n_3565)
);

INVxp67_ASAP7_75t_L g3566 ( 
.A(n_3032),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3350),
.B(n_286),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3353),
.B(n_287),
.Y(n_3568)
);

O2A1O1Ixp33_ASAP7_75t_SL g3569 ( 
.A1(n_3143),
.A2(n_288),
.B(n_289),
.C(n_287),
.Y(n_3569)
);

A2O1A1Ixp33_ASAP7_75t_L g3570 ( 
.A1(n_3540),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3570)
);

OAI22xp5_ASAP7_75t_L g3571 ( 
.A1(n_3364),
.A2(n_289),
.B1(n_290),
.B2(n_288),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3399),
.B(n_288),
.Y(n_3572)
);

HB1xp67_ASAP7_75t_L g3573 ( 
.A(n_2935),
.Y(n_3573)
);

INVx3_ASAP7_75t_L g3574 ( 
.A(n_3015),
.Y(n_3574)
);

AOI21x1_ASAP7_75t_L g3575 ( 
.A1(n_3043),
.A2(n_291),
.B(n_290),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_2930),
.Y(n_3576)
);

OAI321xp33_ASAP7_75t_L g3577 ( 
.A1(n_3256),
.A2(n_3368),
.A3(n_3395),
.B1(n_3383),
.B2(n_3521),
.C(n_3451),
.Y(n_3577)
);

INVx3_ASAP7_75t_L g3578 ( 
.A(n_3015),
.Y(n_3578)
);

INVx3_ASAP7_75t_L g3579 ( 
.A(n_3015),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3408),
.B(n_291),
.Y(n_3580)
);

AOI21x1_ASAP7_75t_L g3581 ( 
.A1(n_3043),
.A2(n_292),
.B(n_291),
.Y(n_3581)
);

A2O1A1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_3417),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3422),
.B(n_292),
.Y(n_3583)
);

AOI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3345),
.A2(n_293),
.B(n_292),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3427),
.B(n_3428),
.Y(n_3585)
);

NAND2xp33_ASAP7_75t_L g3586 ( 
.A(n_3166),
.B(n_3171),
.Y(n_3586)
);

NAND2xp33_ASAP7_75t_L g3587 ( 
.A(n_3166),
.B(n_293),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3435),
.B(n_3440),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3442),
.B(n_295),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_2911),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_3345),
.A2(n_296),
.B(n_295),
.Y(n_3591)
);

AOI21x1_ASAP7_75t_L g3592 ( 
.A1(n_3196),
.A2(n_296),
.B(n_295),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3443),
.B(n_297),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_3447),
.B(n_297),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3466),
.A2(n_298),
.B1(n_299),
.B2(n_297),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3469),
.B(n_298),
.Y(n_3596)
);

NOR2xp33_ASAP7_75t_L g3597 ( 
.A(n_2904),
.B(n_298),
.Y(n_3597)
);

NOR2xp67_ASAP7_75t_L g3598 ( 
.A(n_2896),
.B(n_299),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3472),
.B(n_299),
.Y(n_3599)
);

CKINVDCx5p33_ASAP7_75t_R g3600 ( 
.A(n_3515),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3474),
.B(n_300),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3481),
.B(n_300),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3482),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3500),
.B(n_301),
.Y(n_3604)
);

BUFx2_ASAP7_75t_L g3605 ( 
.A(n_2935),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3504),
.B(n_301),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_SL g3607 ( 
.A(n_3165),
.B(n_301),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3511),
.Y(n_3608)
);

AND2x4_ASAP7_75t_L g3609 ( 
.A(n_3081),
.B(n_302),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3524),
.B(n_303),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3011),
.Y(n_3611)
);

AOI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_2959),
.A2(n_304),
.B1(n_305),
.B2(n_303),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3020),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3370),
.A2(n_305),
.B(n_304),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3375),
.A2(n_3384),
.B(n_3382),
.Y(n_3615)
);

A2O1A1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_3002),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_3616)
);

O2A1O1Ixp33_ASAP7_75t_L g3617 ( 
.A1(n_3004),
.A2(n_2958),
.B(n_3256),
.C(n_3137),
.Y(n_3617)
);

INVx5_ASAP7_75t_L g3618 ( 
.A(n_3514),
.Y(n_3618)
);

AND2x4_ASAP7_75t_L g3619 ( 
.A(n_2896),
.B(n_305),
.Y(n_3619)
);

BUFx6f_ASAP7_75t_L g3620 ( 
.A(n_2984),
.Y(n_3620)
);

HB1xp67_ASAP7_75t_L g3621 ( 
.A(n_2935),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_2937),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2943),
.Y(n_3623)
);

NAND2x1p5_ASAP7_75t_L g3624 ( 
.A(n_3520),
.B(n_306),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_2903),
.B(n_306),
.Y(n_3625)
);

O2A1O1Ixp5_ASAP7_75t_L g3626 ( 
.A1(n_3388),
.A2(n_308),
.B(n_309),
.C(n_307),
.Y(n_3626)
);

HB1xp67_ASAP7_75t_L g3627 ( 
.A(n_2897),
.Y(n_3627)
);

OAI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_3284),
.A2(n_24),
.B(n_26),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_2903),
.B(n_307),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_3524),
.A2(n_308),
.B(n_307),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_2942),
.B(n_309),
.Y(n_3631)
);

NAND2x1p5_ASAP7_75t_L g3632 ( 
.A(n_3520),
.B(n_309),
.Y(n_3632)
);

INVx1_ASAP7_75t_SL g3633 ( 
.A(n_3514),
.Y(n_3633)
);

OAI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_2907),
.A2(n_24),
.B(n_26),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_2887),
.B(n_310),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_2890),
.B(n_310),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_2891),
.B(n_310),
.Y(n_3637)
);

AOI22xp5_ASAP7_75t_L g3638 ( 
.A1(n_3106),
.A2(n_312),
.B1(n_313),
.B2(n_311),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_2908),
.B(n_311),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_L g3640 ( 
.A(n_3121),
.B(n_311),
.Y(n_3640)
);

AND2x4_ASAP7_75t_L g3641 ( 
.A(n_3100),
.B(n_312),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_3196),
.A2(n_314),
.B(n_313),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_2945),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_2919),
.B(n_313),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3195),
.A2(n_315),
.B(n_314),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_2920),
.B(n_314),
.Y(n_3646)
);

AOI21xp5_ASAP7_75t_L g3647 ( 
.A1(n_3304),
.A2(n_316),
.B(n_315),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2963),
.Y(n_3648)
);

AOI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3307),
.A2(n_316),
.B(n_315),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3107),
.B(n_316),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_R g3651 ( 
.A(n_3108),
.B(n_27),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_2977),
.Y(n_3652)
);

INVxp67_ASAP7_75t_L g3653 ( 
.A(n_3506),
.Y(n_3653)
);

AOI22xp5_ASAP7_75t_L g3654 ( 
.A1(n_2957),
.A2(n_318),
.B1(n_319),
.B2(n_317),
.Y(n_3654)
);

INVx3_ASAP7_75t_L g3655 ( 
.A(n_3165),
.Y(n_3655)
);

INVx4_ASAP7_75t_L g3656 ( 
.A(n_3514),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3166),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3023),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_SL g3659 ( 
.A(n_3093),
.B(n_317),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3305),
.B(n_318),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3306),
.B(n_318),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3025),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_3662)
);

NOR2xp67_ASAP7_75t_L g3663 ( 
.A(n_3163),
.B(n_3115),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3316),
.B(n_319),
.Y(n_3664)
);

INVx3_ASAP7_75t_L g3665 ( 
.A(n_3171),
.Y(n_3665)
);

A2O1A1Ixp33_ASAP7_75t_L g3666 ( 
.A1(n_3025),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_3666)
);

INVx2_ASAP7_75t_SL g3667 ( 
.A(n_2912),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3308),
.A2(n_321),
.B(n_319),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3187),
.B(n_321),
.Y(n_3669)
);

OAI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_2907),
.A2(n_28),
.B(n_29),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_2982),
.B(n_321),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3027),
.Y(n_3672)
);

AND2x6_ASAP7_75t_L g3673 ( 
.A(n_3467),
.B(n_322),
.Y(n_3673)
);

OAI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_2909),
.A2(n_28),
.B(n_29),
.Y(n_3674)
);

CKINVDCx20_ASAP7_75t_R g3675 ( 
.A(n_3034),
.Y(n_3675)
);

OAI321xp33_ASAP7_75t_L g3676 ( 
.A1(n_3383),
.A2(n_31),
.A3(n_33),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_2990),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3033),
.Y(n_3678)
);

INVx1_ASAP7_75t_SL g3679 ( 
.A(n_2897),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3037),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3348),
.A2(n_323),
.B(n_322),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_2991),
.B(n_322),
.Y(n_3682)
);

OAI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_2909),
.A2(n_2917),
.B(n_2910),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3169),
.B(n_323),
.Y(n_3684)
);

AOI21xp5_ASAP7_75t_L g3685 ( 
.A1(n_3286),
.A2(n_324),
.B(n_323),
.Y(n_3685)
);

AOI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_3333),
.A2(n_325),
.B(n_324),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3001),
.Y(n_3687)
);

INVx4_ASAP7_75t_L g3688 ( 
.A(n_3171),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3169),
.B(n_326),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3343),
.A2(n_327),
.B(n_326),
.Y(n_3690)
);

AOI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_3344),
.A2(n_327),
.B(n_326),
.Y(n_3691)
);

OAI21xp33_ASAP7_75t_L g3692 ( 
.A1(n_3044),
.A2(n_30),
.B(n_31),
.Y(n_3692)
);

O2A1O1Ixp5_ASAP7_75t_L g3693 ( 
.A1(n_3394),
.A2(n_328),
.B(n_329),
.C(n_327),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3085),
.A2(n_329),
.B(n_328),
.Y(n_3694)
);

OAI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3259),
.A2(n_330),
.B1(n_331),
.B2(n_328),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3024),
.B(n_330),
.Y(n_3696)
);

O2A1O1Ixp33_ASAP7_75t_L g3697 ( 
.A1(n_3450),
.A2(n_331),
.B(n_332),
.C(n_330),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_2910),
.A2(n_2917),
.B(n_2902),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3157),
.A2(n_3271),
.B(n_3261),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3099),
.A2(n_332),
.B(n_331),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3036),
.B(n_333),
.Y(n_3701)
);

AOI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3109),
.A2(n_334),
.B(n_333),
.Y(n_3702)
);

OAI21xp33_ASAP7_75t_L g3703 ( 
.A1(n_3051),
.A2(n_30),
.B(n_31),
.Y(n_3703)
);

OAI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3467),
.A2(n_335),
.B1(n_336),
.B2(n_334),
.Y(n_3704)
);

AOI22xp5_ASAP7_75t_L g3705 ( 
.A1(n_3088),
.A2(n_335),
.B1(n_336),
.B2(n_334),
.Y(n_3705)
);

INVx1_ASAP7_75t_SL g3706 ( 
.A(n_2939),
.Y(n_3706)
);

AOI21x1_ASAP7_75t_L g3707 ( 
.A1(n_2906),
.A2(n_337),
.B(n_336),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_2964),
.B(n_337),
.Y(n_3708)
);

OR2x2_ASAP7_75t_L g3709 ( 
.A(n_3049),
.B(n_337),
.Y(n_3709)
);

BUFx2_ASAP7_75t_SL g3710 ( 
.A(n_3119),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3046),
.B(n_338),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3092),
.B(n_339),
.Y(n_3712)
);

OAI21xp33_ASAP7_75t_L g3713 ( 
.A1(n_3031),
.A2(n_30),
.B(n_31),
.Y(n_3713)
);

OAI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_2900),
.A2(n_32),
.B(n_33),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3035),
.B(n_339),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3475),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3329),
.A2(n_3285),
.B(n_2934),
.Y(n_3717)
);

OAI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_2900),
.A2(n_32),
.B(n_33),
.Y(n_3718)
);

BUFx8_ASAP7_75t_L g3719 ( 
.A(n_3337),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3329),
.A2(n_340),
.B(n_339),
.Y(n_3720)
);

OR2x2_ASAP7_75t_L g3721 ( 
.A(n_2888),
.B(n_340),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_2984),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_2902),
.B(n_3204),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_L g3724 ( 
.A(n_2927),
.B(n_340),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_2905),
.A2(n_342),
.B(n_341),
.Y(n_3725)
);

AOI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_2946),
.A2(n_342),
.B1(n_343),
.B2(n_341),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3169),
.B(n_341),
.Y(n_3727)
);

OAI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_2922),
.A2(n_32),
.B(n_33),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3151),
.A2(n_344),
.B(n_343),
.Y(n_3729)
);

INVx4_ASAP7_75t_L g3730 ( 
.A(n_3198),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3169),
.B(n_344),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3475),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3101),
.A2(n_346),
.B(n_345),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3204),
.B(n_345),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_2953),
.B(n_345),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_3180),
.B(n_346),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3311),
.B(n_346),
.Y(n_3737)
);

O2A1O1Ixp33_ASAP7_75t_SL g3738 ( 
.A1(n_3179),
.A2(n_348),
.B(n_349),
.C(n_347),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3029),
.B(n_347),
.Y(n_3739)
);

OAI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_2922),
.A2(n_34),
.B(n_35),
.Y(n_3740)
);

OAI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3026),
.A2(n_34),
.B(n_35),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_2889),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_SL g3743 ( 
.A(n_3180),
.B(n_349),
.Y(n_3743)
);

INVx3_ASAP7_75t_L g3744 ( 
.A(n_3198),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3312),
.B(n_350),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3118),
.A2(n_351),
.B(n_350),
.Y(n_3746)
);

OAI321xp33_ASAP7_75t_L g3747 ( 
.A1(n_3451),
.A2(n_36),
.A3(n_38),
.B1(n_34),
.B2(n_35),
.C(n_37),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3406),
.A2(n_352),
.B(n_351),
.Y(n_3748)
);

BUFx6f_ASAP7_75t_L g3749 ( 
.A(n_2984),
.Y(n_3749)
);

BUFx8_ASAP7_75t_SL g3750 ( 
.A(n_3423),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3162),
.B(n_353),
.Y(n_3751)
);

A2O1A1Ixp33_ASAP7_75t_L g3752 ( 
.A1(n_3523),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_3752)
);

O2A1O1Ixp33_ASAP7_75t_SL g3753 ( 
.A1(n_2931),
.A2(n_2967),
.B(n_3009),
.C(n_3079),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3073),
.B(n_354),
.Y(n_3754)
);

CKINVDCx10_ASAP7_75t_R g3755 ( 
.A(n_2901),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3478),
.Y(n_3756)
);

AOI21x1_ASAP7_75t_L g3757 ( 
.A1(n_2906),
.A2(n_356),
.B(n_354),
.Y(n_3757)
);

NOR3xp33_ASAP7_75t_L g3758 ( 
.A(n_3420),
.B(n_3468),
.C(n_3053),
.Y(n_3758)
);

O2A1O1Ixp33_ASAP7_75t_L g3759 ( 
.A1(n_3238),
.A2(n_3069),
.B(n_3325),
.C(n_2899),
.Y(n_3759)
);

AOI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_2950),
.A2(n_356),
.B1(n_357),
.B2(n_354),
.Y(n_3760)
);

AO21x1_ASAP7_75t_L g3761 ( 
.A1(n_3460),
.A2(n_358),
.B(n_357),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_2939),
.B(n_357),
.Y(n_3762)
);

O2A1O1Ixp33_ASAP7_75t_L g3763 ( 
.A1(n_2956),
.A2(n_359),
.B(n_360),
.C(n_358),
.Y(n_3763)
);

AOI21xp5_ASAP7_75t_L g3764 ( 
.A1(n_3503),
.A2(n_360),
.B(n_359),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3478),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3479),
.Y(n_3766)
);

CKINVDCx20_ASAP7_75t_R g3767 ( 
.A(n_2928),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3302),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3038),
.B(n_359),
.Y(n_3769)
);

OAI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3072),
.A2(n_36),
.B(n_37),
.Y(n_3770)
);

OAI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3362),
.A2(n_362),
.B1(n_363),
.B2(n_361),
.Y(n_3771)
);

A2O1A1Ixp33_ASAP7_75t_L g3772 ( 
.A1(n_3509),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_3772)
);

BUFx6f_ASAP7_75t_L g3773 ( 
.A(n_2985),
.Y(n_3773)
);

HB1xp67_ASAP7_75t_L g3774 ( 
.A(n_3362),
.Y(n_3774)
);

NAND3xp33_ASAP7_75t_L g3775 ( 
.A(n_3372),
.B(n_362),
.C(n_361),
.Y(n_3775)
);

AOI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3082),
.A2(n_363),
.B(n_362),
.Y(n_3776)
);

BUFx6f_ASAP7_75t_L g3777 ( 
.A(n_2985),
.Y(n_3777)
);

OAI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3082),
.A2(n_37),
.B(n_38),
.Y(n_3778)
);

AOI33xp33_ASAP7_75t_L g3779 ( 
.A1(n_3007),
.A2(n_367),
.A3(n_365),
.B1(n_368),
.B2(n_366),
.B3(n_364),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3164),
.B(n_364),
.Y(n_3780)
);

A2O1A1Ixp33_ASAP7_75t_L g3781 ( 
.A1(n_3288),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_3781)
);

O2A1O1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_2995),
.A2(n_365),
.B(n_366),
.C(n_364),
.Y(n_3782)
);

BUFx4f_ASAP7_75t_L g3783 ( 
.A(n_3362),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_3083),
.A2(n_366),
.B(n_365),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3083),
.A2(n_368),
.B(n_367),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3125),
.B(n_368),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3479),
.Y(n_3787)
);

AOI21x1_ASAP7_75t_L g3788 ( 
.A1(n_3236),
.A2(n_370),
.B(n_369),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3127),
.B(n_369),
.Y(n_3789)
);

O2A1O1Ixp33_ASAP7_75t_SL g3790 ( 
.A1(n_3258),
.A2(n_370),
.B(n_371),
.C(n_369),
.Y(n_3790)
);

AND2x4_ASAP7_75t_L g3791 ( 
.A(n_3398),
.B(n_370),
.Y(n_3791)
);

AOI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3352),
.A2(n_372),
.B(n_371),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3354),
.A2(n_372),
.B(n_371),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3128),
.B(n_372),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3357),
.A2(n_374),
.B(n_373),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3310),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3313),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3483),
.Y(n_3798)
);

AOI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_3359),
.A2(n_374),
.B(n_373),
.Y(n_3799)
);

BUFx3_ASAP7_75t_L g3800 ( 
.A(n_3501),
.Y(n_3800)
);

O2A1O1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_2998),
.A2(n_374),
.B(n_375),
.C(n_373),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_L g3802 ( 
.A(n_3055),
.B(n_375),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3369),
.A2(n_376),
.B(n_375),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_2901),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3322),
.Y(n_3805)
);

AOI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3374),
.A2(n_377),
.B(n_376),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3378),
.A2(n_377),
.B(n_376),
.Y(n_3807)
);

INVx3_ASAP7_75t_L g3808 ( 
.A(n_3198),
.Y(n_3808)
);

O2A1O1Ixp33_ASAP7_75t_L g3809 ( 
.A1(n_2999),
.A2(n_378),
.B(n_379),
.C(n_377),
.Y(n_3809)
);

OAI21x1_ASAP7_75t_L g3810 ( 
.A1(n_3151),
.A2(n_3249),
.B(n_3175),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3111),
.B(n_378),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_3379),
.A2(n_380),
.B(n_379),
.Y(n_3812)
);

HB1xp67_ASAP7_75t_L g3813 ( 
.A(n_2901),
.Y(n_3813)
);

A2O1A1Ixp33_ASAP7_75t_L g3814 ( 
.A1(n_3385),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_3814)
);

O2A1O1Ixp33_ASAP7_75t_L g3815 ( 
.A1(n_3000),
.A2(n_380),
.B(n_381),
.C(n_379),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3146),
.B(n_380),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3129),
.B(n_381),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3483),
.Y(n_3818)
);

NOR2x1p5_ASAP7_75t_L g3819 ( 
.A(n_3131),
.B(n_381),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_2968),
.B(n_382),
.Y(n_3820)
);

AOI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_3052),
.A2(n_383),
.B1(n_384),
.B2(n_382),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3391),
.A2(n_383),
.B(n_382),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3140),
.B(n_383),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3245),
.B(n_384),
.Y(n_3824)
);

NAND2xp33_ASAP7_75t_L g3825 ( 
.A(n_2985),
.B(n_385),
.Y(n_3825)
);

BUFx8_ASAP7_75t_L g3826 ( 
.A(n_3113),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3484),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3400),
.A2(n_3403),
.B(n_3401),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3409),
.A2(n_386),
.B(n_385),
.Y(n_3829)
);

INVx3_ASAP7_75t_L g3830 ( 
.A(n_3115),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3497),
.B(n_385),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_SL g3832 ( 
.A(n_3189),
.B(n_387),
.Y(n_3832)
);

BUFx12f_ASAP7_75t_L g3833 ( 
.A(n_2928),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3142),
.B(n_388),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_3376),
.B(n_389),
.Y(n_3835)
);

OAI21x1_ASAP7_75t_L g3836 ( 
.A1(n_3175),
.A2(n_390),
.B(n_389),
.Y(n_3836)
);

AOI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3056),
.A2(n_390),
.B1(n_391),
.B2(n_389),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3412),
.A2(n_393),
.B(n_392),
.Y(n_3838)
);

AOI21xp5_ASAP7_75t_L g3839 ( 
.A1(n_3414),
.A2(n_393),
.B(n_392),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3421),
.A2(n_393),
.B(n_392),
.Y(n_3840)
);

AOI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_3425),
.A2(n_395),
.B(n_394),
.Y(n_3841)
);

AOI22xp5_ASAP7_75t_L g3842 ( 
.A1(n_3058),
.A2(n_395),
.B1(n_396),
.B2(n_394),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3484),
.Y(n_3843)
);

BUFx12f_ASAP7_75t_L g3844 ( 
.A(n_3097),
.Y(n_3844)
);

OAI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3433),
.A2(n_396),
.B1(n_397),
.B2(n_395),
.Y(n_3845)
);

NOR2xp33_ASAP7_75t_L g3846 ( 
.A(n_3407),
.B(n_396),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3189),
.B(n_397),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3485),
.Y(n_3848)
);

BUFx3_ASAP7_75t_L g3849 ( 
.A(n_3138),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3147),
.B(n_398),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3168),
.B(n_3126),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3149),
.B(n_399),
.Y(n_3852)
);

AOI21xp5_ASAP7_75t_L g3853 ( 
.A1(n_3441),
.A2(n_400),
.B(n_399),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3444),
.A2(n_3536),
.B(n_3534),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3485),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3153),
.B(n_400),
.Y(n_3856)
);

O2A1O1Ixp5_ASAP7_75t_L g3857 ( 
.A1(n_3405),
.A2(n_402),
.B(n_403),
.C(n_401),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3060),
.A2(n_402),
.B1(n_403),
.B2(n_401),
.Y(n_3858)
);

INVx2_ASAP7_75t_SL g3859 ( 
.A(n_3097),
.Y(n_3859)
);

NOR2xp33_ASAP7_75t_L g3860 ( 
.A(n_3513),
.B(n_3116),
.Y(n_3860)
);

O2A1O1Ixp33_ASAP7_75t_L g3861 ( 
.A1(n_3416),
.A2(n_405),
.B(n_406),
.C(n_404),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3253),
.B(n_404),
.Y(n_3862)
);

NOR2xp33_ASAP7_75t_L g3863 ( 
.A(n_2916),
.B(n_405),
.Y(n_3863)
);

CKINVDCx10_ASAP7_75t_R g3864 ( 
.A(n_3335),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3139),
.B(n_405),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3491),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3449),
.A2(n_407),
.B(n_406),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3328),
.B(n_2952),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3214),
.B(n_3221),
.Y(n_3869)
);

NOR2x2_ASAP7_75t_L g3870 ( 
.A(n_3335),
.B(n_406),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_2978),
.B(n_408),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3491),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3201),
.B(n_408),
.Y(n_3873)
);

O2A1O1Ixp33_ASAP7_75t_L g3874 ( 
.A1(n_3418),
.A2(n_410),
.B(n_411),
.C(n_409),
.Y(n_3874)
);

BUFx6f_ASAP7_75t_L g3875 ( 
.A(n_3189),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3452),
.A2(n_410),
.B(n_409),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3455),
.A2(n_412),
.B(n_411),
.Y(n_3877)
);

AOI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_2976),
.A2(n_413),
.B1(n_414),
.B2(n_412),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3456),
.A2(n_414),
.B(n_413),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3194),
.B(n_413),
.Y(n_3880)
);

AOI22xp5_ASAP7_75t_L g3881 ( 
.A1(n_2941),
.A2(n_415),
.B1(n_416),
.B2(n_414),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3458),
.A2(n_416),
.B(n_415),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_2981),
.B(n_3326),
.Y(n_3883)
);

OAI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3057),
.A2(n_39),
.B(n_40),
.Y(n_3884)
);

INVx2_ASAP7_75t_SL g3885 ( 
.A(n_3402),
.Y(n_3885)
);

INVx11_ASAP7_75t_L g3886 ( 
.A(n_3402),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3462),
.A2(n_3539),
.B(n_3537),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3326),
.B(n_415),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3465),
.A2(n_418),
.B(n_417),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3186),
.B(n_418),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3527),
.A2(n_419),
.B(n_418),
.Y(n_3891)
);

BUFx12f_ASAP7_75t_L g3892 ( 
.A(n_3047),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3338),
.B(n_419),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3123),
.B(n_421),
.Y(n_3894)
);

INVx3_ASAP7_75t_L g3895 ( 
.A(n_3240),
.Y(n_3895)
);

OAI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_2965),
.A2(n_41),
.B(n_42),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3339),
.B(n_421),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3182),
.B(n_422),
.Y(n_3898)
);

CKINVDCx20_ASAP7_75t_R g3899 ( 
.A(n_3021),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3351),
.B(n_422),
.Y(n_3900)
);

A2O1A1Ixp33_ASAP7_75t_L g3901 ( 
.A1(n_3543),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3492),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3156),
.B(n_423),
.Y(n_3903)
);

OAI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3335),
.A2(n_424),
.B1(n_425),
.B2(n_423),
.Y(n_3904)
);

NAND2x1_ASAP7_75t_L g3905 ( 
.A(n_3240),
.B(n_423),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3377),
.B(n_3389),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3091),
.A2(n_425),
.B(n_424),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3393),
.B(n_3413),
.Y(n_3908)
);

OAI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_2969),
.A2(n_42),
.B(n_43),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3492),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3415),
.B(n_424),
.Y(n_3911)
);

NOR2xp33_ASAP7_75t_L g3912 ( 
.A(n_3174),
.B(n_426),
.Y(n_3912)
);

AOI22xp5_ASAP7_75t_L g3913 ( 
.A1(n_2997),
.A2(n_427),
.B1(n_428),
.B2(n_426),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3426),
.B(n_427),
.Y(n_3914)
);

BUFx3_ASAP7_75t_L g3915 ( 
.A(n_2921),
.Y(n_3915)
);

A2O1A1Ixp33_ASAP7_75t_L g3916 ( 
.A1(n_3355),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3495),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3495),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3438),
.B(n_427),
.Y(n_3919)
);

HB1xp67_ASAP7_75t_L g3920 ( 
.A(n_3155),
.Y(n_3920)
);

OAI21xp33_ASAP7_75t_L g3921 ( 
.A1(n_3003),
.A2(n_44),
.B(n_45),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3473),
.B(n_428),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3091),
.A2(n_429),
.B(n_428),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3476),
.B(n_429),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3499),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_SL g3926 ( 
.A(n_3240),
.B(n_429),
.Y(n_3926)
);

OAI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_2970),
.A2(n_44),
.B(n_45),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3493),
.B(n_430),
.Y(n_3928)
);

CKINVDCx10_ASAP7_75t_R g3929 ( 
.A(n_3155),
.Y(n_3929)
);

AOI33xp33_ASAP7_75t_L g3930 ( 
.A1(n_3048),
.A2(n_433),
.A3(n_431),
.B1(n_434),
.B2(n_432),
.B3(n_430),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_2971),
.A2(n_432),
.B(n_431),
.Y(n_3931)
);

AOI21x1_ASAP7_75t_L g3932 ( 
.A1(n_2894),
.A2(n_3159),
.B(n_3158),
.Y(n_3932)
);

O2A1O1Ixp33_ASAP7_75t_L g3933 ( 
.A1(n_3437),
.A2(n_432),
.B(n_433),
.C(n_431),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3499),
.Y(n_3934)
);

A2O1A1Ixp33_ASAP7_75t_L g3935 ( 
.A1(n_3148),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3502),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3505),
.B(n_434),
.Y(n_3937)
);

HB1xp67_ASAP7_75t_L g3938 ( 
.A(n_3155),
.Y(n_3938)
);

BUFx6f_ASAP7_75t_L g3939 ( 
.A(n_3323),
.Y(n_3939)
);

OAI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_2973),
.A2(n_45),
.B(n_46),
.Y(n_3940)
);

BUFx4f_ASAP7_75t_L g3941 ( 
.A(n_3184),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_2979),
.A2(n_435),
.B(n_434),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_2988),
.A2(n_436),
.B(n_435),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3507),
.B(n_436),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3173),
.A2(n_437),
.B(n_436),
.Y(n_3945)
);

OAI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3439),
.A2(n_46),
.B(n_47),
.Y(n_3946)
);

AOI21xp5_ASAP7_75t_L g3947 ( 
.A1(n_3173),
.A2(n_438),
.B(n_437),
.Y(n_3947)
);

AOI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3446),
.A2(n_438),
.B(n_437),
.Y(n_3948)
);

OAI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3454),
.A2(n_46),
.B(n_47),
.Y(n_3949)
);

OAI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3457),
.A2(n_48),
.B(n_49),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3528),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3529),
.B(n_438),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3530),
.B(n_439),
.Y(n_3953)
);

OAI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3494),
.A2(n_48),
.B(n_49),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3535),
.B(n_439),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3496),
.A2(n_440),
.B(n_439),
.Y(n_3956)
);

AOI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3498),
.A2(n_441),
.B(n_440),
.Y(n_3957)
);

HB1xp67_ASAP7_75t_L g3958 ( 
.A(n_2886),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3538),
.B(n_440),
.Y(n_3959)
);

AOI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_3533),
.A2(n_3541),
.B(n_3300),
.Y(n_3960)
);

INVx3_ASAP7_75t_L g3961 ( 
.A(n_3323),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3323),
.B(n_441),
.Y(n_3962)
);

AOI21x1_ASAP7_75t_L g3963 ( 
.A1(n_2894),
.A2(n_442),
.B(n_441),
.Y(n_3963)
);

AOI33xp33_ASAP7_75t_L g3964 ( 
.A1(n_3124),
.A2(n_445),
.A3(n_443),
.B1(n_446),
.B2(n_444),
.B3(n_442),
.Y(n_3964)
);

BUFx3_ASAP7_75t_L g3965 ( 
.A(n_2921),
.Y(n_3965)
);

A2O1A1Ixp33_ASAP7_75t_L g3966 ( 
.A1(n_3502),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_3966)
);

AOI21xp5_ASAP7_75t_L g3967 ( 
.A1(n_3059),
.A2(n_444),
.B(n_443),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3065),
.A2(n_446),
.B(n_445),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3078),
.A2(n_447),
.B(n_446),
.Y(n_3969)
);

AND2x2_ASAP7_75t_SL g3970 ( 
.A(n_3297),
.B(n_447),
.Y(n_3970)
);

NOR3xp33_ASAP7_75t_L g3971 ( 
.A(n_3063),
.B(n_448),
.C(n_447),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3508),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3265),
.B(n_448),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_SL g3974 ( 
.A(n_3363),
.B(n_448),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3010),
.B(n_449),
.Y(n_3975)
);

OAI21xp33_ASAP7_75t_L g3976 ( 
.A1(n_3331),
.A2(n_49),
.B(n_50),
.Y(n_3976)
);

INVx3_ASAP7_75t_L g3977 ( 
.A(n_3363),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3508),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_2986),
.B(n_449),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3363),
.B(n_450),
.Y(n_3980)
);

AND2x4_ASAP7_75t_L g3981 ( 
.A(n_3340),
.B(n_450),
.Y(n_3981)
);

O2A1O1Ixp33_ASAP7_75t_L g3982 ( 
.A1(n_3040),
.A2(n_451),
.B(n_452),
.C(n_450),
.Y(n_3982)
);

OAI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3070),
.A2(n_50),
.B(n_51),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_3445),
.B(n_451),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_2994),
.B(n_452),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_SL g3986 ( 
.A(n_3445),
.B(n_452),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3512),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3090),
.A2(n_454),
.B(n_453),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3512),
.Y(n_3989)
);

OAI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_3098),
.A2(n_51),
.B(n_52),
.Y(n_3990)
);

INVx2_ASAP7_75t_L g3991 ( 
.A(n_2992),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3185),
.B(n_453),
.Y(n_3992)
);

AOI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_3297),
.A2(n_454),
.B(n_453),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3445),
.B(n_454),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3190),
.B(n_455),
.Y(n_3995)
);

AO21x1_ASAP7_75t_L g3996 ( 
.A1(n_3521),
.A2(n_3298),
.B(n_3519),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3008),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_2895),
.B(n_455),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3279),
.A2(n_457),
.B(n_456),
.Y(n_3999)
);

BUFx12f_ASAP7_75t_L g4000 ( 
.A(n_3366),
.Y(n_4000)
);

BUFx4f_ASAP7_75t_L g4001 ( 
.A(n_3270),
.Y(n_4001)
);

OAI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3459),
.A2(n_3477),
.B1(n_3488),
.B2(n_3463),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3489),
.A2(n_457),
.B1(n_458),
.B2(n_456),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3176),
.A2(n_458),
.B(n_457),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3176),
.A2(n_460),
.B(n_459),
.Y(n_4005)
);

BUFx6f_ASAP7_75t_L g4006 ( 
.A(n_3532),
.Y(n_4006)
);

OAI321xp33_ASAP7_75t_L g4007 ( 
.A1(n_3387),
.A2(n_53),
.A3(n_55),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_4007)
);

CKINVDCx20_ASAP7_75t_R g4008 ( 
.A(n_2923),
.Y(n_4008)
);

NOR2x1_ASAP7_75t_R g4009 ( 
.A(n_3163),
.B(n_459),
.Y(n_4009)
);

BUFx12f_ASAP7_75t_L g4010 ( 
.A(n_3223),
.Y(n_4010)
);

OAI22x1_ASAP7_75t_L g4011 ( 
.A1(n_3436),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_SL g4012 ( 
.A(n_3532),
.B(n_461),
.Y(n_4012)
);

INVxp67_ASAP7_75t_L g4013 ( 
.A(n_2898),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3177),
.A2(n_462),
.B(n_461),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3177),
.A2(n_463),
.B(n_462),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3519),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3522),
.Y(n_4017)
);

INVx4_ASAP7_75t_L g4018 ( 
.A(n_3340),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3522),
.Y(n_4019)
);

OAI21xp5_ASAP7_75t_L g4020 ( 
.A1(n_3050),
.A2(n_51),
.B(n_52),
.Y(n_4020)
);

INVxp67_ASAP7_75t_L g4021 ( 
.A(n_3210),
.Y(n_4021)
);

NOR3xp33_ASAP7_75t_L g4022 ( 
.A(n_2987),
.B(n_464),
.C(n_463),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3178),
.A2(n_464),
.B(n_463),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3178),
.A2(n_465),
.B(n_464),
.Y(n_4024)
);

AOI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_2885),
.A2(n_466),
.B(n_465),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3532),
.B(n_465),
.Y(n_4026)
);

INVx3_ASAP7_75t_L g4027 ( 
.A(n_3381),
.Y(n_4027)
);

CKINVDCx10_ASAP7_75t_R g4028 ( 
.A(n_2925),
.Y(n_4028)
);

HB1xp67_ASAP7_75t_L g4029 ( 
.A(n_2918),
.Y(n_4029)
);

INVx3_ASAP7_75t_L g4030 ( 
.A(n_3381),
.Y(n_4030)
);

BUFx4f_ASAP7_75t_L g4031 ( 
.A(n_3209),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3199),
.B(n_466),
.Y(n_4032)
);

AOI21xp5_ASAP7_75t_L g4033 ( 
.A1(n_3320),
.A2(n_467),
.B(n_466),
.Y(n_4033)
);

INVx4_ASAP7_75t_L g4034 ( 
.A(n_3518),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_3145),
.A2(n_468),
.B(n_467),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3213),
.B(n_468),
.Y(n_4036)
);

AND2x4_ASAP7_75t_L g4037 ( 
.A(n_3518),
.B(n_468),
.Y(n_4037)
);

NAND2x1p5_ASAP7_75t_L g4038 ( 
.A(n_3208),
.B(n_2947),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3217),
.B(n_469),
.Y(n_4039)
);

INVx3_ASAP7_75t_L g4040 ( 
.A(n_3280),
.Y(n_4040)
);

AO21x1_ASAP7_75t_L g4041 ( 
.A1(n_3298),
.A2(n_470),
.B(n_469),
.Y(n_4041)
);

AOI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3525),
.A2(n_471),
.B(n_470),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3525),
.A2(n_471),
.B(n_470),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3461),
.B(n_3470),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3154),
.B(n_471),
.Y(n_4045)
);

INVxp67_ASAP7_75t_L g4046 ( 
.A(n_3103),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_SL g4047 ( 
.A(n_2996),
.B(n_472),
.Y(n_4047)
);

AOI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_2962),
.A2(n_3075),
.B(n_3067),
.Y(n_4048)
);

OAI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3012),
.A2(n_473),
.B1(n_474),
.B2(n_472),
.Y(n_4049)
);

O2A1O1Ixp33_ASAP7_75t_L g4050 ( 
.A1(n_3042),
.A2(n_474),
.B(n_475),
.C(n_473),
.Y(n_4050)
);

OAI21xp33_ASAP7_75t_L g4051 ( 
.A1(n_3341),
.A2(n_3045),
.B(n_3303),
.Y(n_4051)
);

AOI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3076),
.A2(n_474),
.B(n_473),
.Y(n_4052)
);

INVx2_ASAP7_75t_L g4053 ( 
.A(n_3077),
.Y(n_4053)
);

AOI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3080),
.A2(n_3252),
.B(n_3255),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3112),
.B(n_475),
.Y(n_4055)
);

OAI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_3134),
.A2(n_53),
.B(n_54),
.Y(n_4056)
);

OAI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3135),
.A2(n_53),
.B(n_54),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_2961),
.B(n_476),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_2975),
.B(n_476),
.Y(n_4059)
);

AOI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3267),
.A2(n_477),
.B(n_476),
.Y(n_4060)
);

A2O1A1Ixp33_ASAP7_75t_L g4061 ( 
.A1(n_3283),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_2936),
.B(n_478),
.Y(n_4062)
);

O2A1O1Ixp33_ASAP7_75t_L g4063 ( 
.A1(n_3094),
.A2(n_479),
.B(n_480),
.C(n_478),
.Y(n_4063)
);

AOI21xp33_ASAP7_75t_L g4064 ( 
.A1(n_3332),
.A2(n_480),
.B(n_479),
.Y(n_4064)
);

AOI22xp5_ASAP7_75t_L g4065 ( 
.A1(n_3017),
.A2(n_3022),
.B1(n_2892),
.B2(n_3276),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3234),
.Y(n_4066)
);

AOI21xp5_ASAP7_75t_L g4067 ( 
.A1(n_3358),
.A2(n_481),
.B(n_480),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_2940),
.B(n_481),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3018),
.B(n_482),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3019),
.B(n_483),
.Y(n_4070)
);

AOI21xp5_ASAP7_75t_L g4071 ( 
.A1(n_3218),
.A2(n_486),
.B(n_484),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3248),
.Y(n_4072)
);

OAI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_3225),
.A2(n_55),
.B(n_56),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3222),
.A2(n_486),
.B(n_484),
.Y(n_4074)
);

AOI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_3226),
.A2(n_487),
.B(n_486),
.Y(n_4075)
);

CKINVDCx5p33_ASAP7_75t_R g4076 ( 
.A(n_3086),
.Y(n_4076)
);

OAI321xp33_ASAP7_75t_L g4077 ( 
.A1(n_3167),
.A2(n_57),
.A3(n_59),
.B1(n_55),
.B2(n_56),
.C(n_58),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_3247),
.B(n_487),
.Y(n_4078)
);

NOR2xp33_ASAP7_75t_L g4079 ( 
.A(n_3061),
.B(n_488),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_3227),
.A2(n_489),
.B(n_488),
.Y(n_4080)
);

BUFx2_ASAP7_75t_L g4081 ( 
.A(n_2938),
.Y(n_4081)
);

BUFx3_ASAP7_75t_L g4082 ( 
.A(n_2993),
.Y(n_4082)
);

BUFx3_ASAP7_75t_L g4083 ( 
.A(n_3318),
.Y(n_4083)
);

INVx1_ASAP7_75t_SL g4084 ( 
.A(n_3336),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3110),
.B(n_488),
.Y(n_4085)
);

NOR2xp33_ASAP7_75t_L g4086 ( 
.A(n_2980),
.B(n_489),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3183),
.B(n_490),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3262),
.Y(n_4088)
);

AOI21x1_ASAP7_75t_L g4089 ( 
.A1(n_3275),
.A2(n_491),
.B(n_490),
.Y(n_4089)
);

NAND2x1p5_ASAP7_75t_L g4090 ( 
.A(n_3360),
.B(n_491),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3250),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_3229),
.A2(n_493),
.B(n_492),
.Y(n_4092)
);

AOI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_3233),
.A2(n_494),
.B(n_492),
.Y(n_4093)
);

AOI21xp5_ASAP7_75t_L g4094 ( 
.A1(n_3235),
.A2(n_495),
.B(n_494),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3188),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3349),
.B(n_494),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3041),
.B(n_495),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_2948),
.B(n_496),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_SL g4099 ( 
.A(n_2929),
.B(n_496),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_SL g4100 ( 
.A(n_3152),
.B(n_3373),
.Y(n_4100)
);

INVxp67_ASAP7_75t_L g4101 ( 
.A(n_2933),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_2951),
.B(n_497),
.Y(n_4102)
);

CKINVDCx20_ASAP7_75t_R g4103 ( 
.A(n_3397),
.Y(n_4103)
);

BUFx6f_ASAP7_75t_L g4104 ( 
.A(n_3249),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3272),
.Y(n_4105)
);

INVx3_ASAP7_75t_L g4106 ( 
.A(n_3239),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_3246),
.A2(n_498),
.B(n_497),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3281),
.A2(n_498),
.B(n_497),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3542),
.B(n_499),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3013),
.B(n_499),
.Y(n_4110)
);

OAI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3030),
.A2(n_56),
.B(n_57),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3062),
.B(n_500),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3132),
.Y(n_4113)
);

O2A1O1Ixp33_ASAP7_75t_L g4114 ( 
.A1(n_3096),
.A2(n_501),
.B(n_502),
.C(n_500),
.Y(n_4114)
);

BUFx2_ASAP7_75t_L g4115 ( 
.A(n_3480),
.Y(n_4115)
);

BUFx3_ASAP7_75t_L g4116 ( 
.A(n_3510),
.Y(n_4116)
);

A2O1A1Ixp33_ASAP7_75t_L g4117 ( 
.A1(n_3551),
.A2(n_3314),
.B(n_3220),
.C(n_3161),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3558),
.B(n_3315),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_3669),
.B(n_3411),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3783),
.B(n_3239),
.Y(n_4120)
);

INVx1_ASAP7_75t_SL g4121 ( 
.A(n_4103),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_4105),
.B(n_3557),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3576),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3783),
.B(n_3232),
.Y(n_4124)
);

BUFx2_ASAP7_75t_L g4125 ( 
.A(n_3719),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3547),
.Y(n_4126)
);

AND2x2_ASAP7_75t_SL g4127 ( 
.A(n_3970),
.B(n_3054),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_3973),
.B(n_2983),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_4046),
.B(n_3105),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3828),
.A2(n_3334),
.B(n_3277),
.Y(n_4130)
);

NAND3xp33_ASAP7_75t_SL g4131 ( 
.A(n_3651),
.B(n_3212),
.C(n_3193),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_L g4132 ( 
.A(n_4065),
.B(n_3005),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3585),
.B(n_3317),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3550),
.B(n_3607),
.Y(n_4134)
);

INVx5_ASAP7_75t_L g4135 ( 
.A(n_3833),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3588),
.B(n_3321),
.Y(n_4136)
);

INVx2_ASAP7_75t_SL g4137 ( 
.A(n_4031),
.Y(n_4137)
);

OAI22xp5_ASAP7_75t_L g4138 ( 
.A1(n_3723),
.A2(n_2972),
.B1(n_2955),
.B2(n_3130),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_3688),
.B(n_3095),
.Y(n_4139)
);

O2A1O1Ixp33_ASAP7_75t_L g4140 ( 
.A1(n_4051),
.A2(n_3365),
.B(n_3367),
.C(n_3361),
.Y(n_4140)
);

INVx2_ASAP7_75t_L g4141 ( 
.A(n_3603),
.Y(n_4141)
);

A2O1A1Ixp33_ASAP7_75t_L g4142 ( 
.A1(n_3555),
.A2(n_3294),
.B(n_3211),
.C(n_3230),
.Y(n_4142)
);

A2O1A1Ixp33_ASAP7_75t_L g4143 ( 
.A1(n_3713),
.A2(n_2983),
.B(n_3531),
.C(n_3517),
.Y(n_4143)
);

INVx6_ASAP7_75t_L g4144 ( 
.A(n_3618),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_3608),
.Y(n_4145)
);

A2O1A1Ixp33_ASAP7_75t_L g4146 ( 
.A1(n_3975),
.A2(n_3371),
.B(n_3392),
.C(n_3390),
.Y(n_4146)
);

OR2x2_ASAP7_75t_L g4147 ( 
.A(n_4021),
.B(n_3448),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3622),
.Y(n_4148)
);

OAI21xp33_ASAP7_75t_L g4149 ( 
.A1(n_3863),
.A2(n_3324),
.B(n_3257),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3623),
.Y(n_4150)
);

OAI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_3641),
.A2(n_3356),
.B1(n_3429),
.B2(n_3419),
.Y(n_4151)
);

AOI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_3854),
.A2(n_3278),
.B(n_3203),
.Y(n_4152)
);

BUFx6f_ASAP7_75t_L g4153 ( 
.A(n_3618),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3643),
.Y(n_4154)
);

OAI21xp33_ASAP7_75t_L g4155 ( 
.A1(n_3779),
.A2(n_3410),
.B(n_3404),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3648),
.Y(n_4156)
);

AND2x4_ASAP7_75t_L g4157 ( 
.A(n_3688),
.B(n_3268),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3831),
.B(n_3104),
.Y(n_4158)
);

AOI21xp5_ASAP7_75t_L g4159 ( 
.A1(n_3887),
.A2(n_3224),
.B(n_3197),
.Y(n_4159)
);

OAI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_3641),
.A2(n_3066),
.B1(n_3181),
.B2(n_3207),
.Y(n_4160)
);

AO32x2_ASAP7_75t_L g4161 ( 
.A1(n_3904),
.A2(n_3704),
.A3(n_4002),
.B1(n_3595),
.B2(n_3571),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3652),
.Y(n_4162)
);

BUFx6f_ASAP7_75t_L g4163 ( 
.A(n_3618),
.Y(n_4163)
);

AOI21xp5_ASAP7_75t_L g4164 ( 
.A1(n_3699),
.A2(n_3237),
.B(n_3228),
.Y(n_4164)
);

A2O1A1Ixp33_ASAP7_75t_SL g4165 ( 
.A1(n_3597),
.A2(n_3386),
.B(n_3431),
.C(n_3430),
.Y(n_4165)
);

O2A1O1Ixp33_ASAP7_75t_L g4166 ( 
.A1(n_3851),
.A2(n_3434),
.B(n_3453),
.C(n_3432),
.Y(n_4166)
);

HB1xp67_ASAP7_75t_L g4167 ( 
.A(n_3627),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_3611),
.Y(n_4168)
);

INVx3_ASAP7_75t_L g4169 ( 
.A(n_4031),
.Y(n_4169)
);

AOI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_3758),
.A2(n_3074),
.B1(n_3087),
.B2(n_3064),
.Y(n_4170)
);

CKINVDCx5p33_ASAP7_75t_R g4171 ( 
.A(n_3844),
.Y(n_4171)
);

A2O1A1Ixp33_ASAP7_75t_L g4172 ( 
.A1(n_3921),
.A2(n_3471),
.B(n_3486),
.C(n_3464),
.Y(n_4172)
);

INVx3_ASAP7_75t_SL g4173 ( 
.A(n_3600),
.Y(n_4173)
);

OAI22xp5_ASAP7_75t_SL g4174 ( 
.A1(n_4010),
.A2(n_3192),
.B1(n_3490),
.B2(n_3487),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_3548),
.B(n_2913),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_3753),
.A2(n_3242),
.B(n_3251),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_3673),
.A2(n_3868),
.B1(n_3971),
.B2(n_4058),
.Y(n_4177)
);

AOI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_3717),
.A2(n_3200),
.B(n_3150),
.Y(n_4178)
);

OAI21xp33_ASAP7_75t_L g4179 ( 
.A1(n_3869),
.A2(n_3930),
.B(n_3703),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4091),
.B(n_3089),
.Y(n_4180)
);

BUFx6f_ASAP7_75t_L g4181 ( 
.A(n_3546),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3677),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_3587),
.A2(n_3202),
.B(n_3215),
.Y(n_4183)
);

INVx1_ASAP7_75t_SL g4184 ( 
.A(n_3710),
.Y(n_4184)
);

AND2x2_ASAP7_75t_L g4185 ( 
.A(n_3898),
.B(n_3104),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_SL g4186 ( 
.A(n_3550),
.B(n_3516),
.Y(n_4186)
);

NAND2x2_ASAP7_75t_L g4187 ( 
.A(n_3819),
.B(n_3028),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3716),
.B(n_3006),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_3549),
.B(n_2914),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3613),
.Y(n_4190)
);

OAI22xp5_ASAP7_75t_L g4191 ( 
.A1(n_3883),
.A2(n_3133),
.B1(n_3287),
.B2(n_3293),
.Y(n_4191)
);

O2A1O1Ixp33_ASAP7_75t_SL g4192 ( 
.A1(n_3610),
.A2(n_3141),
.B(n_3216),
.C(n_3299),
.Y(n_4192)
);

BUFx6f_ASAP7_75t_L g4193 ( 
.A(n_3546),
.Y(n_4193)
);

AOI21x1_ASAP7_75t_L g4194 ( 
.A1(n_3996),
.A2(n_3544),
.B(n_3289),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_3960),
.A2(n_3296),
.B(n_3295),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_3615),
.A2(n_3291),
.B(n_3290),
.Y(n_4196)
);

NOR3xp33_ASAP7_75t_L g4197 ( 
.A(n_4009),
.B(n_3553),
.C(n_3759),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3687),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_3732),
.B(n_3205),
.Y(n_4199)
);

AND2x2_ASAP7_75t_SL g4200 ( 
.A(n_3586),
.B(n_3122),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4072),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4066),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3683),
.A2(n_3273),
.B(n_3269),
.Y(n_4203)
);

O2A1O1Ixp33_ASAP7_75t_L g4204 ( 
.A1(n_3617),
.A2(n_2915),
.B(n_3068),
.C(n_3016),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3756),
.B(n_3206),
.Y(n_4205)
);

BUFx2_ASAP7_75t_L g4206 ( 
.A(n_3719),
.Y(n_4206)
);

A2O1A1Ixp33_ASAP7_75t_SL g4207 ( 
.A1(n_3983),
.A2(n_3120),
.B(n_3274),
.C(n_3292),
.Y(n_4207)
);

OAI21xp33_ASAP7_75t_L g4208 ( 
.A1(n_3692),
.A2(n_3241),
.B(n_3219),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_3658),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3765),
.B(n_3243),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3672),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_3678),
.Y(n_4212)
);

BUFx10_ASAP7_75t_L g4213 ( 
.A(n_3565),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3766),
.B(n_3244),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3787),
.B(n_3231),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_3894),
.B(n_3117),
.Y(n_4216)
);

NAND2xp33_ASAP7_75t_R g4217 ( 
.A(n_4076),
.B(n_500),
.Y(n_4217)
);

NOR2xp33_ASAP7_75t_L g4218 ( 
.A(n_3566),
.B(n_3014),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_3680),
.Y(n_4219)
);

INVx2_ASAP7_75t_L g4220 ( 
.A(n_4053),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_L g4221 ( 
.A(n_3653),
.B(n_2893),
.Y(n_4221)
);

CKINVDCx16_ASAP7_75t_R g4222 ( 
.A(n_3675),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_3698),
.A2(n_3260),
.B(n_3191),
.Y(n_4223)
);

O2A1O1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_3616),
.A2(n_3102),
.B(n_2966),
.C(n_2989),
.Y(n_4224)
);

AOI21xp5_ASAP7_75t_L g4225 ( 
.A1(n_3798),
.A2(n_3160),
.B(n_3136),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_3593),
.Y(n_4226)
);

OAI21x1_ASAP7_75t_L g4227 ( 
.A1(n_3810),
.A2(n_3114),
.B(n_3170),
.Y(n_4227)
);

OAI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_3605),
.A2(n_3172),
.B1(n_2949),
.B2(n_3254),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3818),
.B(n_3827),
.Y(n_4229)
);

NOR2xp33_ASAP7_75t_L g4230 ( 
.A(n_3755),
.B(n_2924),
.Y(n_4230)
);

A2O1A1Ixp33_ASAP7_75t_L g4231 ( 
.A1(n_3748),
.A2(n_3264),
.B(n_3263),
.C(n_3266),
.Y(n_4231)
);

A2O1A1Ixp33_ASAP7_75t_L g4232 ( 
.A1(n_3764),
.A2(n_3282),
.B(n_2932),
.C(n_2926),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_3742),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_3843),
.B(n_501),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_3594),
.Y(n_4235)
);

NOR2xp33_ASAP7_75t_L g4236 ( 
.A(n_3864),
.B(n_501),
.Y(n_4236)
);

CKINVDCx16_ASAP7_75t_R g4237 ( 
.A(n_3767),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_3848),
.B(n_502),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3855),
.B(n_502),
.Y(n_4239)
);

OR2x2_ASAP7_75t_L g4240 ( 
.A(n_3679),
.B(n_503),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_3638),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.Y(n_4241)
);

OAI22xp5_ASAP7_75t_L g4242 ( 
.A1(n_3866),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_3872),
.A2(n_506),
.B(n_505),
.Y(n_4243)
);

AOI21xp5_ASAP7_75t_L g4244 ( 
.A1(n_3902),
.A2(n_507),
.B(n_506),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_SL g4245 ( 
.A(n_3550),
.B(n_506),
.Y(n_4245)
);

OR2x2_ASAP7_75t_L g4246 ( 
.A(n_3706),
.B(n_3709),
.Y(n_4246)
);

BUFx3_ASAP7_75t_L g4247 ( 
.A(n_3826),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_R g4248 ( 
.A(n_3929),
.B(n_507),
.Y(n_4248)
);

O2A1O1Ixp33_ASAP7_75t_SL g4249 ( 
.A1(n_3662),
.A2(n_1117),
.B(n_1118),
.C(n_1116),
.Y(n_4249)
);

O2A1O1Ixp33_ASAP7_75t_L g4250 ( 
.A1(n_3736),
.A2(n_508),
.B(n_509),
.C(n_507),
.Y(n_4250)
);

BUFx6f_ASAP7_75t_L g4251 ( 
.A(n_3546),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_3550),
.B(n_508),
.Y(n_4252)
);

OAI21xp33_ASAP7_75t_L g4253 ( 
.A1(n_3561),
.A2(n_56),
.B(n_58),
.Y(n_4253)
);

OAI21xp33_ASAP7_75t_L g4254 ( 
.A1(n_3964),
.A2(n_58),
.B(n_59),
.Y(n_4254)
);

O2A1O1Ixp33_ASAP7_75t_L g4255 ( 
.A1(n_3743),
.A2(n_509),
.B(n_510),
.C(n_508),
.Y(n_4255)
);

NOR3xp33_ASAP7_75t_L g4256 ( 
.A(n_3820),
.B(n_511),
.C(n_509),
.Y(n_4256)
);

INVx3_ASAP7_75t_SL g4257 ( 
.A(n_3870),
.Y(n_4257)
);

CKINVDCx6p67_ASAP7_75t_R g4258 ( 
.A(n_4028),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_3910),
.B(n_3917),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_3918),
.A2(n_512),
.B(n_511),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_3824),
.B(n_1108),
.Y(n_4261)
);

INVxp67_ASAP7_75t_L g4262 ( 
.A(n_4081),
.Y(n_4262)
);

HB1xp67_ASAP7_75t_L g4263 ( 
.A(n_3573),
.Y(n_4263)
);

AOI221xp5_ASAP7_75t_L g4264 ( 
.A1(n_4110),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.C(n_512),
.Y(n_4264)
);

AND2x2_ASAP7_75t_SL g4265 ( 
.A(n_3730),
.B(n_512),
.Y(n_4265)
);

O2A1O1Ixp33_ASAP7_75t_L g4266 ( 
.A1(n_4087),
.A2(n_514),
.B(n_515),
.C(n_513),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3599),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_3635),
.Y(n_4268)
);

INVx4_ASAP7_75t_L g4269 ( 
.A(n_3886),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_R g4270 ( 
.A(n_3826),
.B(n_515),
.Y(n_4270)
);

OAI22xp5_ASAP7_75t_L g4271 ( 
.A1(n_3925),
.A2(n_517),
.B1(n_518),
.B2(n_516),
.Y(n_4271)
);

AND2x6_ASAP7_75t_L g4272 ( 
.A(n_3655),
.B(n_517),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_3768),
.Y(n_4273)
);

NOR2xp33_ASAP7_75t_L g4274 ( 
.A(n_4101),
.B(n_517),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3906),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_3934),
.A2(n_3972),
.B(n_3936),
.Y(n_4276)
);

BUFx6f_ASAP7_75t_L g4277 ( 
.A(n_3656),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_3978),
.A2(n_520),
.B(n_519),
.Y(n_4278)
);

NOR2xp33_ASAP7_75t_L g4279 ( 
.A(n_3804),
.B(n_519),
.Y(n_4279)
);

A2O1A1Ixp33_ASAP7_75t_L g4280 ( 
.A1(n_3634),
.A2(n_520),
.B(n_521),
.C(n_519),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_3708),
.B(n_1116),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_3796),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_3797),
.Y(n_4283)
);

NOR2xp33_ASAP7_75t_R g4284 ( 
.A(n_3899),
.B(n_520),
.Y(n_4284)
);

INVx2_ASAP7_75t_SL g4285 ( 
.A(n_3941),
.Y(n_4285)
);

BUFx4f_ASAP7_75t_L g4286 ( 
.A(n_4000),
.Y(n_4286)
);

OAI21xp33_ASAP7_75t_SL g4287 ( 
.A1(n_3729),
.A2(n_522),
.B(n_521),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_3987),
.A2(n_522),
.B(n_521),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_3559),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_3730),
.B(n_522),
.Y(n_4290)
);

NOR2xp33_ASAP7_75t_L g4291 ( 
.A(n_3813),
.B(n_523),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_3805),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_3908),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3951),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_3903),
.B(n_1120),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3989),
.B(n_523),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_SL g4297 ( 
.A(n_3656),
.B(n_523),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_3609),
.B(n_1121),
.Y(n_4298)
);

HB1xp67_ASAP7_75t_L g4299 ( 
.A(n_3621),
.Y(n_4299)
);

BUFx8_ASAP7_75t_L g4300 ( 
.A(n_3859),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_3991),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4016),
.B(n_524),
.Y(n_4302)
);

OA22x2_ASAP7_75t_L g4303 ( 
.A1(n_4011),
.A2(n_3705),
.B1(n_3938),
.B2(n_3920),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_SL g4304 ( 
.A(n_3550),
.B(n_524),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_SL g4305 ( 
.A(n_3830),
.B(n_525),
.Y(n_4305)
);

O2A1O1Ixp33_ASAP7_75t_L g4306 ( 
.A1(n_3659),
.A2(n_526),
.B(n_527),
.C(n_525),
.Y(n_4306)
);

BUFx2_ASAP7_75t_L g4307 ( 
.A(n_3849),
.Y(n_4307)
);

OAI21xp33_ASAP7_75t_SL g4308 ( 
.A1(n_3598),
.A2(n_526),
.B(n_525),
.Y(n_4308)
);

INVx1_ASAP7_75t_SL g4309 ( 
.A(n_3633),
.Y(n_4309)
);

INVx2_ASAP7_75t_SL g4310 ( 
.A(n_3941),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4017),
.B(n_527),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3997),
.Y(n_4312)
);

AOI21xp5_ASAP7_75t_L g4313 ( 
.A1(n_4019),
.A2(n_529),
.B(n_528),
.Y(n_4313)
);

BUFx6f_ASAP7_75t_L g4314 ( 
.A(n_3559),
.Y(n_4314)
);

NAND2x1_ASAP7_75t_L g4315 ( 
.A(n_3655),
.B(n_3559),
.Y(n_4315)
);

OAI22xp5_ASAP7_75t_L g4316 ( 
.A1(n_3612),
.A2(n_529),
.B1(n_530),
.B2(n_528),
.Y(n_4316)
);

BUFx12f_ASAP7_75t_L g4317 ( 
.A(n_3885),
.Y(n_4317)
);

OR2x2_ASAP7_75t_L g4318 ( 
.A(n_3762),
.B(n_528),
.Y(n_4318)
);

OAI21x1_ASAP7_75t_L g4319 ( 
.A1(n_3575),
.A2(n_531),
.B(n_529),
.Y(n_4319)
);

AOI33xp33_ASAP7_75t_L g4320 ( 
.A1(n_4109),
.A2(n_62),
.A3(n_64),
.B1(n_60),
.B2(n_61),
.B3(n_63),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_SL g4321 ( 
.A(n_3830),
.B(n_531),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_3654),
.A2(n_532),
.B1(n_533),
.B2(n_531),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4085),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4088),
.B(n_533),
.Y(n_4324)
);

AOI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_3577),
.A2(n_534),
.B(n_533),
.Y(n_4325)
);

AOI21xp5_ASAP7_75t_L g4326 ( 
.A1(n_4054),
.A2(n_535),
.B(n_534),
.Y(n_4326)
);

BUFx2_ASAP7_75t_L g4327 ( 
.A(n_4008),
.Y(n_4327)
);

BUFx3_ASAP7_75t_L g4328 ( 
.A(n_3800),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4095),
.B(n_536),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3734),
.B(n_536),
.Y(n_4330)
);

AOI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_3628),
.A2(n_538),
.B(n_537),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3737),
.B(n_537),
.Y(n_4332)
);

O2A1O1Ixp33_ASAP7_75t_L g4333 ( 
.A1(n_3935),
.A2(n_539),
.B(n_540),
.C(n_537),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_SL g4334 ( 
.A(n_3774),
.B(n_4106),
.Y(n_4334)
);

OR2x6_ASAP7_75t_L g4335 ( 
.A(n_3892),
.B(n_540),
.Y(n_4335)
);

NOR2xp67_ASAP7_75t_L g4336 ( 
.A(n_3663),
.B(n_540),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_3609),
.B(n_541),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4113),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_3745),
.B(n_541),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4048),
.A2(n_542),
.B(n_541),
.Y(n_4340)
);

O2A1O1Ixp33_ASAP7_75t_L g4341 ( 
.A1(n_3697),
.A2(n_543),
.B(n_544),
.C(n_542),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3888),
.B(n_542),
.Y(n_4342)
);

OAI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_3626),
.A2(n_544),
.B(n_543),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_3625),
.B(n_545),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_3650),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3636),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_3629),
.B(n_4097),
.Y(n_4347)
);

OAI22xp5_ASAP7_75t_L g4348 ( 
.A1(n_3821),
.A2(n_546),
.B1(n_547),
.B2(n_545),
.Y(n_4348)
);

CKINVDCx16_ASAP7_75t_R g4349 ( 
.A(n_4100),
.Y(n_4349)
);

AND2x4_ASAP7_75t_L g4350 ( 
.A(n_4106),
.B(n_545),
.Y(n_4350)
);

AOI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_3673),
.A2(n_547),
.B1(n_548),
.B2(n_546),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3637),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_R g4353 ( 
.A(n_4001),
.B(n_546),
.Y(n_4353)
);

O2A1O1Ixp33_ASAP7_75t_SL g4354 ( 
.A1(n_3666),
.A2(n_1114),
.B(n_1115),
.C(n_1113),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_3751),
.B(n_3780),
.Y(n_4355)
);

NOR2xp33_ASAP7_75t_L g4356 ( 
.A(n_4013),
.B(n_549),
.Y(n_4356)
);

NOR2xp33_ASAP7_75t_L g4357 ( 
.A(n_3860),
.B(n_549),
.Y(n_4357)
);

AOI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3825),
.A2(n_550),
.B(n_549),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3786),
.B(n_550),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_3789),
.B(n_550),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_3794),
.B(n_551),
.Y(n_4361)
);

BUFx6f_ASAP7_75t_L g4362 ( 
.A(n_3590),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_3790),
.A2(n_4044),
.B(n_3630),
.Y(n_4363)
);

OAI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_3837),
.A2(n_552),
.B1(n_553),
.B2(n_551),
.Y(n_4364)
);

NOR3xp33_ASAP7_75t_SL g4365 ( 
.A(n_4099),
.B(n_1118),
.C(n_1117),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_3569),
.A2(n_552),
.B(n_551),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_3639),
.Y(n_4367)
);

INVx1_ASAP7_75t_SL g4368 ( 
.A(n_3750),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3644),
.Y(n_4369)
);

OAI21xp33_ASAP7_75t_SL g4370 ( 
.A1(n_3836),
.A2(n_553),
.B(n_552),
.Y(n_4370)
);

BUFx6f_ASAP7_75t_L g4371 ( 
.A(n_3590),
.Y(n_4371)
);

AOI21xp5_ASAP7_75t_L g4372 ( 
.A1(n_3738),
.A2(n_554),
.B(n_553),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_3817),
.B(n_554),
.Y(n_4373)
);

BUFx6f_ASAP7_75t_L g4374 ( 
.A(n_3590),
.Y(n_4374)
);

BUFx2_ASAP7_75t_L g4375 ( 
.A(n_3673),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_3739),
.B(n_1121),
.Y(n_4376)
);

OAI22xp5_ASAP7_75t_L g4377 ( 
.A1(n_3842),
.A2(n_555),
.B1(n_556),
.B2(n_554),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_3823),
.B(n_3834),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_3963),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_3850),
.B(n_555),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_SL g4381 ( 
.A(n_3761),
.B(n_4018),
.Y(n_4381)
);

CKINVDCx6p67_ASAP7_75t_R g4382 ( 
.A(n_3673),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_3728),
.A2(n_556),
.B(n_555),
.Y(n_4383)
);

A2O1A1Ixp33_ASAP7_75t_SL g4384 ( 
.A1(n_3990),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_4384)
);

INVx3_ASAP7_75t_L g4385 ( 
.A(n_4001),
.Y(n_4385)
);

OAI22xp5_ASAP7_75t_L g4386 ( 
.A1(n_3858),
.A2(n_558),
.B1(n_559),
.B2(n_557),
.Y(n_4386)
);

NOR2xp33_ASAP7_75t_R g4387 ( 
.A(n_3574),
.B(n_3578),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_3890),
.B(n_1106),
.Y(n_4388)
);

A2O1A1Ixp33_ASAP7_75t_L g4389 ( 
.A1(n_3670),
.A2(n_558),
.B(n_560),
.C(n_557),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_3646),
.Y(n_4390)
);

INVxp67_ASAP7_75t_L g4391 ( 
.A(n_4115),
.Y(n_4391)
);

O2A1O1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_4112),
.A2(n_558),
.B(n_560),
.C(n_557),
.Y(n_4392)
);

OAI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_3693),
.A2(n_561),
.B(n_560),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_3740),
.A2(n_562),
.B(n_561),
.Y(n_4394)
);

O2A1O1Ixp33_ASAP7_75t_L g4395 ( 
.A1(n_4078),
.A2(n_563),
.B(n_564),
.C(n_562),
.Y(n_4395)
);

NOR2xp33_ASAP7_75t_R g4396 ( 
.A(n_3574),
.B(n_562),
.Y(n_4396)
);

OAI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_3913),
.A2(n_565),
.B1(n_566),
.B2(n_564),
.Y(n_4397)
);

AOI21xp5_ASAP7_75t_L g4398 ( 
.A1(n_3684),
.A2(n_565),
.B(n_564),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_3865),
.B(n_566),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_3707),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_3757),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_3721),
.B(n_567),
.Y(n_4402)
);

BUFx6f_ASAP7_75t_L g4403 ( 
.A(n_3620),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_3660),
.B(n_567),
.Y(n_4404)
);

INVx1_ASAP7_75t_SL g4405 ( 
.A(n_4082),
.Y(n_4405)
);

OAI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_3726),
.A2(n_568),
.B1(n_569),
.B2(n_567),
.Y(n_4406)
);

BUFx2_ASAP7_75t_L g4407 ( 
.A(n_4083),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_3661),
.B(n_568),
.Y(n_4408)
);

BUFx8_ASAP7_75t_L g4409 ( 
.A(n_3816),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_3791),
.B(n_1119),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_3664),
.B(n_568),
.Y(n_4411)
);

OR2x6_ASAP7_75t_L g4412 ( 
.A(n_3624),
.B(n_569),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_3856),
.B(n_569),
.Y(n_4413)
);

NOR2xp33_ASAP7_75t_L g4414 ( 
.A(n_3862),
.B(n_570),
.Y(n_4414)
);

NOR2xp67_ASAP7_75t_L g4415 ( 
.A(n_3667),
.B(n_570),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_3581),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_3671),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_4018),
.B(n_571),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_3682),
.Y(n_4419)
);

NOR3xp33_ASAP7_75t_SL g4420 ( 
.A(n_4007),
.B(n_1105),
.C(n_1104),
.Y(n_4420)
);

O2A1O1Ixp33_ASAP7_75t_L g4421 ( 
.A1(n_4047),
.A2(n_573),
.B(n_574),
.C(n_572),
.Y(n_4421)
);

BUFx12f_ASAP7_75t_L g4422 ( 
.A(n_4038),
.Y(n_4422)
);

NOR3xp33_ASAP7_75t_L g4423 ( 
.A(n_3998),
.B(n_573),
.C(n_572),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_3592),
.Y(n_4424)
);

O2A1O1Ixp33_ASAP7_75t_L g4425 ( 
.A1(n_3562),
.A2(n_574),
.B(n_575),
.C(n_572),
.Y(n_4425)
);

AOI21x1_ASAP7_75t_L g4426 ( 
.A1(n_3932),
.A2(n_575),
.B(n_574),
.Y(n_4426)
);

BUFx3_ASAP7_75t_L g4427 ( 
.A(n_4116),
.Y(n_4427)
);

AO21x1_ASAP7_75t_L g4428 ( 
.A1(n_3771),
.A2(n_577),
.B(n_576),
.Y(n_4428)
);

A2O1A1Ixp33_ASAP7_75t_L g4429 ( 
.A1(n_3674),
.A2(n_577),
.B(n_578),
.C(n_576),
.Y(n_4429)
);

OAI22xp5_ASAP7_75t_L g4430 ( 
.A1(n_3760),
.A2(n_577),
.B1(n_578),
.B2(n_576),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_3578),
.B(n_579),
.Y(n_4431)
);

NOR2xp33_ASAP7_75t_L g4432 ( 
.A(n_4084),
.B(n_579),
.Y(n_4432)
);

AND2x4_ASAP7_75t_L g4433 ( 
.A(n_3579),
.B(n_580),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_3715),
.B(n_580),
.Y(n_4434)
);

A2O1A1Ixp33_ASAP7_75t_SL g4435 ( 
.A1(n_3741),
.A2(n_3770),
.B(n_3909),
.C(n_3896),
.Y(n_4435)
);

AOI22x1_ASAP7_75t_L g4436 ( 
.A1(n_3552),
.A2(n_582),
.B1(n_583),
.B2(n_581),
.Y(n_4436)
);

AOI21xp5_ASAP7_75t_L g4437 ( 
.A1(n_3689),
.A2(n_582),
.B(n_581),
.Y(n_4437)
);

INVx3_ASAP7_75t_SL g4438 ( 
.A(n_3791),
.Y(n_4438)
);

A2O1A1Ixp33_ASAP7_75t_L g4439 ( 
.A1(n_3714),
.A2(n_582),
.B(n_583),
.C(n_581),
.Y(n_4439)
);

INVx4_ASAP7_75t_L g4440 ( 
.A(n_3619),
.Y(n_4440)
);

BUFx2_ASAP7_75t_L g4441 ( 
.A(n_3915),
.Y(n_4441)
);

A2O1A1Ixp33_ASAP7_75t_L g4442 ( 
.A1(n_3718),
.A2(n_585),
.B(n_586),
.C(n_584),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_3560),
.B(n_584),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3696),
.Y(n_4444)
);

AOI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_3727),
.A2(n_585),
.B(n_584),
.Y(n_4445)
);

HB1xp67_ASAP7_75t_L g4446 ( 
.A(n_3958),
.Y(n_4446)
);

INVx1_ASAP7_75t_SL g4447 ( 
.A(n_4029),
.Y(n_4447)
);

AOI21xp5_ASAP7_75t_L g4448 ( 
.A1(n_3731),
.A2(n_587),
.B(n_586),
.Y(n_4448)
);

OR2x2_ASAP7_75t_L g4449 ( 
.A(n_3554),
.B(n_587),
.Y(n_4449)
);

AO32x1_ASAP7_75t_L g4450 ( 
.A1(n_4003),
.A2(n_590),
.A3(n_591),
.B1(n_589),
.B2(n_588),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_3564),
.B(n_588),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_3701),
.Y(n_4452)
);

AOI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_3642),
.A2(n_3778),
.B(n_3772),
.Y(n_4453)
);

AO32x1_ASAP7_75t_L g4454 ( 
.A1(n_3556),
.A2(n_591),
.A3(n_592),
.B1(n_590),
.B2(n_589),
.Y(n_4454)
);

NOR2xp33_ASAP7_75t_L g4455 ( 
.A(n_3912),
.B(n_589),
.Y(n_4455)
);

OAI22xp5_ASAP7_75t_L g4456 ( 
.A1(n_3545),
.A2(n_591),
.B1(n_592),
.B2(n_590),
.Y(n_4456)
);

OAI22xp5_ASAP7_75t_L g4457 ( 
.A1(n_3881),
.A2(n_593),
.B1(n_594),
.B2(n_592),
.Y(n_4457)
);

INVx4_ASAP7_75t_L g4458 ( 
.A(n_3619),
.Y(n_4458)
);

INVx5_ASAP7_75t_L g4459 ( 
.A(n_3620),
.Y(n_4459)
);

BUFx2_ASAP7_75t_L g4460 ( 
.A(n_3965),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_SL g4461 ( 
.A(n_4034),
.B(n_593),
.Y(n_4461)
);

OAI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_3632),
.A2(n_595),
.B1(n_596),
.B2(n_594),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_3788),
.Y(n_4463)
);

AOI21xp5_ASAP7_75t_L g4464 ( 
.A1(n_3832),
.A2(n_595),
.B(n_594),
.Y(n_4464)
);

O2A1O1Ixp33_ASAP7_75t_L g4465 ( 
.A1(n_3781),
.A2(n_596),
.B(n_597),
.C(n_595),
.Y(n_4465)
);

INVxp67_ASAP7_75t_L g4466 ( 
.A(n_3724),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4089),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_3878),
.A2(n_597),
.B1(n_598),
.B2(n_596),
.Y(n_4468)
);

OAI22xp5_ASAP7_75t_L g4469 ( 
.A1(n_4096),
.A2(n_600),
.B1(n_601),
.B2(n_599),
.Y(n_4469)
);

NOR2xp33_ASAP7_75t_L g4470 ( 
.A(n_3631),
.B(n_599),
.Y(n_4470)
);

INVx2_ASAP7_75t_L g4471 ( 
.A(n_3893),
.Y(n_4471)
);

AND2x4_ASAP7_75t_L g4472 ( 
.A(n_3579),
.B(n_600),
.Y(n_4472)
);

NOR2xp33_ASAP7_75t_L g4473 ( 
.A(n_3640),
.B(n_600),
.Y(n_4473)
);

INVxp67_ASAP7_75t_SL g4474 ( 
.A(n_3620),
.Y(n_4474)
);

OAI22xp5_ASAP7_75t_L g4475 ( 
.A1(n_4111),
.A2(n_602),
.B1(n_603),
.B2(n_601),
.Y(n_4475)
);

NOR2xp33_ASAP7_75t_L g4476 ( 
.A(n_3735),
.B(n_601),
.Y(n_4476)
);

OR2x6_ASAP7_75t_L g4477 ( 
.A(n_4090),
.B(n_602),
.Y(n_4477)
);

OR2x6_ASAP7_75t_L g4478 ( 
.A(n_3657),
.B(n_603),
.Y(n_4478)
);

AND2x2_ASAP7_75t_SL g4479 ( 
.A(n_3981),
.B(n_603),
.Y(n_4479)
);

AND2x2_ASAP7_75t_SL g4480 ( 
.A(n_3981),
.B(n_604),
.Y(n_4480)
);

INVx2_ASAP7_75t_SL g4481 ( 
.A(n_4037),
.Y(n_4481)
);

A2O1A1Ixp33_ASAP7_75t_L g4482 ( 
.A1(n_3725),
.A2(n_605),
.B(n_606),
.C(n_604),
.Y(n_4482)
);

NOR2xp33_ASAP7_75t_L g4483 ( 
.A(n_3769),
.B(n_605),
.Y(n_4483)
);

AND2x6_ASAP7_75t_L g4484 ( 
.A(n_3657),
.B(n_605),
.Y(n_4484)
);

OAI22xp5_ASAP7_75t_L g4485 ( 
.A1(n_3884),
.A2(n_607),
.B1(n_608),
.B2(n_606),
.Y(n_4485)
);

BUFx2_ASAP7_75t_L g4486 ( 
.A(n_4034),
.Y(n_4486)
);

HB1xp67_ASAP7_75t_L g4487 ( 
.A(n_4037),
.Y(n_4487)
);

O2A1O1Ixp33_ASAP7_75t_L g4488 ( 
.A1(n_3754),
.A2(n_607),
.B(n_608),
.C(n_606),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_3847),
.A2(n_609),
.B(n_608),
.Y(n_4489)
);

AND2x4_ASAP7_75t_L g4490 ( 
.A(n_3665),
.B(n_3744),
.Y(n_4490)
);

AOI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_3926),
.A2(n_610),
.B(n_609),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_3567),
.B(n_609),
.Y(n_4492)
);

AOI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_3962),
.A2(n_612),
.B(n_611),
.Y(n_4493)
);

AOI21x1_ASAP7_75t_L g4494 ( 
.A1(n_3905),
.A2(n_612),
.B(n_611),
.Y(n_4494)
);

BUFx8_ASAP7_75t_L g4495 ( 
.A(n_4104),
.Y(n_4495)
);

OAI22xp5_ASAP7_75t_L g4496 ( 
.A1(n_3927),
.A2(n_614),
.B1(n_616),
.B2(n_613),
.Y(n_4496)
);

AOI22xp33_ASAP7_75t_L g4497 ( 
.A1(n_4022),
.A2(n_616),
.B1(n_617),
.B2(n_613),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_3897),
.Y(n_4498)
);

OAI22xp5_ASAP7_75t_L g4499 ( 
.A1(n_3940),
.A2(n_616),
.B1(n_617),
.B2(n_613),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4020),
.A2(n_3568),
.B1(n_3580),
.B2(n_3572),
.Y(n_4500)
);

O2A1O1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_3871),
.A2(n_618),
.B(n_619),
.C(n_617),
.Y(n_4501)
);

OAI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_3583),
.A2(n_619),
.B1(n_620),
.B2(n_618),
.Y(n_4502)
);

A2O1A1Ixp33_ASAP7_75t_L g4503 ( 
.A1(n_3733),
.A2(n_619),
.B(n_620),
.C(n_618),
.Y(n_4503)
);

NAND3xp33_ASAP7_75t_SL g4504 ( 
.A(n_3763),
.B(n_60),
.C(n_61),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_3711),
.Y(n_4505)
);

OR2x6_ASAP7_75t_L g4506 ( 
.A(n_3665),
.B(n_620),
.Y(n_4506)
);

AOI21xp5_ASAP7_75t_L g4507 ( 
.A1(n_3974),
.A2(n_622),
.B(n_621),
.Y(n_4507)
);

NAND3xp33_ASAP7_75t_L g4508 ( 
.A(n_3752),
.B(n_1105),
.C(n_1104),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_SL g4509 ( 
.A(n_3722),
.B(n_621),
.Y(n_4509)
);

NOR2xp67_ASAP7_75t_L g4510 ( 
.A(n_4040),
.B(n_622),
.Y(n_4510)
);

AOI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_3980),
.A2(n_624),
.B(n_623),
.Y(n_4511)
);

NOR2x1_ASAP7_75t_L g4512 ( 
.A(n_3744),
.B(n_623),
.Y(n_4512)
);

INVx2_ASAP7_75t_SL g4513 ( 
.A(n_3808),
.Y(n_4513)
);

NOR2xp33_ASAP7_75t_SL g4514 ( 
.A(n_3808),
.B(n_624),
.Y(n_4514)
);

AOI21x1_ASAP7_75t_L g4515 ( 
.A1(n_3984),
.A2(n_625),
.B(n_624),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_R g4516 ( 
.A(n_3895),
.B(n_625),
.Y(n_4516)
);

BUFx6f_ASAP7_75t_L g4517 ( 
.A(n_3722),
.Y(n_4517)
);

NOR2xp33_ASAP7_75t_R g4518 ( 
.A(n_3895),
.B(n_3961),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_3589),
.B(n_625),
.Y(n_4519)
);

O2A1O1Ixp33_ASAP7_75t_L g4520 ( 
.A1(n_4068),
.A2(n_627),
.B(n_628),
.C(n_626),
.Y(n_4520)
);

O2A1O1Ixp33_ASAP7_75t_SL g4521 ( 
.A1(n_3966),
.A2(n_1110),
.B(n_1111),
.C(n_1109),
.Y(n_4521)
);

INVx3_ASAP7_75t_L g4522 ( 
.A(n_4040),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_3986),
.A2(n_627),
.B(n_626),
.Y(n_4523)
);

OR2x6_ASAP7_75t_L g4524 ( 
.A(n_3563),
.B(n_626),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3992),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_3900),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_SL g4527 ( 
.A(n_3722),
.B(n_627),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_SL g4528 ( 
.A(n_3749),
.B(n_3773),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_3911),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3995),
.Y(n_4530)
);

OR2x2_ASAP7_75t_L g4531 ( 
.A(n_3596),
.B(n_628),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_3994),
.A2(n_630),
.B(n_629),
.Y(n_4532)
);

AOI22xp5_ASAP7_75t_L g4533 ( 
.A1(n_3802),
.A2(n_630),
.B1(n_631),
.B2(n_629),
.Y(n_4533)
);

AOI221xp5_ASAP7_75t_L g4534 ( 
.A1(n_4086),
.A2(n_632),
.B1(n_633),
.B2(n_631),
.C(n_630),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4032),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_3914),
.Y(n_4536)
);

AOI21xp5_ASAP7_75t_L g4537 ( 
.A1(n_4012),
.A2(n_633),
.B(n_632),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_3919),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_3601),
.B(n_3602),
.Y(n_4539)
);

INVx5_ASAP7_75t_L g4540 ( 
.A(n_3749),
.Y(n_4540)
);

A2O1A1Ixp33_ASAP7_75t_SL g4541 ( 
.A1(n_3747),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_4541)
);

AOI221xp5_ASAP7_75t_SL g4542 ( 
.A1(n_4049),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_4542)
);

AOI21x1_ASAP7_75t_L g4543 ( 
.A1(n_4026),
.A2(n_633),
.B(n_632),
.Y(n_4543)
);

OR2x2_ASAP7_75t_L g4544 ( 
.A(n_3604),
.B(n_634),
.Y(n_4544)
);

OA22x2_ASAP7_75t_L g4545 ( 
.A1(n_3976),
.A2(n_635),
.B1(n_636),
.B2(n_634),
.Y(n_4545)
);

AOI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_3606),
.A2(n_635),
.B(n_634),
.Y(n_4546)
);

A2O1A1Ixp33_ASAP7_75t_L g4547 ( 
.A1(n_3746),
.A2(n_637),
.B(n_638),
.C(n_636),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_4027),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4036),
.Y(n_4549)
);

AO21x2_ASAP7_75t_L g4550 ( 
.A1(n_3946),
.A2(n_637),
.B(n_636),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_3811),
.B(n_3835),
.Y(n_4551)
);

AND2x4_ASAP7_75t_L g4552 ( 
.A(n_3961),
.B(n_637),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_3712),
.B(n_638),
.Y(n_4553)
);

AOI21xp5_ASAP7_75t_L g4554 ( 
.A1(n_3880),
.A2(n_639),
.B(n_638),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4045),
.B(n_639),
.Y(n_4555)
);

CKINVDCx16_ASAP7_75t_R g4556 ( 
.A(n_4079),
.Y(n_4556)
);

NOR2x1_ASAP7_75t_R g4557 ( 
.A(n_4062),
.B(n_639),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_3922),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_3846),
.B(n_1111),
.Y(n_4559)
);

OR2x6_ASAP7_75t_SL g4560 ( 
.A(n_3695),
.B(n_3845),
.Y(n_4560)
);

BUFx2_ASAP7_75t_L g4561 ( 
.A(n_3977),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4056),
.B(n_1112),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_3924),
.Y(n_4563)
);

OAI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_3857),
.A2(n_641),
.B(n_640),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_SL g4565 ( 
.A(n_3749),
.B(n_640),
.Y(n_4565)
);

OAI21xp33_ASAP7_75t_L g4566 ( 
.A1(n_4098),
.A2(n_63),
.B(n_64),
.Y(n_4566)
);

INVx2_ASAP7_75t_SL g4567 ( 
.A(n_4027),
.Y(n_4567)
);

A2O1A1Ixp33_ASAP7_75t_L g4568 ( 
.A1(n_4050),
.A2(n_641),
.B(n_642),
.C(n_640),
.Y(n_4568)
);

O2A1O1Ixp33_ASAP7_75t_L g4569 ( 
.A1(n_4061),
.A2(n_642),
.B(n_643),
.C(n_641),
.Y(n_4569)
);

BUFx4f_ASAP7_75t_SL g4570 ( 
.A(n_4030),
.Y(n_4570)
);

AOI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4055),
.A2(n_645),
.B1(n_646),
.B2(n_643),
.Y(n_4571)
);

NAND2x1p5_ASAP7_75t_L g4572 ( 
.A(n_3773),
.B(n_3777),
.Y(n_4572)
);

BUFx6f_ASAP7_75t_L g4573 ( 
.A(n_3773),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_3928),
.Y(n_4574)
);

AND2x4_ASAP7_75t_L g4575 ( 
.A(n_3977),
.B(n_643),
.Y(n_4575)
);

AOI21xp5_ASAP7_75t_L g4576 ( 
.A1(n_3720),
.A2(n_646),
.B(n_645),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_3937),
.Y(n_4577)
);

NOR2xp33_ASAP7_75t_L g4578 ( 
.A(n_3979),
.B(n_645),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_SL g4579 ( 
.A(n_3777),
.B(n_647),
.Y(n_4579)
);

AOI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_3873),
.A2(n_648),
.B1(n_649),
.B2(n_647),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_SL g4581 ( 
.A(n_3777),
.B(n_3875),
.Y(n_4581)
);

AOI21xp5_ASAP7_75t_L g4582 ( 
.A1(n_4059),
.A2(n_648),
.B(n_647),
.Y(n_4582)
);

INVx2_ASAP7_75t_L g4583 ( 
.A(n_3944),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_3952),
.Y(n_4584)
);

NOR2xp33_ASAP7_75t_L g4585 ( 
.A(n_3985),
.B(n_648),
.Y(n_4585)
);

AO32x1_ASAP7_75t_L g4586 ( 
.A1(n_4041),
.A2(n_651),
.A3(n_652),
.B1(n_650),
.B2(n_649),
.Y(n_4586)
);

AOI21xp5_ASAP7_75t_L g4587 ( 
.A1(n_3852),
.A2(n_650),
.B(n_649),
.Y(n_4587)
);

O2A1O1Ixp33_ASAP7_75t_L g4588 ( 
.A1(n_3814),
.A2(n_651),
.B(n_652),
.C(n_650),
.Y(n_4588)
);

OAI22xp5_ASAP7_75t_L g4589 ( 
.A1(n_3949),
.A2(n_653),
.B1(n_654),
.B2(n_651),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4069),
.B(n_653),
.Y(n_4590)
);

AOI21xp5_ASAP7_75t_L g4591 ( 
.A1(n_3584),
.A2(n_3591),
.B(n_3875),
.Y(n_4591)
);

AOI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_3875),
.A2(n_654),
.B(n_653),
.Y(n_4592)
);

NOR3xp33_ASAP7_75t_SL g4593 ( 
.A(n_3676),
.B(n_1112),
.C(n_1109),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4039),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4070),
.B(n_4102),
.Y(n_4595)
);

NOR2xp33_ASAP7_75t_R g4596 ( 
.A(n_3939),
.B(n_655),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_3939),
.A2(n_4006),
.B(n_3993),
.Y(n_4597)
);

NAND2x1_ASAP7_75t_L g4598 ( 
.A(n_3939),
.B(n_655),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_3953),
.Y(n_4599)
);

NOR2xp33_ASAP7_75t_L g4600 ( 
.A(n_4030),
.B(n_655),
.Y(n_4600)
);

OAI22xp5_ASAP7_75t_L g4601 ( 
.A1(n_3950),
.A2(n_657),
.B1(n_658),
.B2(n_656),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_SL g4602 ( 
.A(n_4006),
.B(n_656),
.Y(n_4602)
);

OAI22xp5_ASAP7_75t_L g4603 ( 
.A1(n_3954),
.A2(n_658),
.B1(n_659),
.B2(n_657),
.Y(n_4603)
);

AOI21xp5_ASAP7_75t_L g4604 ( 
.A1(n_4006),
.A2(n_658),
.B(n_657),
.Y(n_4604)
);

BUFx2_ASAP7_75t_L g4605 ( 
.A(n_4104),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_3955),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4057),
.B(n_659),
.Y(n_4607)
);

AOI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_4035),
.A2(n_661),
.B(n_660),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_3959),
.Y(n_4609)
);

NOR2xp33_ASAP7_75t_L g4610 ( 
.A(n_4025),
.B(n_660),
.Y(n_4610)
);

AND2x6_ASAP7_75t_L g4611 ( 
.A(n_4104),
.B(n_661),
.Y(n_4611)
);

HB1xp67_ASAP7_75t_L g4612 ( 
.A(n_4073),
.Y(n_4612)
);

HB1xp67_ASAP7_75t_L g4613 ( 
.A(n_3775),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_3776),
.B(n_662),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_3784),
.B(n_662),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_3907),
.Y(n_4616)
);

A2O1A1Ixp33_ASAP7_75t_L g4617 ( 
.A1(n_3982),
.A2(n_4114),
.B(n_4063),
.C(n_3874),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_3923),
.Y(n_4618)
);

AOI21x1_ASAP7_75t_L g4619 ( 
.A1(n_4033),
.A2(n_663),
.B(n_662),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_3570),
.Y(n_4620)
);

BUFx2_ASAP7_75t_SL g4621 ( 
.A(n_4042),
.Y(n_4621)
);

BUFx6f_ASAP7_75t_L g4622 ( 
.A(n_4077),
.Y(n_4622)
);

AOI22xp5_ASAP7_75t_L g4623 ( 
.A1(n_3785),
.A2(n_664),
.B1(n_665),
.B2(n_663),
.Y(n_4623)
);

AND3x2_ASAP7_75t_L g4624 ( 
.A(n_3582),
.B(n_664),
.C(n_663),
.Y(n_4624)
);

CKINVDCx6p67_ASAP7_75t_R g4625 ( 
.A(n_3901),
.Y(n_4625)
);

AOI21xp5_ASAP7_75t_L g4626 ( 
.A1(n_3686),
.A2(n_666),
.B(n_665),
.Y(n_4626)
);

HB1xp67_ASAP7_75t_L g4627 ( 
.A(n_4043),
.Y(n_4627)
);

OAI22xp5_ASAP7_75t_L g4628 ( 
.A1(n_3916),
.A2(n_666),
.B1(n_667),
.B2(n_665),
.Y(n_4628)
);

AND2x4_ASAP7_75t_L g4629 ( 
.A(n_3795),
.B(n_666),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_3945),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_3782),
.B(n_667),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_3799),
.B(n_667),
.Y(n_4632)
);

AOI22xp5_ASAP7_75t_L g4633 ( 
.A1(n_3948),
.A2(n_669),
.B1(n_670),
.B2(n_668),
.Y(n_4633)
);

NOR3xp33_ASAP7_75t_SL g4634 ( 
.A(n_3803),
.B(n_1107),
.C(n_1106),
.Y(n_4634)
);

AOI21xp5_ASAP7_75t_L g4635 ( 
.A1(n_3690),
.A2(n_669),
.B(n_668),
.Y(n_4635)
);

AOI21xp5_ASAP7_75t_L g4636 ( 
.A1(n_3691),
.A2(n_669),
.B(n_668),
.Y(n_4636)
);

OAI22xp5_ASAP7_75t_L g4637 ( 
.A1(n_4004),
.A2(n_671),
.B1(n_673),
.B2(n_670),
.Y(n_4637)
);

INVx4_ASAP7_75t_L g4638 ( 
.A(n_4005),
.Y(n_4638)
);

OAI22xp5_ASAP7_75t_L g4639 ( 
.A1(n_4014),
.A2(n_671),
.B1(n_673),
.B2(n_670),
.Y(n_4639)
);

AOI21xp5_ASAP7_75t_L g4640 ( 
.A1(n_3806),
.A2(n_675),
.B(n_674),
.Y(n_4640)
);

A2O1A1Ixp33_ASAP7_75t_SL g4641 ( 
.A1(n_3801),
.A2(n_66),
.B(n_63),
.C(n_65),
.Y(n_4641)
);

OAI22x1_ASAP7_75t_L g4642 ( 
.A1(n_3809),
.A2(n_675),
.B1(n_676),
.B2(n_674),
.Y(n_4642)
);

AOI21xp5_ASAP7_75t_L g4643 ( 
.A1(n_3807),
.A2(n_676),
.B(n_675),
.Y(n_4643)
);

INVx6_ASAP7_75t_L g4644 ( 
.A(n_3861),
.Y(n_4644)
);

OR2x6_ASAP7_75t_L g4645 ( 
.A(n_4015),
.B(n_676),
.Y(n_4645)
);

BUFx6f_ASAP7_75t_L g4646 ( 
.A(n_4064),
.Y(n_4646)
);

AOI21xp5_ASAP7_75t_L g4647 ( 
.A1(n_3812),
.A2(n_678),
.B(n_677),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_SL g4648 ( 
.A(n_3815),
.B(n_677),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_3822),
.B(n_679),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_3829),
.Y(n_4650)
);

INVx3_ASAP7_75t_L g4651 ( 
.A(n_4023),
.Y(n_4651)
);

BUFx6f_ASAP7_75t_L g4652 ( 
.A(n_3700),
.Y(n_4652)
);

INVx3_ASAP7_75t_L g4653 ( 
.A(n_4024),
.Y(n_4653)
);

NOR3xp33_ASAP7_75t_L g4654 ( 
.A(n_3933),
.B(n_680),
.C(n_679),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_3947),
.Y(n_4655)
);

O2A1O1Ixp33_ASAP7_75t_L g4656 ( 
.A1(n_3838),
.A2(n_680),
.B(n_681),
.C(n_679),
.Y(n_4656)
);

AO22x1_ASAP7_75t_L g4657 ( 
.A1(n_4052),
.A2(n_682),
.B1(n_683),
.B2(n_681),
.Y(n_4657)
);

BUFx4f_ASAP7_75t_L g4658 ( 
.A(n_4108),
.Y(n_4658)
);

AOI21xp5_ASAP7_75t_L g4659 ( 
.A1(n_3839),
.A2(n_683),
.B(n_682),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_3840),
.B(n_682),
.Y(n_4660)
);

AOI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_3956),
.A2(n_684),
.B1(n_685),
.B2(n_683),
.Y(n_4661)
);

OAI22xp5_ASAP7_75t_L g4662 ( 
.A1(n_3957),
.A2(n_685),
.B1(n_686),
.B2(n_684),
.Y(n_4662)
);

NAND3xp33_ASAP7_75t_L g4663 ( 
.A(n_3841),
.B(n_1108),
.C(n_1107),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_SL g4664 ( 
.A(n_3853),
.B(n_684),
.Y(n_4664)
);

O2A1O1Ixp33_ASAP7_75t_L g4665 ( 
.A1(n_3867),
.A2(n_686),
.B(n_687),
.C(n_685),
.Y(n_4665)
);

INVx4_ASAP7_75t_L g4666 ( 
.A(n_3876),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_3877),
.Y(n_4667)
);

A2O1A1Ixp33_ASAP7_75t_SL g4668 ( 
.A1(n_3879),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_4668)
);

NOR2xp33_ASAP7_75t_R g4669 ( 
.A(n_3882),
.B(n_686),
.Y(n_4669)
);

AOI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_3889),
.A2(n_688),
.B(n_687),
.Y(n_4670)
);

NOR2xp67_ASAP7_75t_SL g4671 ( 
.A(n_3792),
.B(n_688),
.Y(n_4671)
);

BUFx3_ASAP7_75t_L g4672 ( 
.A(n_4071),
.Y(n_4672)
);

OR2x2_ASAP7_75t_L g4673 ( 
.A(n_3891),
.B(n_689),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_SL g4674 ( 
.A(n_3793),
.B(n_689),
.Y(n_4674)
);

INVx3_ASAP7_75t_L g4675 ( 
.A(n_3614),
.Y(n_4675)
);

A2O1A1Ixp33_ASAP7_75t_L g4676 ( 
.A1(n_3645),
.A2(n_690),
.B(n_691),
.C(n_689),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_3931),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_3694),
.B(n_1100),
.Y(n_4678)
);

INVx4_ASAP7_75t_L g4679 ( 
.A(n_3967),
.Y(n_4679)
);

INVx4_ASAP7_75t_L g4680 ( 
.A(n_3968),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_3942),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4376),
.B(n_4281),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4122),
.B(n_3969),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4123),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4148),
.Y(n_4685)
);

AOI21xp5_ASAP7_75t_L g4686 ( 
.A1(n_4134),
.A2(n_3702),
.B(n_4067),
.Y(n_4686)
);

BUFx3_ASAP7_75t_L g4687 ( 
.A(n_4247),
.Y(n_4687)
);

AOI21x1_ASAP7_75t_L g4688 ( 
.A1(n_4194),
.A2(n_4060),
.B(n_3943),
.Y(n_4688)
);

OAI21x1_ASAP7_75t_L g4689 ( 
.A1(n_4597),
.A2(n_4075),
.B(n_4074),
.Y(n_4689)
);

AOI21x1_ASAP7_75t_L g4690 ( 
.A1(n_4426),
.A2(n_3988),
.B(n_3649),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4226),
.B(n_3647),
.Y(n_4691)
);

BUFx12f_ASAP7_75t_L g4692 ( 
.A(n_4135),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4150),
.Y(n_4693)
);

AO31x2_ASAP7_75t_L g4694 ( 
.A1(n_4416),
.A2(n_4080),
.A3(n_4093),
.B(n_4092),
.Y(n_4694)
);

AOI22xp5_ASAP7_75t_L g4695 ( 
.A1(n_4479),
.A2(n_3681),
.B1(n_3668),
.B2(n_3999),
.Y(n_4695)
);

OAI21x1_ASAP7_75t_L g4696 ( 
.A1(n_4379),
.A2(n_4107),
.B(n_4094),
.Y(n_4696)
);

OAI21xp5_ASAP7_75t_L g4697 ( 
.A1(n_4146),
.A2(n_3685),
.B(n_691),
.Y(n_4697)
);

BUFx6f_ASAP7_75t_L g4698 ( 
.A(n_4277),
.Y(n_4698)
);

OAI21x1_ASAP7_75t_L g4699 ( 
.A1(n_4591),
.A2(n_4401),
.B(n_4400),
.Y(n_4699)
);

OAI21xp5_ASAP7_75t_L g4700 ( 
.A1(n_4172),
.A2(n_691),
.B(n_690),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4154),
.Y(n_4701)
);

A2O1A1Ixp33_ASAP7_75t_L g4702 ( 
.A1(n_4415),
.A2(n_4297),
.B(n_4336),
.C(n_4365),
.Y(n_4702)
);

OAI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4143),
.A2(n_692),
.B(n_690),
.Y(n_4703)
);

OA21x2_ASAP7_75t_L g4704 ( 
.A1(n_4424),
.A2(n_693),
.B(n_692),
.Y(n_4704)
);

A2O1A1Ixp33_ASAP7_75t_L g4705 ( 
.A1(n_4308),
.A2(n_693),
.B(n_694),
.C(n_692),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4235),
.B(n_693),
.Y(n_4706)
);

AOI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4130),
.A2(n_695),
.B(n_694),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4220),
.Y(n_4708)
);

AND3x4_ASAP7_75t_L g4709 ( 
.A(n_4197),
.B(n_697),
.C(n_696),
.Y(n_4709)
);

AOI21xp5_ASAP7_75t_L g4710 ( 
.A1(n_4363),
.A2(n_698),
.B(n_696),
.Y(n_4710)
);

AOI21xp5_ASAP7_75t_L g4711 ( 
.A1(n_4528),
.A2(n_4581),
.B(n_4435),
.Y(n_4711)
);

A2O1A1Ixp33_ASAP7_75t_L g4712 ( 
.A1(n_4341),
.A2(n_698),
.B(n_699),
.C(n_696),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4126),
.Y(n_4713)
);

AOI21xp5_ASAP7_75t_L g4714 ( 
.A1(n_4453),
.A2(n_699),
.B(n_698),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4267),
.B(n_4229),
.Y(n_4715)
);

OA21x2_ASAP7_75t_L g4716 ( 
.A1(n_4467),
.A2(n_700),
.B(n_699),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4156),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4246),
.B(n_700),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4259),
.B(n_4275),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_4293),
.B(n_4276),
.Y(n_4720)
);

AO21x1_ASAP7_75t_L g4721 ( 
.A1(n_4381),
.A2(n_701),
.B(n_700),
.Y(n_4721)
);

NOR4xp25_ASAP7_75t_L g4722 ( 
.A(n_4320),
.B(n_702),
.C(n_703),
.D(n_701),
.Y(n_4722)
);

AOI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4480),
.A2(n_1119),
.B1(n_1120),
.B2(n_1117),
.Y(n_4723)
);

OAI21x1_ASAP7_75t_L g4724 ( 
.A1(n_4463),
.A2(n_703),
.B(n_702),
.Y(n_4724)
);

INVx5_ASAP7_75t_L g4725 ( 
.A(n_4135),
.Y(n_4725)
);

NAND2xp33_ASAP7_75t_SL g4726 ( 
.A(n_4596),
.B(n_702),
.Y(n_4726)
);

OAI21x1_ASAP7_75t_L g4727 ( 
.A1(n_4203),
.A2(n_704),
.B(n_703),
.Y(n_4727)
);

OR2x2_ASAP7_75t_L g4728 ( 
.A(n_4167),
.B(n_704),
.Y(n_4728)
);

NOR2xp33_ASAP7_75t_SL g4729 ( 
.A(n_4135),
.B(n_704),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4141),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4162),
.B(n_705),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_L g4732 ( 
.A1(n_4191),
.A2(n_706),
.B(n_705),
.Y(n_4732)
);

AOI21xp5_ASAP7_75t_L g4733 ( 
.A1(n_4152),
.A2(n_706),
.B(n_705),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4182),
.B(n_4198),
.Y(n_4734)
);

OAI21x1_ASAP7_75t_L g4735 ( 
.A1(n_4196),
.A2(n_707),
.B(n_706),
.Y(n_4735)
);

OR2x2_ASAP7_75t_L g4736 ( 
.A(n_4202),
.B(n_707),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4201),
.Y(n_4737)
);

AOI21xp5_ASAP7_75t_L g4738 ( 
.A1(n_4500),
.A2(n_708),
.B(n_707),
.Y(n_4738)
);

BUFx2_ASAP7_75t_L g4739 ( 
.A(n_4495),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4145),
.Y(n_4740)
);

A2O1A1Ixp33_ASAP7_75t_L g4741 ( 
.A1(n_4588),
.A2(n_709),
.B(n_710),
.C(n_708),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4345),
.B(n_709),
.Y(n_4742)
);

OAI22xp5_ASAP7_75t_L g4743 ( 
.A1(n_4382),
.A2(n_4187),
.B1(n_4375),
.B2(n_4560),
.Y(n_4743)
);

OAI21x1_ASAP7_75t_L g4744 ( 
.A1(n_4164),
.A2(n_711),
.B(n_710),
.Y(n_4744)
);

OAI21x1_ASAP7_75t_L g4745 ( 
.A1(n_4651),
.A2(n_712),
.B(n_711),
.Y(n_4745)
);

OAI21x1_ASAP7_75t_L g4746 ( 
.A1(n_4653),
.A2(n_713),
.B(n_712),
.Y(n_4746)
);

OA21x2_ASAP7_75t_L g4747 ( 
.A1(n_4319),
.A2(n_713),
.B(n_712),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_SL g4748 ( 
.A1(n_4440),
.A2(n_715),
.B(n_714),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4118),
.B(n_4268),
.Y(n_4749)
);

AND2x2_ASAP7_75t_L g4750 ( 
.A(n_4298),
.B(n_4337),
.Y(n_4750)
);

AOI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4178),
.A2(n_715),
.B(n_714),
.Y(n_4751)
);

OAI21xp33_ASAP7_75t_L g4752 ( 
.A1(n_4149),
.A2(n_716),
.B(n_714),
.Y(n_4752)
);

AO31x2_ASAP7_75t_L g4753 ( 
.A1(n_4679),
.A2(n_717),
.A3(n_718),
.B(n_716),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4211),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4323),
.B(n_716),
.Y(n_4755)
);

NOR2xp33_ASAP7_75t_L g4756 ( 
.A(n_4257),
.B(n_717),
.Y(n_4756)
);

OAI22x1_ASAP7_75t_L g4757 ( 
.A1(n_4438),
.A2(n_4125),
.B1(n_4206),
.B2(n_4184),
.Y(n_4757)
);

INVx2_ASAP7_75t_L g4758 ( 
.A(n_4168),
.Y(n_4758)
);

A2O1A1Ixp33_ASAP7_75t_L g4759 ( 
.A1(n_4465),
.A2(n_719),
.B(n_720),
.C(n_717),
.Y(n_4759)
);

INVx2_ASAP7_75t_SL g4760 ( 
.A(n_4300),
.Y(n_4760)
);

NAND2xp33_ASAP7_75t_L g4761 ( 
.A(n_4353),
.B(n_719),
.Y(n_4761)
);

OAI21xp33_ASAP7_75t_L g4762 ( 
.A1(n_4303),
.A2(n_721),
.B(n_720),
.Y(n_4762)
);

A2O1A1Ixp33_ASAP7_75t_L g4763 ( 
.A1(n_4569),
.A2(n_722),
.B(n_723),
.C(n_721),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4294),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4190),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4346),
.B(n_721),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4352),
.B(n_722),
.Y(n_4767)
);

AOI221xp5_ASAP7_75t_SL g4768 ( 
.A1(n_4140),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4367),
.B(n_722),
.Y(n_4769)
);

OAI21x1_ASAP7_75t_L g4770 ( 
.A1(n_4572),
.A2(n_724),
.B(n_723),
.Y(n_4770)
);

INVxp67_ASAP7_75t_SL g4771 ( 
.A(n_4487),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4369),
.B(n_723),
.Y(n_4772)
);

A2O1A1Ixp33_ASAP7_75t_L g4773 ( 
.A1(n_4333),
.A2(n_725),
.B(n_726),
.C(n_724),
.Y(n_4773)
);

OAI21x1_ASAP7_75t_L g4774 ( 
.A1(n_4159),
.A2(n_725),
.B(n_724),
.Y(n_4774)
);

AND2x4_ASAP7_75t_L g4775 ( 
.A(n_4458),
.B(n_726),
.Y(n_4775)
);

OAI21x1_ASAP7_75t_SL g4776 ( 
.A1(n_4428),
.A2(n_728),
.B(n_727),
.Y(n_4776)
);

A2O1A1Ixp33_ASAP7_75t_L g4777 ( 
.A1(n_4425),
.A2(n_728),
.B(n_729),
.C(n_727),
.Y(n_4777)
);

INVx3_ASAP7_75t_SL g4778 ( 
.A(n_4269),
.Y(n_4778)
);

INVx3_ASAP7_75t_L g4779 ( 
.A(n_4422),
.Y(n_4779)
);

A2O1A1Ixp33_ASAP7_75t_L g4780 ( 
.A1(n_4420),
.A2(n_729),
.B(n_730),
.C(n_728),
.Y(n_4780)
);

OAI21xp5_ASAP7_75t_L g4781 ( 
.A1(n_4142),
.A2(n_730),
.B(n_729),
.Y(n_4781)
);

AOI21xp5_ASAP7_75t_L g4782 ( 
.A1(n_4245),
.A2(n_731),
.B(n_730),
.Y(n_4782)
);

OAI22xp5_ASAP7_75t_L g4783 ( 
.A1(n_4177),
.A2(n_732),
.B1(n_733),
.B2(n_731),
.Y(n_4783)
);

BUFx10_ASAP7_75t_L g4784 ( 
.A(n_4171),
.Y(n_4784)
);

OAI21xp5_ASAP7_75t_L g4785 ( 
.A1(n_4166),
.A2(n_734),
.B(n_733),
.Y(n_4785)
);

NAND2xp33_ASAP7_75t_R g4786 ( 
.A(n_4396),
.B(n_1119),
.Y(n_4786)
);

AOI211x1_ASAP7_75t_L g4787 ( 
.A1(n_4131),
.A2(n_735),
.B(n_736),
.C(n_734),
.Y(n_4787)
);

OAI21x1_ASAP7_75t_L g4788 ( 
.A1(n_4655),
.A2(n_737),
.B(n_736),
.Y(n_4788)
);

AOI21x1_ASAP7_75t_L g4789 ( 
.A1(n_4486),
.A2(n_737),
.B(n_736),
.Y(n_4789)
);

BUFx6f_ASAP7_75t_L g4790 ( 
.A(n_4277),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4301),
.Y(n_4791)
);

OAI21xp5_ASAP7_75t_L g4792 ( 
.A1(n_4383),
.A2(n_739),
.B(n_738),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_4216),
.B(n_4410),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4390),
.B(n_738),
.Y(n_4794)
);

OAI22xp5_ASAP7_75t_L g4795 ( 
.A1(n_4265),
.A2(n_740),
.B1(n_741),
.B2(n_739),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4312),
.Y(n_4796)
);

INVx6_ASAP7_75t_SL g4797 ( 
.A(n_4412),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4417),
.B(n_741),
.Y(n_4798)
);

OAI22x1_ASAP7_75t_L g4799 ( 
.A1(n_4236),
.A2(n_742),
.B1(n_743),
.B2(n_741),
.Y(n_4799)
);

CKINVDCx16_ASAP7_75t_R g4800 ( 
.A(n_4222),
.Y(n_4800)
);

AOI21xp33_ASAP7_75t_L g4801 ( 
.A1(n_4207),
.A2(n_743),
.B(n_742),
.Y(n_4801)
);

OAI22x1_ASAP7_75t_L g4802 ( 
.A1(n_4327),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4209),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4419),
.B(n_4444),
.Y(n_4804)
);

INVxp67_ASAP7_75t_L g4805 ( 
.A(n_4446),
.Y(n_4805)
);

AO22x2_ASAP7_75t_L g4806 ( 
.A1(n_4160),
.A2(n_745),
.B1(n_746),
.B2(n_744),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_4252),
.A2(n_4304),
.B(n_4186),
.Y(n_4807)
);

OAI21x1_ASAP7_75t_L g4808 ( 
.A1(n_4677),
.A2(n_746),
.B(n_745),
.Y(n_4808)
);

BUFx6f_ASAP7_75t_L g4809 ( 
.A(n_4153),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4616),
.A2(n_747),
.B(n_746),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4212),
.Y(n_4811)
);

AO31x2_ASAP7_75t_L g4812 ( 
.A1(n_4680),
.A2(n_748),
.A3(n_749),
.B(n_747),
.Y(n_4812)
);

OAI21x1_ASAP7_75t_L g4813 ( 
.A1(n_4675),
.A2(n_748),
.B(n_747),
.Y(n_4813)
);

OAI21xp5_ASAP7_75t_L g4814 ( 
.A1(n_4394),
.A2(n_750),
.B(n_749),
.Y(n_4814)
);

AO31x2_ASAP7_75t_L g4815 ( 
.A1(n_4630),
.A2(n_752),
.A3(n_753),
.B(n_751),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_SL g4816 ( 
.A(n_4349),
.B(n_752),
.Y(n_4816)
);

NAND2x1p5_ASAP7_75t_L g4817 ( 
.A(n_4153),
.B(n_753),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4219),
.Y(n_4818)
);

INVx1_ASAP7_75t_SL g4819 ( 
.A(n_4121),
.Y(n_4819)
);

AO21x1_ASAP7_75t_L g4820 ( 
.A1(n_4514),
.A2(n_754),
.B(n_753),
.Y(n_4820)
);

INVxp67_ASAP7_75t_SL g4821 ( 
.A(n_4474),
.Y(n_4821)
);

AND2x4_ASAP7_75t_L g4822 ( 
.A(n_4307),
.B(n_754),
.Y(n_4822)
);

AND2x4_ASAP7_75t_L g4823 ( 
.A(n_4412),
.B(n_755),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4233),
.Y(n_4824)
);

OAI21x1_ASAP7_75t_L g4825 ( 
.A1(n_4227),
.A2(n_757),
.B(n_756),
.Y(n_4825)
);

AOI21xp5_ASAP7_75t_L g4826 ( 
.A1(n_4618),
.A2(n_757),
.B(n_756),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4176),
.A2(n_758),
.B(n_756),
.Y(n_4827)
);

NOR4xp25_ASAP7_75t_L g4828 ( 
.A(n_4155),
.B(n_759),
.C(n_760),
.D(n_758),
.Y(n_4828)
);

A2O1A1Ixp33_ASAP7_75t_L g4829 ( 
.A1(n_4306),
.A2(n_760),
.B(n_761),
.C(n_758),
.Y(n_4829)
);

A2O1A1Ixp33_ASAP7_75t_L g4830 ( 
.A1(n_4593),
.A2(n_761),
.B(n_762),
.C(n_760),
.Y(n_4830)
);

NAND3x1_ASAP7_75t_L g4831 ( 
.A(n_4284),
.B(n_763),
.C(n_762),
.Y(n_4831)
);

OAI21x1_ASAP7_75t_L g4832 ( 
.A1(n_4315),
.A2(n_4681),
.B(n_4195),
.Y(n_4832)
);

BUFx2_ASAP7_75t_L g4833 ( 
.A(n_4495),
.Y(n_4833)
);

O2A1O1Ixp33_ASAP7_75t_SL g4834 ( 
.A1(n_4541),
.A2(n_763),
.B(n_764),
.C(n_762),
.Y(n_4834)
);

AOI21xp5_ASAP7_75t_L g4835 ( 
.A1(n_4667),
.A2(n_764),
.B(n_763),
.Y(n_4835)
);

AOI221xp5_ASAP7_75t_SL g4836 ( 
.A1(n_4466),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_4836)
);

AOI21xp5_ASAP7_75t_L g4837 ( 
.A1(n_4627),
.A2(n_4192),
.B(n_4658),
.Y(n_4837)
);

NOR2xp33_ASAP7_75t_SL g4838 ( 
.A(n_4237),
.B(n_1115),
.Y(n_4838)
);

OAI21x1_ASAP7_75t_L g4839 ( 
.A1(n_4494),
.A2(n_765),
.B(n_764),
.Y(n_4839)
);

BUFx6f_ASAP7_75t_L g4840 ( 
.A(n_4153),
.Y(n_4840)
);

A2O1A1Ixp33_ASAP7_75t_L g4841 ( 
.A1(n_4510),
.A2(n_766),
.B(n_767),
.C(n_765),
.Y(n_4841)
);

OAI21x1_ASAP7_75t_L g4842 ( 
.A1(n_4223),
.A2(n_767),
.B(n_766),
.Y(n_4842)
);

BUFx8_ASAP7_75t_L g4843 ( 
.A(n_4317),
.Y(n_4843)
);

OAI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_4170),
.A2(n_768),
.B(n_766),
.Y(n_4844)
);

AOI21xp5_ASAP7_75t_L g4845 ( 
.A1(n_4612),
.A2(n_769),
.B(n_768),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4273),
.Y(n_4846)
);

BUFx2_ASAP7_75t_L g4847 ( 
.A(n_4518),
.Y(n_4847)
);

AO21x1_ASAP7_75t_L g4848 ( 
.A1(n_4462),
.A2(n_770),
.B(n_769),
.Y(n_4848)
);

OAI21xp5_ASAP7_75t_L g4849 ( 
.A1(n_4568),
.A2(n_771),
.B(n_770),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4452),
.B(n_770),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4505),
.B(n_771),
.Y(n_4851)
);

O2A1O1Ixp33_ASAP7_75t_SL g4852 ( 
.A1(n_4120),
.A2(n_773),
.B(n_774),
.C(n_772),
.Y(n_4852)
);

AO31x2_ASAP7_75t_L g4853 ( 
.A1(n_4638),
.A2(n_773),
.A3(n_774),
.B(n_772),
.Y(n_4853)
);

INVx1_ASAP7_75t_SL g4854 ( 
.A(n_4328),
.Y(n_4854)
);

OAI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_4663),
.A2(n_773),
.B(n_772),
.Y(n_4855)
);

INVx4_ASAP7_75t_L g4856 ( 
.A(n_4163),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4282),
.Y(n_4857)
);

AO31x2_ASAP7_75t_L g4858 ( 
.A1(n_4666),
.A2(n_775),
.A3(n_776),
.B(n_774),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_SL g4859 ( 
.A(n_4516),
.B(n_775),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4283),
.Y(n_4860)
);

INVxp67_ASAP7_75t_SL g4861 ( 
.A(n_4181),
.Y(n_4861)
);

AOI21xp5_ASAP7_75t_SL g4862 ( 
.A1(n_4545),
.A2(n_776),
.B(n_775),
.Y(n_4862)
);

O2A1O1Ixp5_ASAP7_75t_L g4863 ( 
.A1(n_4631),
.A2(n_777),
.B(n_778),
.C(n_776),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4292),
.Y(n_4864)
);

AOI221x1_ASAP7_75t_L g4865 ( 
.A1(n_4325),
.A2(n_779),
.B1(n_780),
.B2(n_778),
.C(n_777),
.Y(n_4865)
);

OAI21x1_ASAP7_75t_L g4866 ( 
.A1(n_4619),
.A2(n_778),
.B(n_777),
.Y(n_4866)
);

BUFx2_ASAP7_75t_L g4867 ( 
.A(n_4163),
.Y(n_4867)
);

AOI21xp5_ASAP7_75t_L g4868 ( 
.A1(n_4183),
.A2(n_4331),
.B(n_4355),
.Y(n_4868)
);

INVx3_ASAP7_75t_SL g4869 ( 
.A(n_4173),
.Y(n_4869)
);

NOR4xp25_ASAP7_75t_L g4870 ( 
.A(n_4179),
.B(n_780),
.C(n_781),
.D(n_779),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4525),
.B(n_780),
.Y(n_4871)
);

OAI22xp5_ASAP7_75t_L g4872 ( 
.A1(n_4625),
.A2(n_782),
.B1(n_783),
.B2(n_781),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4338),
.Y(n_4873)
);

A2O1A1Ixp33_ASAP7_75t_L g4874 ( 
.A1(n_4266),
.A2(n_782),
.B(n_783),
.C(n_781),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4530),
.B(n_783),
.Y(n_4875)
);

AO21x2_ASAP7_75t_L g4876 ( 
.A1(n_4504),
.A2(n_785),
.B(n_784),
.Y(n_4876)
);

AOI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4378),
.A2(n_787),
.B(n_784),
.Y(n_4877)
);

NOR3xp33_ASAP7_75t_L g4878 ( 
.A(n_4174),
.B(n_795),
.C(n_787),
.Y(n_4878)
);

AOI21x1_ASAP7_75t_L g4879 ( 
.A1(n_4124),
.A2(n_787),
.B(n_784),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_L g4880 ( 
.A(n_4132),
.B(n_788),
.Y(n_4880)
);

AOI21xp5_ASAP7_75t_L g4881 ( 
.A1(n_4370),
.A2(n_789),
.B(n_788),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4215),
.Y(n_4882)
);

AOI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_4617),
.A2(n_791),
.B(n_790),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4350),
.Y(n_4884)
);

OAI21x1_ASAP7_75t_L g4885 ( 
.A1(n_4225),
.A2(n_791),
.B(n_790),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4350),
.Y(n_4886)
);

BUFx3_ASAP7_75t_L g4887 ( 
.A(n_4300),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4535),
.B(n_790),
.Y(n_4888)
);

O2A1O1Ixp33_ASAP7_75t_SL g4889 ( 
.A1(n_4280),
.A2(n_793),
.B(n_794),
.C(n_792),
.Y(n_4889)
);

AO31x2_ASAP7_75t_L g4890 ( 
.A1(n_4642),
.A2(n_793),
.A3(n_794),
.B(n_792),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_L g4891 ( 
.A(n_4549),
.B(n_792),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4240),
.Y(n_4892)
);

CKINVDCx5p33_ASAP7_75t_R g4893 ( 
.A(n_4258),
.Y(n_4893)
);

OAI21xp5_ASAP7_75t_L g4894 ( 
.A1(n_4508),
.A2(n_794),
.B(n_793),
.Y(n_4894)
);

OAI21x1_ASAP7_75t_L g4895 ( 
.A1(n_4515),
.A2(n_796),
.B(n_795),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4324),
.Y(n_4896)
);

OAI22xp33_ASAP7_75t_L g4897 ( 
.A1(n_4477),
.A2(n_797),
.B1(n_798),
.B2(n_796),
.Y(n_4897)
);

BUFx8_ASAP7_75t_SL g4898 ( 
.A(n_4286),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4594),
.B(n_797),
.Y(n_4899)
);

INVx2_ASAP7_75t_L g4900 ( 
.A(n_4471),
.Y(n_4900)
);

NAND2x1p5_ASAP7_75t_L g4901 ( 
.A(n_4163),
.B(n_797),
.Y(n_4901)
);

OAI21x1_ASAP7_75t_L g4902 ( 
.A1(n_4543),
.A2(n_799),
.B(n_798),
.Y(n_4902)
);

OR2x2_ASAP7_75t_L g4903 ( 
.A(n_4447),
.B(n_799),
.Y(n_4903)
);

AOI21xp5_ASAP7_75t_L g4904 ( 
.A1(n_4539),
.A2(n_801),
.B(n_800),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4234),
.Y(n_4905)
);

AOI21xp5_ASAP7_75t_L g4906 ( 
.A1(n_4384),
.A2(n_801),
.B(n_800),
.Y(n_4906)
);

OAI21x1_ASAP7_75t_L g4907 ( 
.A1(n_4598),
.A2(n_802),
.B(n_800),
.Y(n_4907)
);

NOR3xp33_ASAP7_75t_L g4908 ( 
.A(n_4557),
.B(n_811),
.C(n_803),
.Y(n_4908)
);

BUFx2_ASAP7_75t_R g4909 ( 
.A(n_4169),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4238),
.Y(n_4910)
);

BUFx2_ASAP7_75t_L g4911 ( 
.A(n_4387),
.Y(n_4911)
);

AOI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4595),
.A2(n_803),
.B(n_802),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4239),
.Y(n_4913)
);

CKINVDCx6p67_ASAP7_75t_R g4914 ( 
.A(n_4335),
.Y(n_4914)
);

OAI21x1_ASAP7_75t_L g4915 ( 
.A1(n_4326),
.A2(n_803),
.B(n_802),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4296),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4261),
.B(n_804),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4498),
.Y(n_4918)
);

CKINVDCx20_ASAP7_75t_R g4919 ( 
.A(n_4270),
.Y(n_4919)
);

INVx3_ASAP7_75t_L g4920 ( 
.A(n_4144),
.Y(n_4920)
);

NAND2x1p5_ASAP7_75t_L g4921 ( 
.A(n_4385),
.B(n_804),
.Y(n_4921)
);

AOI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4620),
.A2(n_805),
.B(n_804),
.Y(n_4922)
);

INVx2_ASAP7_75t_L g4923 ( 
.A(n_4526),
.Y(n_4923)
);

INVx2_ASAP7_75t_SL g4924 ( 
.A(n_4137),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4133),
.B(n_805),
.Y(n_4925)
);

AO31x2_ASAP7_75t_L g4926 ( 
.A1(n_4561),
.A2(n_807),
.A3(n_808),
.B(n_806),
.Y(n_4926)
);

AOI21xp5_ASAP7_75t_L g4927 ( 
.A1(n_4613),
.A2(n_4648),
.B(n_4334),
.Y(n_4927)
);

AOI21xp5_ASAP7_75t_L g4928 ( 
.A1(n_4287),
.A2(n_807),
.B(n_806),
.Y(n_4928)
);

AND2x2_ASAP7_75t_SL g4929 ( 
.A(n_4200),
.B(n_807),
.Y(n_4929)
);

AND2x4_ASAP7_75t_L g4930 ( 
.A(n_4427),
.B(n_808),
.Y(n_4930)
);

AO31x2_ASAP7_75t_L g4931 ( 
.A1(n_4529),
.A2(n_809),
.A3(n_810),
.B(n_808),
.Y(n_4931)
);

OA21x2_ASAP7_75t_L g4932 ( 
.A1(n_4343),
.A2(n_810),
.B(n_809),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4136),
.B(n_4295),
.Y(n_4933)
);

AOI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4127),
.A2(n_1112),
.B1(n_1113),
.B2(n_1107),
.Y(n_4934)
);

AO31x2_ASAP7_75t_L g4935 ( 
.A1(n_4536),
.A2(n_812),
.A3(n_813),
.B(n_810),
.Y(n_4935)
);

OAI21x1_ASAP7_75t_L g4936 ( 
.A1(n_4393),
.A2(n_813),
.B(n_812),
.Y(n_4936)
);

AOI21xp5_ASAP7_75t_L g4937 ( 
.A1(n_4652),
.A2(n_813),
.B(n_812),
.Y(n_4937)
);

OAI21x1_ASAP7_75t_L g4938 ( 
.A1(n_4564),
.A2(n_815),
.B(n_814),
.Y(n_4938)
);

NOR4xp25_ASAP7_75t_L g4939 ( 
.A(n_4254),
.B(n_815),
.C(n_816),
.D(n_814),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4302),
.Y(n_4940)
);

BUFx6f_ASAP7_75t_L g4941 ( 
.A(n_4144),
.Y(n_4941)
);

AO31x2_ASAP7_75t_L g4942 ( 
.A1(n_4538),
.A2(n_815),
.A3(n_816),
.B(n_814),
.Y(n_4942)
);

NOR2xp67_ASAP7_75t_L g4943 ( 
.A(n_4285),
.B(n_817),
.Y(n_4943)
);

CKINVDCx11_ASAP7_75t_R g4944 ( 
.A(n_4213),
.Y(n_4944)
);

A2O1A1Ixp33_ASAP7_75t_L g4945 ( 
.A1(n_4250),
.A2(n_817),
.B(n_818),
.C(n_816),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4311),
.Y(n_4946)
);

BUFx12f_ASAP7_75t_L g4947 ( 
.A(n_4335),
.Y(n_4947)
);

OR2x6_ASAP7_75t_L g4948 ( 
.A(n_4477),
.B(n_817),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4119),
.B(n_818),
.Y(n_4949)
);

INVxp67_ASAP7_75t_SL g4950 ( 
.A(n_4181),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_SL g4951 ( 
.A(n_4459),
.B(n_818),
.Y(n_4951)
);

AO32x2_ASAP7_75t_L g4952 ( 
.A1(n_4151),
.A2(n_821),
.A3(n_822),
.B1(n_820),
.B2(n_819),
.Y(n_4952)
);

INVx5_ASAP7_75t_L g4953 ( 
.A(n_4611),
.Y(n_4953)
);

NOR2xp33_ASAP7_75t_L g4954 ( 
.A(n_4556),
.B(n_819),
.Y(n_4954)
);

NAND3x1_ASAP7_75t_L g4955 ( 
.A(n_4230),
.B(n_4351),
.C(n_4512),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4329),
.Y(n_4956)
);

NOR4xp25_ASAP7_75t_L g4957 ( 
.A(n_4262),
.B(n_820),
.C(n_822),
.D(n_819),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_4562),
.B(n_4609),
.Y(n_4958)
);

OAI21xp5_ASAP7_75t_L g4959 ( 
.A1(n_4389),
.A2(n_824),
.B(n_823),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4552),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4552),
.Y(n_4961)
);

INVx2_ASAP7_75t_SL g4962 ( 
.A(n_4310),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4575),
.Y(n_4963)
);

OAI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_4478),
.A2(n_824),
.B1(n_825),
.B2(n_823),
.Y(n_4964)
);

A2O1A1Ixp33_ASAP7_75t_L g4965 ( 
.A1(n_4255),
.A2(n_825),
.B(n_826),
.C(n_824),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4575),
.Y(n_4966)
);

AOI21xp5_ASAP7_75t_L g4967 ( 
.A1(n_4652),
.A2(n_826),
.B(n_825),
.Y(n_4967)
);

BUFx2_ASAP7_75t_R g4968 ( 
.A(n_4180),
.Y(n_4968)
);

AOI22xp33_ASAP7_75t_L g4969 ( 
.A1(n_4644),
.A2(n_827),
.B1(n_828),
.B2(n_826),
.Y(n_4969)
);

AND2x4_ASAP7_75t_L g4970 ( 
.A(n_4478),
.B(n_827),
.Y(n_4970)
);

NAND2xp33_ASAP7_75t_L g4971 ( 
.A(n_4272),
.B(n_4611),
.Y(n_4971)
);

NAND3x1_ASAP7_75t_L g4972 ( 
.A(n_4248),
.B(n_828),
.C(n_827),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4551),
.B(n_828),
.Y(n_4973)
);

AND2x4_ASAP7_75t_L g4974 ( 
.A(n_4506),
.B(n_829),
.Y(n_4974)
);

AOI21xp5_ASAP7_75t_L g4975 ( 
.A1(n_4249),
.A2(n_830),
.B(n_829),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4199),
.B(n_829),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4205),
.B(n_830),
.Y(n_4977)
);

O2A1O1Ixp33_ASAP7_75t_SL g4978 ( 
.A1(n_4429),
.A2(n_831),
.B(n_832),
.C(n_830),
.Y(n_4978)
);

BUFx3_ASAP7_75t_L g4979 ( 
.A(n_4407),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4263),
.Y(n_4980)
);

O2A1O1Ixp5_ASAP7_75t_L g4981 ( 
.A1(n_4671),
.A2(n_833),
.B(n_834),
.C(n_832),
.Y(n_4981)
);

NOR2x1_ASAP7_75t_SL g4982 ( 
.A(n_4506),
.B(n_832),
.Y(n_4982)
);

BUFx6f_ASAP7_75t_L g4983 ( 
.A(n_4459),
.Y(n_4983)
);

A2O1A1Ixp33_ASAP7_75t_L g4984 ( 
.A1(n_4253),
.A2(n_834),
.B(n_835),
.C(n_833),
.Y(n_4984)
);

NOR2xp33_ASAP7_75t_SL g4985 ( 
.A(n_4368),
.B(n_1100),
.Y(n_4985)
);

AOI221xp5_ASAP7_75t_SL g4986 ( 
.A1(n_4138),
.A2(n_4357),
.B1(n_4476),
.B2(n_4483),
.C(n_4534),
.Y(n_4986)
);

INVx2_ASAP7_75t_SL g4987 ( 
.A(n_4441),
.Y(n_4987)
);

OAI21x1_ASAP7_75t_L g4988 ( 
.A1(n_4558),
.A2(n_835),
.B(n_833),
.Y(n_4988)
);

AO31x2_ASAP7_75t_L g4989 ( 
.A1(n_4563),
.A2(n_836),
.A3(n_837),
.B(n_835),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4210),
.B(n_836),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4214),
.B(n_837),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4299),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4481),
.B(n_837),
.Y(n_4993)
);

AOI221x1_ASAP7_75t_L g4994 ( 
.A1(n_4423),
.A2(n_840),
.B1(n_841),
.B2(n_839),
.C(n_838),
.Y(n_4994)
);

NAND3x1_ASAP7_75t_L g4995 ( 
.A(n_4432),
.B(n_839),
.C(n_838),
.Y(n_4995)
);

OAI21x1_ASAP7_75t_L g4996 ( 
.A1(n_4574),
.A2(n_839),
.B(n_838),
.Y(n_4996)
);

NOR2xp33_ASAP7_75t_SL g4997 ( 
.A(n_4611),
.B(n_1105),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4188),
.B(n_840),
.Y(n_4998)
);

INVx5_ASAP7_75t_L g4999 ( 
.A(n_4272),
.Y(n_4999)
);

BUFx3_ASAP7_75t_L g5000 ( 
.A(n_4460),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_4577),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4388),
.B(n_840),
.Y(n_5002)
);

AO31x2_ASAP7_75t_L g5003 ( 
.A1(n_4583),
.A2(n_842),
.A3(n_843),
.B(n_841),
.Y(n_5003)
);

NOR2x1_ASAP7_75t_SL g5004 ( 
.A(n_4524),
.B(n_841),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4318),
.Y(n_5005)
);

INVx8_ASAP7_75t_L g5006 ( 
.A(n_4484),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4128),
.B(n_842),
.Y(n_5007)
);

OAI21xp5_ASAP7_75t_L g5008 ( 
.A1(n_4439),
.A2(n_4442),
.B(n_4358),
.Y(n_5008)
);

BUFx3_ASAP7_75t_L g5009 ( 
.A(n_4405),
.Y(n_5009)
);

BUFx3_ASAP7_75t_L g5010 ( 
.A(n_4309),
.Y(n_5010)
);

AOI21xp5_ASAP7_75t_L g5011 ( 
.A1(n_4354),
.A2(n_844),
.B(n_842),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4147),
.B(n_844),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4185),
.B(n_844),
.Y(n_5013)
);

AOI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_4584),
.A2(n_846),
.B(n_845),
.Y(n_5014)
);

AOI21xp5_ASAP7_75t_L g5015 ( 
.A1(n_4599),
.A2(n_846),
.B(n_845),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4431),
.Y(n_5016)
);

OAI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_4482),
.A2(n_847),
.B(n_845),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4431),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4414),
.B(n_4606),
.Y(n_5019)
);

AOI221xp5_ASAP7_75t_SL g5020 ( 
.A1(n_4228),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4433),
.Y(n_5021)
);

OAI21x1_ASAP7_75t_L g5022 ( 
.A1(n_4436),
.A2(n_848),
.B(n_847),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4158),
.B(n_848),
.Y(n_5023)
);

AOI21xp5_ASAP7_75t_L g5024 ( 
.A1(n_4117),
.A2(n_849),
.B(n_848),
.Y(n_5024)
);

INVxp67_ASAP7_75t_SL g5025 ( 
.A(n_4181),
.Y(n_5025)
);

OA21x2_ASAP7_75t_L g5026 ( 
.A1(n_4542),
.A2(n_850),
.B(n_849),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4433),
.Y(n_5027)
);

OAI21x1_ASAP7_75t_L g5028 ( 
.A1(n_4548),
.A2(n_851),
.B(n_850),
.Y(n_5028)
);

OAI21x1_ASAP7_75t_L g5029 ( 
.A1(n_4674),
.A2(n_4340),
.B(n_4664),
.Y(n_5029)
);

BUFx3_ASAP7_75t_L g5030 ( 
.A(n_4409),
.Y(n_5030)
);

NAND2xp33_ASAP7_75t_R g5031 ( 
.A(n_4669),
.B(n_1102),
.Y(n_5031)
);

OAI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_4503),
.A2(n_852),
.B(n_851),
.Y(n_5032)
);

AOI21x1_ASAP7_75t_L g5033 ( 
.A1(n_4418),
.A2(n_853),
.B(n_852),
.Y(n_5033)
);

A2O1A1Ixp33_ASAP7_75t_L g5034 ( 
.A1(n_4395),
.A2(n_854),
.B(n_855),
.C(n_853),
.Y(n_5034)
);

INVxp67_ASAP7_75t_L g5035 ( 
.A(n_4129),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4472),
.Y(n_5036)
);

BUFx6f_ASAP7_75t_L g5037 ( 
.A(n_4459),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_4347),
.B(n_853),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4641),
.A2(n_855),
.B(n_854),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4402),
.B(n_856),
.Y(n_5040)
);

OAI21xp5_ASAP7_75t_L g5041 ( 
.A1(n_4547),
.A2(n_857),
.B(n_856),
.Y(n_5041)
);

OAI22xp5_ASAP7_75t_L g5042 ( 
.A1(n_4645),
.A2(n_857),
.B1(n_858),
.B2(n_856),
.Y(n_5042)
);

OAI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4634),
.A2(n_859),
.B(n_858),
.Y(n_5043)
);

OAI22x1_ASAP7_75t_L g5044 ( 
.A1(n_4290),
.A2(n_859),
.B1(n_860),
.B2(n_858),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_4559),
.B(n_860),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_SL g5046 ( 
.A(n_4540),
.B(n_861),
.Y(n_5046)
);

OAI21x1_ASAP7_75t_SL g5047 ( 
.A1(n_4501),
.A2(n_862),
.B(n_861),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_4332),
.B(n_862),
.Y(n_5048)
);

AND3x4_ASAP7_75t_L g5049 ( 
.A(n_4290),
.B(n_863),
.C(n_862),
.Y(n_5049)
);

AOI221x1_ASAP7_75t_L g5050 ( 
.A1(n_4566),
.A2(n_865),
.B1(n_866),
.B2(n_864),
.C(n_863),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_4403),
.Y(n_5051)
);

AND2x4_ASAP7_75t_L g5052 ( 
.A(n_4472),
.B(n_863),
.Y(n_5052)
);

AO22x1_ASAP7_75t_L g5053 ( 
.A1(n_4272),
.A2(n_865),
.B1(n_867),
.B2(n_864),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_SL g5054 ( 
.A1(n_4392),
.A2(n_4520),
.B(n_4607),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4339),
.B(n_864),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4578),
.B(n_865),
.Y(n_5056)
);

OAI21x1_ASAP7_75t_L g5057 ( 
.A1(n_4608),
.A2(n_868),
.B(n_867),
.Y(n_5057)
);

OAI21x1_ASAP7_75t_L g5058 ( 
.A1(n_4592),
.A2(n_869),
.B(n_868),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4585),
.B(n_868),
.Y(n_5059)
);

OAI22xp5_ASAP7_75t_L g5060 ( 
.A1(n_4645),
.A2(n_870),
.B1(n_871),
.B2(n_869),
.Y(n_5060)
);

BUFx12f_ASAP7_75t_L g5061 ( 
.A(n_4409),
.Y(n_5061)
);

OAI21x1_ASAP7_75t_L g5062 ( 
.A1(n_4604),
.A2(n_872),
.B(n_870),
.Y(n_5062)
);

A2O1A1Ixp33_ASAP7_75t_L g5063 ( 
.A1(n_4656),
.A2(n_874),
.B(n_876),
.C(n_873),
.Y(n_5063)
);

OAI22x1_ASAP7_75t_L g5064 ( 
.A1(n_4391),
.A2(n_874),
.B1(n_876),
.B2(n_873),
.Y(n_5064)
);

AOI22xp5_ASAP7_75t_L g5065 ( 
.A1(n_4650),
.A2(n_877),
.B1(n_878),
.B2(n_873),
.Y(n_5065)
);

BUFx2_ASAP7_75t_L g5066 ( 
.A(n_4570),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_4449),
.B(n_877),
.Y(n_5067)
);

AOI21x1_ASAP7_75t_L g5068 ( 
.A1(n_4461),
.A2(n_878),
.B(n_877),
.Y(n_5068)
);

OAI21x1_ASAP7_75t_L g5069 ( 
.A1(n_4509),
.A2(n_879),
.B(n_878),
.Y(n_5069)
);

OAI21xp33_ASAP7_75t_L g5070 ( 
.A1(n_4274),
.A2(n_4455),
.B(n_4356),
.Y(n_5070)
);

INVx4_ASAP7_75t_L g5071 ( 
.A(n_4484),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4600),
.Y(n_5072)
);

NOR3xp33_ASAP7_75t_L g5073 ( 
.A(n_4224),
.B(n_880),
.C(n_879),
.Y(n_5073)
);

INVx5_ASAP7_75t_L g5074 ( 
.A(n_4484),
.Y(n_5074)
);

OAI21xp5_ASAP7_75t_L g5075 ( 
.A1(n_4665),
.A2(n_880),
.B(n_879),
.Y(n_5075)
);

AOI22xp5_ASAP7_75t_L g5076 ( 
.A1(n_4473),
.A2(n_881),
.B1(n_882),
.B2(n_880),
.Y(n_5076)
);

NOR2xp33_ASAP7_75t_L g5077 ( 
.A(n_4221),
.B(n_881),
.Y(n_5077)
);

OAI21x1_ASAP7_75t_L g5078 ( 
.A1(n_4527),
.A2(n_883),
.B(n_882),
.Y(n_5078)
);

OAI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_4576),
.A2(n_884),
.B(n_883),
.Y(n_5079)
);

AOI21xp5_ASAP7_75t_L g5080 ( 
.A1(n_4521),
.A2(n_885),
.B(n_884),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_4403),
.Y(n_5081)
);

OAI21x1_ASAP7_75t_L g5082 ( 
.A1(n_4565),
.A2(n_885),
.B(n_884),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4470),
.B(n_885),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_L g5084 ( 
.A(n_4660),
.B(n_886),
.Y(n_5084)
);

OAI22xp5_ASAP7_75t_L g5085 ( 
.A1(n_4524),
.A2(n_887),
.B1(n_888),
.B2(n_886),
.Y(n_5085)
);

O2A1O1Ixp5_ASAP7_75t_L g5086 ( 
.A1(n_4485),
.A2(n_887),
.B(n_888),
.C(n_886),
.Y(n_5086)
);

AO31x2_ASAP7_75t_L g5087 ( 
.A1(n_4475),
.A2(n_888),
.A3(n_889),
.B(n_887),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4522),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4279),
.B(n_889),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4531),
.Y(n_5090)
);

OAI21x1_ASAP7_75t_L g5091 ( 
.A1(n_4579),
.A2(n_891),
.B(n_890),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_4193),
.Y(n_5092)
);

O2A1O1Ixp5_ASAP7_75t_SL g5093 ( 
.A1(n_4602),
.A2(n_892),
.B(n_893),
.C(n_891),
.Y(n_5093)
);

OAI21x1_ASAP7_75t_L g5094 ( 
.A1(n_4398),
.A2(n_893),
.B(n_892),
.Y(n_5094)
);

NAND3xp33_ASAP7_75t_L g5095 ( 
.A(n_4264),
.B(n_4654),
.C(n_4256),
.Y(n_5095)
);

INVx4_ASAP7_75t_L g5096 ( 
.A(n_4139),
.Y(n_5096)
);

INVx2_ASAP7_75t_L g5097 ( 
.A(n_4193),
.Y(n_5097)
);

OAI21xp5_ASAP7_75t_L g5098 ( 
.A1(n_4640),
.A2(n_894),
.B(n_893),
.Y(n_5098)
);

OA22x2_ASAP7_75t_L g5099 ( 
.A1(n_4533),
.A2(n_895),
.B1(n_896),
.B2(n_894),
.Y(n_5099)
);

O2A1O1Ixp33_ASAP7_75t_SL g5100 ( 
.A1(n_4668),
.A2(n_895),
.B(n_896),
.C(n_894),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4193),
.Y(n_5101)
);

INVx2_ASAP7_75t_L g5102 ( 
.A(n_4251),
.Y(n_5102)
);

OAI21x1_ASAP7_75t_L g5103 ( 
.A1(n_4437),
.A2(n_896),
.B(n_895),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4291),
.B(n_897),
.Y(n_5104)
);

NOR2x1_ASAP7_75t_L g5105 ( 
.A(n_4305),
.B(n_897),
.Y(n_5105)
);

AOI21xp5_ASAP7_75t_L g5106 ( 
.A1(n_4251),
.A2(n_899),
.B(n_898),
.Y(n_5106)
);

OA21x2_ASAP7_75t_L g5107 ( 
.A1(n_4231),
.A2(n_899),
.B(n_898),
.Y(n_5107)
);

OAI21x1_ASAP7_75t_L g5108 ( 
.A1(n_4445),
.A2(n_4448),
.B(n_4626),
.Y(n_5108)
);

AOI21xp5_ASAP7_75t_L g5109 ( 
.A1(n_4251),
.A2(n_900),
.B(n_898),
.Y(n_5109)
);

AOI21xp5_ASAP7_75t_L g5110 ( 
.A1(n_4289),
.A2(n_901),
.B(n_900),
.Y(n_5110)
);

OAI21x1_ASAP7_75t_L g5111 ( 
.A1(n_4635),
.A2(n_902),
.B(n_901),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4544),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4289),
.Y(n_5113)
);

AOI221xp5_ASAP7_75t_L g5114 ( 
.A1(n_4241),
.A2(n_904),
.B1(n_905),
.B2(n_903),
.C(n_902),
.Y(n_5114)
);

O2A1O1Ixp33_ASAP7_75t_L g5115 ( 
.A1(n_4165),
.A2(n_4204),
.B(n_4232),
.C(n_4590),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4289),
.A2(n_903),
.B(n_902),
.Y(n_5116)
);

A2O1A1Ixp33_ASAP7_75t_L g5117 ( 
.A1(n_4421),
.A2(n_905),
.B(n_906),
.C(n_904),
.Y(n_5117)
);

OAI21x1_ASAP7_75t_SL g5118 ( 
.A1(n_4496),
.A2(n_905),
.B(n_904),
.Y(n_5118)
);

OAI21x1_ASAP7_75t_L g5119 ( 
.A1(n_4636),
.A2(n_907),
.B(n_906),
.Y(n_5119)
);

BUFx3_ASAP7_75t_L g5120 ( 
.A(n_4139),
.Y(n_5120)
);

OAI21x1_ASAP7_75t_L g5121 ( 
.A1(n_4366),
.A2(n_909),
.B(n_908),
.Y(n_5121)
);

NOR2xp33_ASAP7_75t_L g5122 ( 
.A(n_4175),
.B(n_910),
.Y(n_5122)
);

AND2x2_ASAP7_75t_L g5123 ( 
.A(n_4629),
.B(n_910),
.Y(n_5123)
);

O2A1O1Ixp5_ASAP7_75t_SL g5124 ( 
.A1(n_4321),
.A2(n_911),
.B(n_912),
.C(n_910),
.Y(n_5124)
);

INVx5_ASAP7_75t_L g5125 ( 
.A(n_4540),
.Y(n_5125)
);

HB1xp67_ASAP7_75t_L g5126 ( 
.A(n_4605),
.Y(n_5126)
);

OAI21x1_ASAP7_75t_L g5127 ( 
.A1(n_4372),
.A2(n_912),
.B(n_911),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_L g5128 ( 
.A(n_4678),
.B(n_912),
.Y(n_5128)
);

AO31x2_ASAP7_75t_L g5129 ( 
.A1(n_4499),
.A2(n_914),
.A3(n_915),
.B(n_913),
.Y(n_5129)
);

AOI21xp5_ASAP7_75t_L g5130 ( 
.A1(n_4314),
.A2(n_914),
.B(n_913),
.Y(n_5130)
);

OAI21x1_ASAP7_75t_L g5131 ( 
.A1(n_4614),
.A2(n_914),
.B(n_913),
.Y(n_5131)
);

OAI21xp5_ASAP7_75t_L g5132 ( 
.A1(n_4643),
.A2(n_916),
.B(n_915),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_SL g5133 ( 
.A(n_4540),
.B(n_916),
.Y(n_5133)
);

A2O1A1Ixp33_ASAP7_75t_L g5134 ( 
.A1(n_4488),
.A2(n_917),
.B(n_918),
.C(n_916),
.Y(n_5134)
);

NOR2xp33_ASAP7_75t_L g5135 ( 
.A(n_4189),
.B(n_917),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_4344),
.B(n_917),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_SL g5137 ( 
.A(n_4622),
.B(n_918),
.Y(n_5137)
);

AND2x4_ASAP7_75t_L g5138 ( 
.A(n_4490),
.B(n_918),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_4330),
.B(n_919),
.Y(n_5139)
);

OAI22xp5_ASAP7_75t_L g5140 ( 
.A1(n_4622),
.A2(n_920),
.B1(n_921),
.B2(n_919),
.Y(n_5140)
);

AND2x2_ASAP7_75t_L g5141 ( 
.A(n_4629),
.B(n_919),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4673),
.Y(n_5142)
);

O2A1O1Ixp5_ASAP7_75t_L g5143 ( 
.A1(n_4657),
.A2(n_921),
.B(n_922),
.C(n_920),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4161),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_4434),
.B(n_4342),
.Y(n_5145)
);

NOR2xp33_ASAP7_75t_L g5146 ( 
.A(n_4218),
.B(n_921),
.Y(n_5146)
);

CKINVDCx11_ASAP7_75t_R g5147 ( 
.A(n_4490),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4314),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_4555),
.B(n_922),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_4359),
.B(n_922),
.Y(n_5150)
);

AOI21x1_ASAP7_75t_SL g5151 ( 
.A1(n_4360),
.A2(n_924),
.B(n_923),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_4361),
.B(n_923),
.Y(n_5152)
);

OAI21x1_ASAP7_75t_L g5153 ( 
.A1(n_4615),
.A2(n_925),
.B(n_924),
.Y(n_5153)
);

CKINVDCx6p67_ASAP7_75t_R g5154 ( 
.A(n_4157),
.Y(n_5154)
);

AO22x2_ASAP7_75t_L g5155 ( 
.A1(n_4589),
.A2(n_925),
.B1(n_926),
.B2(n_924),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_4373),
.B(n_925),
.Y(n_5156)
);

AOI21x1_ASAP7_75t_L g5157 ( 
.A1(n_4789),
.A2(n_4157),
.B(n_4601),
.Y(n_5157)
);

OAI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4761),
.A2(n_4582),
.B(n_4554),
.Y(n_5158)
);

OAI21x1_ASAP7_75t_L g5159 ( 
.A1(n_4699),
.A2(n_4507),
.B(n_4489),
.Y(n_5159)
);

OAI22xp5_ASAP7_75t_L g5160 ( 
.A1(n_5049),
.A2(n_4622),
.B1(n_4497),
.B2(n_4644),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_SL g5161 ( 
.A(n_5074),
.B(n_4517),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_4758),
.Y(n_5162)
);

NOR2xp33_ASAP7_75t_L g5163 ( 
.A(n_4854),
.B(n_4513),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4684),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_4882),
.B(n_4580),
.Y(n_5165)
);

AOI221xp5_ASAP7_75t_L g5166 ( 
.A1(n_4957),
.A2(n_4468),
.B1(n_4348),
.B2(n_4386),
.C(n_4377),
.Y(n_5166)
);

OAI21x1_ASAP7_75t_L g5167 ( 
.A1(n_4832),
.A2(n_4837),
.B(n_4711),
.Y(n_5167)
);

NAND3xp33_ASAP7_75t_L g5168 ( 
.A(n_4762),
.B(n_4610),
.C(n_4217),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4685),
.Y(n_5169)
);

OAI21x1_ASAP7_75t_L g5170 ( 
.A1(n_4689),
.A2(n_4686),
.B(n_4696),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_4971),
.A2(n_4208),
.B(n_4362),
.Y(n_5171)
);

A2O1A1Ixp33_ASAP7_75t_L g5172 ( 
.A1(n_4726),
.A2(n_4244),
.B(n_4260),
.C(n_4243),
.Y(n_5172)
);

AOI22xp33_ASAP7_75t_SL g5173 ( 
.A1(n_5006),
.A2(n_4621),
.B1(n_4603),
.B2(n_4550),
.Y(n_5173)
);

AOI22xp33_ASAP7_75t_SL g5174 ( 
.A1(n_5006),
.A2(n_4646),
.B1(n_4397),
.B2(n_4406),
.Y(n_5174)
);

OAI21x1_ASAP7_75t_L g5175 ( 
.A1(n_4688),
.A2(n_4537),
.B(n_4491),
.Y(n_5175)
);

INVx8_ASAP7_75t_L g5176 ( 
.A(n_4725),
.Y(n_5176)
);

AOI22xp33_ASAP7_75t_L g5177 ( 
.A1(n_4878),
.A2(n_4646),
.B1(n_4672),
.B2(n_4457),
.Y(n_5177)
);

BUFx6f_ASAP7_75t_L g5178 ( 
.A(n_4698),
.Y(n_5178)
);

NAND2x1_ASAP7_75t_L g5179 ( 
.A(n_5071),
.B(n_4314),
.Y(n_5179)
);

AO21x2_ASAP7_75t_L g5180 ( 
.A1(n_4721),
.A2(n_4399),
.B(n_4380),
.Y(n_5180)
);

INVx2_ASAP7_75t_L g5181 ( 
.A(n_4765),
.Y(n_5181)
);

OR2x2_ASAP7_75t_L g5182 ( 
.A(n_4682),
.B(n_4567),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4693),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_4701),
.Y(n_5184)
);

NOR2xp33_ASAP7_75t_L g5185 ( 
.A(n_4914),
.B(n_69),
.Y(n_5185)
);

AO31x2_ASAP7_75t_L g5186 ( 
.A1(n_5050),
.A2(n_4242),
.A3(n_4271),
.B(n_4637),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_4717),
.Y(n_5187)
);

OAI21x1_ASAP7_75t_L g5188 ( 
.A1(n_4690),
.A2(n_4493),
.B(n_4464),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_4900),
.B(n_4571),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4737),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4734),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4754),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_4857),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4764),
.Y(n_5194)
);

AO21x2_ASAP7_75t_L g5195 ( 
.A1(n_4927),
.A2(n_4408),
.B(n_4404),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4791),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_4918),
.B(n_4923),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_4796),
.Y(n_5198)
);

OAI21x1_ASAP7_75t_L g5199 ( 
.A1(n_4788),
.A2(n_4807),
.B(n_4808),
.Y(n_5199)
);

AOI21x1_ASAP7_75t_L g5200 ( 
.A1(n_4757),
.A2(n_4288),
.B(n_4278),
.Y(n_5200)
);

INVx2_ASAP7_75t_L g5201 ( 
.A(n_4860),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_4793),
.B(n_4161),
.Y(n_5202)
);

OAI21x1_ASAP7_75t_SL g5203 ( 
.A1(n_5004),
.A2(n_4313),
.B(n_4587),
.Y(n_5203)
);

OR2x2_ASAP7_75t_L g5204 ( 
.A(n_4980),
.B(n_4443),
.Y(n_5204)
);

OAI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_4908),
.A2(n_4546),
.B(n_4523),
.Y(n_5205)
);

OAI21x1_ASAP7_75t_L g5206 ( 
.A1(n_4724),
.A2(n_4532),
.B(n_4511),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4992),
.Y(n_5207)
);

NAND2x1_ASAP7_75t_L g5208 ( 
.A(n_5096),
.B(n_4362),
.Y(n_5208)
);

OAI21x1_ASAP7_75t_L g5209 ( 
.A1(n_4745),
.A2(n_4659),
.B(n_4647),
.Y(n_5209)
);

A2O1A1Ixp33_ASAP7_75t_L g5210 ( 
.A1(n_4702),
.A2(n_4670),
.B(n_4623),
.C(n_4676),
.Y(n_5210)
);

AND2x4_ASAP7_75t_L g5211 ( 
.A(n_5120),
.B(n_4362),
.Y(n_5211)
);

NAND2xp5_ASAP7_75t_L g5212 ( 
.A(n_5001),
.B(n_4411),
.Y(n_5212)
);

AOI22xp33_ASAP7_75t_L g5213 ( 
.A1(n_4929),
.A2(n_4646),
.B1(n_4430),
.B2(n_4364),
.Y(n_5213)
);

NAND2xp5_ASAP7_75t_L g5214 ( 
.A(n_5142),
.B(n_4413),
.Y(n_5214)
);

NAND3xp33_ASAP7_75t_L g5215 ( 
.A(n_5137),
.B(n_4661),
.C(n_4633),
.Y(n_5215)
);

BUFx2_ASAP7_75t_L g5216 ( 
.A(n_4797),
.Y(n_5216)
);

OA21x2_ASAP7_75t_L g5217 ( 
.A1(n_4868),
.A2(n_4649),
.B(n_4632),
.Y(n_5217)
);

AOI22xp33_ASAP7_75t_L g5218 ( 
.A1(n_4709),
.A2(n_4316),
.B1(n_4322),
.B2(n_4456),
.Y(n_5218)
);

BUFx6f_ASAP7_75t_L g5219 ( 
.A(n_4698),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_L g5220 ( 
.A(n_5005),
.B(n_4451),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_4740),
.Y(n_5221)
);

INVx1_ASAP7_75t_SL g5222 ( 
.A(n_5147),
.Y(n_5222)
);

NAND2xp5_ASAP7_75t_L g5223 ( 
.A(n_4892),
.B(n_4492),
.Y(n_5223)
);

OAI21xp5_ASAP7_75t_L g5224 ( 
.A1(n_5143),
.A2(n_4553),
.B(n_4519),
.Y(n_5224)
);

NAND2x1p5_ASAP7_75t_L g5225 ( 
.A(n_4725),
.B(n_4371),
.Y(n_5225)
);

OAI21x1_ASAP7_75t_L g5226 ( 
.A1(n_4746),
.A2(n_4639),
.B(n_4662),
.Y(n_5226)
);

NOR2xp33_ASAP7_75t_L g5227 ( 
.A(n_4838),
.B(n_71),
.Y(n_5227)
);

AND2x2_ASAP7_75t_L g5228 ( 
.A(n_4750),
.B(n_4161),
.Y(n_5228)
);

OR2x6_ASAP7_75t_L g5229 ( 
.A(n_4948),
.B(n_4371),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_SL g5230 ( 
.A(n_5074),
.B(n_4371),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4958),
.B(n_4624),
.Y(n_5231)
);

OAI21x1_ASAP7_75t_L g5232 ( 
.A1(n_4813),
.A2(n_4469),
.B(n_4502),
.Y(n_5232)
);

OAI22xp33_ASAP7_75t_L g5233 ( 
.A1(n_4997),
.A2(n_4628),
.B1(n_4517),
.B2(n_4573),
.Y(n_5233)
);

AOI21xp5_ASAP7_75t_L g5234 ( 
.A1(n_5115),
.A2(n_4517),
.B(n_4374),
.Y(n_5234)
);

AOI22xp33_ASAP7_75t_L g5235 ( 
.A1(n_4948),
.A2(n_4573),
.B1(n_4374),
.B2(n_4450),
.Y(n_5235)
);

INVxp67_ASAP7_75t_L g5236 ( 
.A(n_5000),
.Y(n_5236)
);

OAI21x1_ASAP7_75t_L g5237 ( 
.A1(n_5029),
.A2(n_4573),
.B(n_4374),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_4864),
.Y(n_5238)
);

AO21x2_ASAP7_75t_L g5239 ( 
.A1(n_4828),
.A2(n_4586),
.B(n_4454),
.Y(n_5239)
);

OAI21x1_ASAP7_75t_L g5240 ( 
.A1(n_4774),
.A2(n_4586),
.B(n_4454),
.Y(n_5240)
);

AND2x4_ASAP7_75t_L g5241 ( 
.A(n_4887),
.B(n_926),
.Y(n_5241)
);

HB1xp67_ASAP7_75t_L g5242 ( 
.A(n_4805),
.Y(n_5242)
);

INVxp67_ASAP7_75t_L g5243 ( 
.A(n_4979),
.Y(n_5243)
);

OAI221xp5_ASAP7_75t_SL g5244 ( 
.A1(n_4723),
.A2(n_4450),
.B1(n_928),
.B2(n_929),
.C(n_927),
.Y(n_5244)
);

A2O1A1Ixp33_ASAP7_75t_L g5245 ( 
.A1(n_4943),
.A2(n_4729),
.B(n_4844),
.C(n_4823),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_4803),
.Y(n_5246)
);

AO31x2_ASAP7_75t_L g5247 ( 
.A1(n_5144),
.A2(n_927),
.A3(n_928),
.B(n_926),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_4708),
.Y(n_5248)
);

AOI222xp33_ASAP7_75t_L g5249 ( 
.A1(n_4799),
.A2(n_930),
.B1(n_928),
.B2(n_931),
.C1(n_929),
.C2(n_927),
.Y(n_5249)
);

INVx2_ASAP7_75t_L g5250 ( 
.A(n_4713),
.Y(n_5250)
);

NOR2xp33_ASAP7_75t_L g5251 ( 
.A(n_4947),
.B(n_71),
.Y(n_5251)
);

AOI21xp33_ASAP7_75t_SL g5252 ( 
.A1(n_4760),
.A2(n_931),
.B(n_930),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_4811),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4818),
.Y(n_5254)
);

OAI22xp5_ASAP7_75t_SL g5255 ( 
.A1(n_4919),
.A2(n_932),
.B1(n_933),
.B2(n_930),
.Y(n_5255)
);

OA21x2_ASAP7_75t_L g5256 ( 
.A1(n_4720),
.A2(n_934),
.B(n_932),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_4730),
.Y(n_5257)
);

OAI21x1_ASAP7_75t_L g5258 ( 
.A1(n_4744),
.A2(n_5151),
.B(n_4735),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_SL g5259 ( 
.A(n_5074),
.B(n_934),
.Y(n_5259)
);

BUFx2_ASAP7_75t_L g5260 ( 
.A(n_4797),
.Y(n_5260)
);

CKINVDCx5p33_ASAP7_75t_R g5261 ( 
.A(n_4898),
.Y(n_5261)
);

OA21x2_ASAP7_75t_L g5262 ( 
.A1(n_4781),
.A2(n_935),
.B(n_934),
.Y(n_5262)
);

AOI22xp5_ASAP7_75t_L g5263 ( 
.A1(n_5031),
.A2(n_936),
.B1(n_937),
.B2(n_935),
.Y(n_5263)
);

BUFx3_ASAP7_75t_L g5264 ( 
.A(n_4692),
.Y(n_5264)
);

OAI21x1_ASAP7_75t_L g5265 ( 
.A1(n_4839),
.A2(n_936),
.B(n_935),
.Y(n_5265)
);

INVx2_ASAP7_75t_L g5266 ( 
.A(n_4824),
.Y(n_5266)
);

OAI21x1_ASAP7_75t_L g5267 ( 
.A1(n_5022),
.A2(n_937),
.B(n_936),
.Y(n_5267)
);

AOI21xp5_ASAP7_75t_L g5268 ( 
.A1(n_4999),
.A2(n_938),
.B(n_937),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_4846),
.Y(n_5269)
);

BUFx12f_ASAP7_75t_L g5270 ( 
.A(n_4843),
.Y(n_5270)
);

OAI21x1_ASAP7_75t_L g5271 ( 
.A1(n_4825),
.A2(n_939),
.B(n_938),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_4873),
.Y(n_5272)
);

OAI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_4955),
.A2(n_940),
.B(n_939),
.Y(n_5273)
);

OAI21x1_ASAP7_75t_L g5274 ( 
.A1(n_4727),
.A2(n_941),
.B(n_940),
.Y(n_5274)
);

INVx2_ASAP7_75t_SL g5275 ( 
.A(n_4725),
.Y(n_5275)
);

OAI21x1_ASAP7_75t_L g5276 ( 
.A1(n_4895),
.A2(n_941),
.B(n_940),
.Y(n_5276)
);

A2O1A1Ixp33_ASAP7_75t_L g5277 ( 
.A1(n_5073),
.A2(n_943),
.B(n_944),
.C(n_942),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_4719),
.Y(n_5278)
);

OR2x6_ASAP7_75t_L g5279 ( 
.A(n_4911),
.B(n_942),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4804),
.Y(n_5280)
);

HB1xp67_ASAP7_75t_L g5281 ( 
.A(n_5126),
.Y(n_5281)
);

NOR2xp33_ASAP7_75t_L g5282 ( 
.A(n_5009),
.B(n_71),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4771),
.Y(n_5283)
);

OR2x2_ASAP7_75t_L g5284 ( 
.A(n_4933),
.B(n_942),
.Y(n_5284)
);

AOI21x1_ASAP7_75t_L g5285 ( 
.A1(n_4743),
.A2(n_944),
.B(n_943),
.Y(n_5285)
);

OA21x2_ASAP7_75t_L g5286 ( 
.A1(n_4703),
.A2(n_944),
.B(n_943),
.Y(n_5286)
);

NAND2x1_ASAP7_75t_L g5287 ( 
.A(n_4847),
.B(n_945),
.Y(n_5287)
);

NOR2xp33_ASAP7_75t_L g5288 ( 
.A(n_4985),
.B(n_71),
.Y(n_5288)
);

AOI22xp5_ASAP7_75t_L g5289 ( 
.A1(n_4786),
.A2(n_946),
.B1(n_947),
.B2(n_945),
.Y(n_5289)
);

OA21x2_ASAP7_75t_L g5290 ( 
.A1(n_4710),
.A2(n_946),
.B(n_945),
.Y(n_5290)
);

NOR2xp33_ASAP7_75t_L g5291 ( 
.A(n_5035),
.B(n_72),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4715),
.Y(n_5292)
);

OA21x2_ASAP7_75t_L g5293 ( 
.A1(n_4866),
.A2(n_949),
.B(n_947),
.Y(n_5293)
);

AO21x1_ASAP7_75t_L g5294 ( 
.A1(n_4970),
.A2(n_949),
.B(n_947),
.Y(n_5294)
);

INVx2_ASAP7_75t_L g5295 ( 
.A(n_5092),
.Y(n_5295)
);

OAI22xp5_ASAP7_75t_L g5296 ( 
.A1(n_4999),
.A2(n_950),
.B1(n_952),
.B2(n_949),
.Y(n_5296)
);

OAI21x1_ASAP7_75t_L g5297 ( 
.A1(n_4902),
.A2(n_953),
.B(n_950),
.Y(n_5297)
);

BUFx5_ASAP7_75t_L g5298 ( 
.A(n_5016),
.Y(n_5298)
);

OA21x2_ASAP7_75t_L g5299 ( 
.A1(n_4894),
.A2(n_954),
.B(n_950),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_4728),
.Y(n_5300)
);

A2O1A1Ixp33_ASAP7_75t_L g5301 ( 
.A1(n_4780),
.A2(n_955),
.B(n_956),
.C(n_954),
.Y(n_5301)
);

OA21x2_ASAP7_75t_L g5302 ( 
.A1(n_4700),
.A2(n_955),
.B(n_954),
.Y(n_5302)
);

OAI21x1_ASAP7_75t_L g5303 ( 
.A1(n_4842),
.A2(n_957),
.B(n_956),
.Y(n_5303)
);

AOI22xp33_ASAP7_75t_L g5304 ( 
.A1(n_5070),
.A2(n_5095),
.B1(n_5099),
.B2(n_4974),
.Y(n_5304)
);

BUFx2_ASAP7_75t_L g5305 ( 
.A(n_4867),
.Y(n_5305)
);

OAI21x1_ASAP7_75t_L g5306 ( 
.A1(n_5108),
.A2(n_957),
.B(n_956),
.Y(n_5306)
);

AOI22xp33_ASAP7_75t_L g5307 ( 
.A1(n_4806),
.A2(n_959),
.B1(n_960),
.B2(n_958),
.Y(n_5307)
);

AND2x4_ASAP7_75t_L g5308 ( 
.A(n_4999),
.B(n_958),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_4749),
.Y(n_5309)
);

OAI21x1_ASAP7_75t_L g5310 ( 
.A1(n_5097),
.A2(n_960),
.B(n_959),
.Y(n_5310)
);

OAI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_4981),
.A2(n_962),
.B(n_961),
.Y(n_5311)
);

CKINVDCx11_ASAP7_75t_R g5312 ( 
.A(n_4778),
.Y(n_5312)
);

CKINVDCx6p67_ASAP7_75t_R g5313 ( 
.A(n_5061),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_5101),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5090),
.B(n_1120),
.Y(n_5315)
);

OAI21x1_ASAP7_75t_L g5316 ( 
.A1(n_5102),
.A2(n_963),
.B(n_962),
.Y(n_5316)
);

INVx1_ASAP7_75t_SL g5317 ( 
.A(n_4687),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_5112),
.Y(n_5318)
);

OAI21x1_ASAP7_75t_L g5319 ( 
.A1(n_5113),
.A2(n_963),
.B(n_962),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_5088),
.Y(n_5320)
);

OR2x2_ASAP7_75t_L g5321 ( 
.A(n_4987),
.B(n_4718),
.Y(n_5321)
);

OAI21x1_ASAP7_75t_L g5322 ( 
.A1(n_5148),
.A2(n_964),
.B(n_963),
.Y(n_5322)
);

NOR2x1_ASAP7_75t_R g5323 ( 
.A(n_5030),
.B(n_964),
.Y(n_5323)
);

NAND3xp33_ASAP7_75t_L g5324 ( 
.A(n_4880),
.B(n_965),
.C(n_964),
.Y(n_5324)
);

OA21x2_ASAP7_75t_L g5325 ( 
.A1(n_4865),
.A2(n_966),
.B(n_965),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_4905),
.B(n_966),
.Y(n_5326)
);

OAI21x1_ASAP7_75t_L g5327 ( 
.A1(n_4988),
.A2(n_968),
.B(n_967),
.Y(n_5327)
);

OAI21x1_ASAP7_75t_L g5328 ( 
.A1(n_4996),
.A2(n_969),
.B(n_968),
.Y(n_5328)
);

OAI21x1_ASAP7_75t_L g5329 ( 
.A1(n_4885),
.A2(n_970),
.B(n_969),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_4903),
.Y(n_5330)
);

AO21x2_ASAP7_75t_L g5331 ( 
.A1(n_4870),
.A2(n_971),
.B(n_969),
.Y(n_5331)
);

BUFx2_ASAP7_75t_L g5332 ( 
.A(n_5154),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_5051),
.Y(n_5333)
);

OAI21x1_ASAP7_75t_L g5334 ( 
.A1(n_4936),
.A2(n_972),
.B(n_971),
.Y(n_5334)
);

OAI21x1_ASAP7_75t_L g5335 ( 
.A1(n_4938),
.A2(n_972),
.B(n_971),
.Y(n_5335)
);

OA21x2_ASAP7_75t_L g5336 ( 
.A1(n_4707),
.A2(n_973),
.B(n_972),
.Y(n_5336)
);

AOI21xp33_ASAP7_75t_SL g5337 ( 
.A1(n_4869),
.A2(n_974),
.B(n_973),
.Y(n_5337)
);

INVx3_ASAP7_75t_L g5338 ( 
.A(n_4790),
.Y(n_5338)
);

BUFx3_ASAP7_75t_L g5339 ( 
.A(n_4779),
.Y(n_5339)
);

HB1xp67_ASAP7_75t_L g5340 ( 
.A(n_4821),
.Y(n_5340)
);

AO31x2_ASAP7_75t_L g5341 ( 
.A1(n_4820),
.A2(n_1113),
.A3(n_974),
.B(n_975),
.Y(n_5341)
);

OAI21x1_ASAP7_75t_L g5342 ( 
.A1(n_4733),
.A2(n_975),
.B(n_973),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4736),
.Y(n_5343)
);

OAI21xp5_ASAP7_75t_L g5344 ( 
.A1(n_5086),
.A2(n_976),
.B(n_975),
.Y(n_5344)
);

AND2x4_ASAP7_75t_L g5345 ( 
.A(n_4953),
.B(n_977),
.Y(n_5345)
);

AOI22xp33_ASAP7_75t_L g5346 ( 
.A1(n_4806),
.A2(n_978),
.B1(n_979),
.B2(n_977),
.Y(n_5346)
);

OAI21x1_ASAP7_75t_L g5347 ( 
.A1(n_5121),
.A2(n_980),
.B(n_979),
.Y(n_5347)
);

NOR2xp33_ASAP7_75t_L g5348 ( 
.A(n_4968),
.B(n_72),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4884),
.Y(n_5349)
);

OAI21x1_ASAP7_75t_L g5350 ( 
.A1(n_5127),
.A2(n_980),
.B(n_979),
.Y(n_5350)
);

O2A1O1Ixp33_ASAP7_75t_SL g5351 ( 
.A1(n_4859),
.A2(n_982),
.B(n_983),
.C(n_981),
.Y(n_5351)
);

O2A1O1Ixp33_ASAP7_75t_L g5352 ( 
.A1(n_4795),
.A2(n_982),
.B(n_983),
.C(n_981),
.Y(n_5352)
);

AOI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_4986),
.A2(n_982),
.B1(n_984),
.B2(n_981),
.Y(n_5353)
);

NAND3xp33_ASAP7_75t_L g5354 ( 
.A(n_4787),
.B(n_985),
.C(n_984),
.Y(n_5354)
);

AND2x2_ASAP7_75t_L g5355 ( 
.A(n_4917),
.B(n_72),
.Y(n_5355)
);

OR2x2_ASAP7_75t_L g5356 ( 
.A(n_5010),
.B(n_1104),
.Y(n_5356)
);

INVx4_ASAP7_75t_L g5357 ( 
.A(n_4790),
.Y(n_5357)
);

OAI22xp33_ASAP7_75t_L g5358 ( 
.A1(n_4953),
.A2(n_985),
.B1(n_986),
.B2(n_984),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_4910),
.B(n_1103),
.Y(n_5359)
);

NAND3xp33_ASAP7_75t_L g5360 ( 
.A(n_4768),
.B(n_986),
.C(n_985),
.Y(n_5360)
);

NAND2xp5_ASAP7_75t_L g5361 ( 
.A(n_4913),
.B(n_4916),
.Y(n_5361)
);

OAI21x1_ASAP7_75t_L g5362 ( 
.A1(n_5033),
.A2(n_987),
.B(n_986),
.Y(n_5362)
);

INVx2_ASAP7_75t_SL g5363 ( 
.A(n_4739),
.Y(n_5363)
);

CKINVDCx11_ASAP7_75t_R g5364 ( 
.A(n_4784),
.Y(n_5364)
);

INVx2_ASAP7_75t_L g5365 ( 
.A(n_5081),
.Y(n_5365)
);

OAI21x1_ASAP7_75t_L g5366 ( 
.A1(n_5068),
.A2(n_988),
.B(n_987),
.Y(n_5366)
);

INVx2_ASAP7_75t_L g5367 ( 
.A(n_4704),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_4886),
.Y(n_5368)
);

AOI22xp33_ASAP7_75t_SL g5369 ( 
.A1(n_4982),
.A2(n_988),
.B1(n_989),
.B2(n_987),
.Y(n_5369)
);

AOI211xp5_ASAP7_75t_L g5370 ( 
.A1(n_4748),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_5370)
);

OA21x2_ASAP7_75t_L g5371 ( 
.A1(n_4785),
.A2(n_989),
.B(n_988),
.Y(n_5371)
);

AOI22xp33_ASAP7_75t_L g5372 ( 
.A1(n_4848),
.A2(n_990),
.B1(n_991),
.B2(n_989),
.Y(n_5372)
);

AOI21xp5_ASAP7_75t_L g5373 ( 
.A1(n_4953),
.A2(n_992),
.B(n_990),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5018),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_5021),
.Y(n_5375)
);

AOI21x1_ASAP7_75t_L g5376 ( 
.A1(n_5053),
.A2(n_994),
.B(n_993),
.Y(n_5376)
);

BUFx6f_ASAP7_75t_L g5377 ( 
.A(n_4983),
.Y(n_5377)
);

AND2x2_ASAP7_75t_L g5378 ( 
.A(n_5002),
.B(n_73),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5027),
.Y(n_5379)
);

BUFx12f_ASAP7_75t_L g5380 ( 
.A(n_4944),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_4704),
.Y(n_5381)
);

HB1xp67_ASAP7_75t_L g5382 ( 
.A(n_5036),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_4896),
.Y(n_5383)
);

AND2x2_ASAP7_75t_L g5384 ( 
.A(n_5023),
.B(n_73),
.Y(n_5384)
);

NAND3xp33_ASAP7_75t_L g5385 ( 
.A(n_4836),
.B(n_995),
.C(n_994),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_4940),
.B(n_994),
.Y(n_5386)
);

NOR2xp33_ASAP7_75t_L g5387 ( 
.A(n_4800),
.B(n_74),
.Y(n_5387)
);

OAI21xp5_ASAP7_75t_L g5388 ( 
.A1(n_4830),
.A2(n_997),
.B(n_996),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_4956),
.Y(n_5389)
);

BUFx6f_ASAP7_75t_L g5390 ( 
.A(n_4983),
.Y(n_5390)
);

CKINVDCx6p67_ASAP7_75t_R g5391 ( 
.A(n_4833),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_4731),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_4946),
.Y(n_5393)
);

AOI22xp33_ASAP7_75t_L g5394 ( 
.A1(n_5155),
.A2(n_997),
.B1(n_998),
.B2(n_996),
.Y(n_5394)
);

OAI21x1_ASAP7_75t_L g5395 ( 
.A1(n_4907),
.A2(n_998),
.B(n_997),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4960),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_4961),
.Y(n_5397)
);

OAI22xp5_ASAP7_75t_L g5398 ( 
.A1(n_4934),
.A2(n_1000),
.B1(n_1001),
.B2(n_999),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_4963),
.Y(n_5399)
);

INVxp67_ASAP7_75t_SL g5400 ( 
.A(n_4861),
.Y(n_5400)
);

INVx2_ASAP7_75t_SL g5401 ( 
.A(n_5066),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_4716),
.Y(n_5402)
);

OAI21x1_ASAP7_75t_L g5403 ( 
.A1(n_4950),
.A2(n_1000),
.B(n_999),
.Y(n_5403)
);

OAI21x1_ASAP7_75t_L g5404 ( 
.A1(n_5025),
.A2(n_4879),
.B(n_5028),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_4716),
.Y(n_5405)
);

AOI21xp33_ASAP7_75t_L g5406 ( 
.A1(n_5054),
.A2(n_4752),
.B(n_5020),
.Y(n_5406)
);

INVx1_ASAP7_75t_L g5407 ( 
.A(n_4966),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_4893),
.Y(n_5408)
);

BUFx6f_ASAP7_75t_L g5409 ( 
.A(n_5037),
.Y(n_5409)
);

AO31x2_ASAP7_75t_L g5410 ( 
.A1(n_4994),
.A2(n_1102),
.A3(n_1001),
.B(n_1002),
.Y(n_5410)
);

AO21x2_ASAP7_75t_L g5411 ( 
.A1(n_4776),
.A2(n_1001),
.B(n_999),
.Y(n_5411)
);

OR2x2_ASAP7_75t_L g5412 ( 
.A(n_5019),
.B(n_1102),
.Y(n_5412)
);

AND2x2_ASAP7_75t_L g5413 ( 
.A(n_5123),
.B(n_5141),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_SL g5414 ( 
.A(n_5125),
.B(n_1002),
.Y(n_5414)
);

OAI21xp5_ASAP7_75t_L g5415 ( 
.A1(n_4883),
.A2(n_1003),
.B(n_1002),
.Y(n_5415)
);

OAI21x1_ASAP7_75t_L g5416 ( 
.A1(n_5131),
.A2(n_1004),
.B(n_1003),
.Y(n_5416)
);

OAI21xp5_ASAP7_75t_L g5417 ( 
.A1(n_4841),
.A2(n_1004),
.B(n_1003),
.Y(n_5417)
);

AO21x1_ASAP7_75t_L g5418 ( 
.A1(n_4897),
.A2(n_1005),
.B(n_1004),
.Y(n_5418)
);

OAI22xp33_ASAP7_75t_L g5419 ( 
.A1(n_5044),
.A2(n_1006),
.B1(n_1007),
.B2(n_1005),
.Y(n_5419)
);

A2O1A1Ixp33_ASAP7_75t_L g5420 ( 
.A1(n_4738),
.A2(n_1007),
.B(n_1008),
.C(n_1006),
.Y(n_5420)
);

OAI21x1_ASAP7_75t_L g5421 ( 
.A1(n_5153),
.A2(n_1007),
.B(n_1006),
.Y(n_5421)
);

OAI21x1_ASAP7_75t_L g5422 ( 
.A1(n_5107),
.A2(n_1009),
.B(n_1008),
.Y(n_5422)
);

INVxp67_ASAP7_75t_SL g5423 ( 
.A(n_5105),
.Y(n_5423)
);

AND2x4_ASAP7_75t_L g5424 ( 
.A(n_4856),
.B(n_1009),
.Y(n_5424)
);

NOR2xp67_ASAP7_75t_SL g5425 ( 
.A(n_5125),
.B(n_1010),
.Y(n_5425)
);

NOR2x1_ASAP7_75t_R g5426 ( 
.A(n_5125),
.B(n_1010),
.Y(n_5426)
);

AO32x2_ASAP7_75t_L g5427 ( 
.A1(n_5085),
.A2(n_1012),
.A3(n_1013),
.B1(n_1011),
.B2(n_1010),
.Y(n_5427)
);

OAI21x1_ASAP7_75t_SL g5428 ( 
.A1(n_5118),
.A2(n_1012),
.B(n_1011),
.Y(n_5428)
);

AND2x4_ASAP7_75t_L g5429 ( 
.A(n_4809),
.B(n_1013),
.Y(n_5429)
);

AO31x2_ASAP7_75t_L g5430 ( 
.A1(n_4984),
.A2(n_1015),
.A3(n_1016),
.B(n_1014),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_4931),
.Y(n_5431)
);

INVx3_ASAP7_75t_SL g5432 ( 
.A(n_4819),
.Y(n_5432)
);

AO21x2_ASAP7_75t_L g5433 ( 
.A1(n_4801),
.A2(n_1015),
.B(n_1014),
.Y(n_5433)
);

AOI22xp33_ASAP7_75t_L g5434 ( 
.A1(n_5155),
.A2(n_1016),
.B1(n_1017),
.B2(n_1014),
.Y(n_5434)
);

AOI21xp5_ASAP7_75t_L g5435 ( 
.A1(n_4732),
.A2(n_1017),
.B(n_1016),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_4931),
.Y(n_5436)
);

OAI21x1_ASAP7_75t_L g5437 ( 
.A1(n_5107),
.A2(n_1018),
.B(n_1017),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_4809),
.Y(n_5438)
);

BUFx6f_ASAP7_75t_L g5439 ( 
.A(n_5037),
.Y(n_5439)
);

AND2x4_ASAP7_75t_L g5440 ( 
.A(n_4840),
.B(n_1018),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_4935),
.Y(n_5441)
);

CKINVDCx20_ASAP7_75t_R g5442 ( 
.A(n_4756),
.Y(n_5442)
);

AND2x2_ASAP7_75t_L g5443 ( 
.A(n_5072),
.B(n_74),
.Y(n_5443)
);

AOI221xp5_ASAP7_75t_L g5444 ( 
.A1(n_4722),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.C(n_78),
.Y(n_5444)
);

A2O1A1Ixp33_ASAP7_75t_L g5445 ( 
.A1(n_4792),
.A2(n_1020),
.B(n_1021),
.C(n_1019),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_L g5446 ( 
.A(n_5145),
.B(n_1101),
.Y(n_5446)
);

AOI222xp33_ASAP7_75t_L g5447 ( 
.A1(n_4802),
.A2(n_1023),
.B1(n_1021),
.B2(n_1024),
.C1(n_1022),
.C2(n_1020),
.Y(n_5447)
);

OAI22xp5_ASAP7_75t_L g5448 ( 
.A1(n_4831),
.A2(n_1021),
.B1(n_1022),
.B2(n_1020),
.Y(n_5448)
);

AOI21xp5_ASAP7_75t_L g5449 ( 
.A1(n_5100),
.A2(n_1025),
.B(n_1024),
.Y(n_5449)
);

INVx2_ASAP7_75t_L g5450 ( 
.A(n_4840),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_4706),
.B(n_4949),
.Y(n_5451)
);

OAI21xp5_ASAP7_75t_L g5452 ( 
.A1(n_4939),
.A2(n_1026),
.B(n_1025),
.Y(n_5452)
);

INVx2_ASAP7_75t_L g5453 ( 
.A(n_4935),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_4942),
.Y(n_5454)
);

OAI21x1_ASAP7_75t_L g5455 ( 
.A1(n_5069),
.A2(n_1027),
.B(n_1026),
.Y(n_5455)
);

OAI21x1_ASAP7_75t_L g5456 ( 
.A1(n_5078),
.A2(n_1027),
.B(n_1026),
.Y(n_5456)
);

INVx2_ASAP7_75t_SL g5457 ( 
.A(n_4941),
.Y(n_5457)
);

OAI21x1_ASAP7_75t_L g5458 ( 
.A1(n_5082),
.A2(n_1029),
.B(n_1028),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5052),
.B(n_75),
.Y(n_5459)
);

INVx6_ASAP7_75t_SL g5460 ( 
.A(n_4930),
.Y(n_5460)
);

OAI21x1_ASAP7_75t_L g5461 ( 
.A1(n_5091),
.A2(n_1030),
.B(n_1028),
.Y(n_5461)
);

AO21x2_ASAP7_75t_L g5462 ( 
.A1(n_4855),
.A2(n_1031),
.B(n_1030),
.Y(n_5462)
);

BUFx6f_ASAP7_75t_L g5463 ( 
.A(n_4941),
.Y(n_5463)
);

INVx1_ASAP7_75t_SL g5464 ( 
.A(n_4909),
.Y(n_5464)
);

INVx2_ASAP7_75t_SL g5465 ( 
.A(n_4924),
.Y(n_5465)
);

AOI21xp5_ASAP7_75t_L g5466 ( 
.A1(n_4834),
.A2(n_1031),
.B(n_1030),
.Y(n_5466)
);

OAI21xp5_ASAP7_75t_L g5467 ( 
.A1(n_4705),
.A2(n_1032),
.B(n_1031),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_4942),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_4989),
.Y(n_5469)
);

AOI22xp33_ASAP7_75t_L g5470 ( 
.A1(n_4954),
.A2(n_1034),
.B1(n_1035),
.B2(n_1033),
.Y(n_5470)
);

OAI22xp33_ASAP7_75t_L g5471 ( 
.A1(n_5042),
.A2(n_1034),
.B1(n_1035),
.B2(n_1033),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_5202),
.B(n_5012),
.Y(n_5472)
);

OAI21xp5_ASAP7_75t_L g5473 ( 
.A1(n_5245),
.A2(n_4972),
.B(n_5273),
.Y(n_5473)
);

NAND2xp5_ASAP7_75t_L g5474 ( 
.A(n_5228),
.B(n_4973),
.Y(n_5474)
);

INVx1_ASAP7_75t_SL g5475 ( 
.A(n_5317),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5292),
.B(n_4691),
.Y(n_5476)
);

INVx3_ASAP7_75t_SL g5477 ( 
.A(n_5391),
.Y(n_5477)
);

OAI21x1_ASAP7_75t_L g5478 ( 
.A1(n_5167),
.A2(n_4901),
.B(n_4817),
.Y(n_5478)
);

NAND2xp5_ASAP7_75t_L g5479 ( 
.A(n_5278),
.B(n_5038),
.Y(n_5479)
);

OAI21x1_ASAP7_75t_L g5480 ( 
.A1(n_5237),
.A2(n_4770),
.B(n_5093),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5164),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_5309),
.B(n_5146),
.Y(n_5482)
);

OAI21x1_ASAP7_75t_L g5483 ( 
.A1(n_5170),
.A2(n_4683),
.B(n_5124),
.Y(n_5483)
);

OAI21x1_ASAP7_75t_L g5484 ( 
.A1(n_5199),
.A2(n_4967),
.B(n_4937),
.Y(n_5484)
);

INVx2_ASAP7_75t_L g5485 ( 
.A(n_5340),
.Y(n_5485)
);

AOI21xp5_ASAP7_75t_L g5486 ( 
.A1(n_5171),
.A2(n_4978),
.B(n_4889),
.Y(n_5486)
);

AO31x2_ASAP7_75t_L g5487 ( 
.A1(n_5431),
.A2(n_5064),
.A3(n_5060),
.B(n_4964),
.Y(n_5487)
);

A2O1A1Ixp33_ASAP7_75t_L g5488 ( 
.A1(n_5287),
.A2(n_4775),
.B(n_4816),
.C(n_4822),
.Y(n_5488)
);

OAI21x1_ASAP7_75t_L g5489 ( 
.A1(n_5157),
.A2(n_4747),
.B(n_4810),
.Y(n_5489)
);

AOI21xp5_ASAP7_75t_L g5490 ( 
.A1(n_5234),
.A2(n_4852),
.B(n_4862),
.Y(n_5490)
);

AO21x2_ASAP7_75t_L g5491 ( 
.A1(n_5423),
.A2(n_5046),
.B(n_4951),
.Y(n_5491)
);

AND2x2_ASAP7_75t_L g5492 ( 
.A(n_5413),
.B(n_5281),
.Y(n_5492)
);

AOI21xp5_ASAP7_75t_L g5493 ( 
.A1(n_5233),
.A2(n_5008),
.B(n_5133),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_5162),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5169),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_5181),
.Y(n_5496)
);

BUFx2_ASAP7_75t_L g5497 ( 
.A(n_5460),
.Y(n_5497)
);

INVx4_ASAP7_75t_L g5498 ( 
.A(n_5312),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_5280),
.B(n_5077),
.Y(n_5499)
);

HB1xp67_ASAP7_75t_L g5500 ( 
.A(n_5305),
.Y(n_5500)
);

AOI21xp33_ASAP7_75t_SL g5501 ( 
.A1(n_5176),
.A2(n_4921),
.B(n_4872),
.Y(n_5501)
);

INVx4_ASAP7_75t_SL g5502 ( 
.A(n_5270),
.Y(n_5502)
);

OAI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_5369),
.A2(n_4995),
.B(n_5024),
.Y(n_5503)
);

OA21x2_ASAP7_75t_L g5504 ( 
.A1(n_5367),
.A2(n_4755),
.B(n_4742),
.Y(n_5504)
);

AO21x2_ASAP7_75t_L g5505 ( 
.A1(n_5452),
.A2(n_4767),
.B(n_4766),
.Y(n_5505)
);

AOI21xp5_ASAP7_75t_L g5506 ( 
.A1(n_5208),
.A2(n_4881),
.B(n_4928),
.Y(n_5506)
);

OAI21x1_ASAP7_75t_L g5507 ( 
.A1(n_5404),
.A2(n_4747),
.B(n_4826),
.Y(n_5507)
);

NOR2xp33_ASAP7_75t_L g5508 ( 
.A(n_5432),
.B(n_5363),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_5191),
.B(n_5318),
.Y(n_5509)
);

NOR2xp33_ASAP7_75t_L g5510 ( 
.A(n_5222),
.B(n_4962),
.Y(n_5510)
);

BUFx2_ASAP7_75t_L g5511 ( 
.A(n_5176),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_5193),
.Y(n_5512)
);

AOI21xp5_ASAP7_75t_L g5513 ( 
.A1(n_5161),
.A2(n_5026),
.B(n_5075),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_5201),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_5238),
.Y(n_5515)
);

NAND2x1p5_ASAP7_75t_L g5516 ( 
.A(n_5339),
.B(n_5138),
.Y(n_5516)
);

OAI21x1_ASAP7_75t_L g5517 ( 
.A1(n_5258),
.A2(n_5039),
.B(n_4906),
.Y(n_5517)
);

INVxp67_ASAP7_75t_L g5518 ( 
.A(n_5332),
.Y(n_5518)
);

OAI21x1_ASAP7_75t_L g5519 ( 
.A1(n_5453),
.A2(n_4835),
.B(n_4975),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5183),
.Y(n_5520)
);

OAI21x1_ASAP7_75t_SL g5521 ( 
.A1(n_5294),
.A2(n_5043),
.B(n_4814),
.Y(n_5521)
);

INVx4_ASAP7_75t_L g5522 ( 
.A(n_5313),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5184),
.Y(n_5523)
);

BUFx3_ASAP7_75t_L g5524 ( 
.A(n_5264),
.Y(n_5524)
);

AOI21xp5_ASAP7_75t_L g5525 ( 
.A1(n_5230),
.A2(n_5026),
.B(n_4874),
.Y(n_5525)
);

AND2x4_ASAP7_75t_L g5526 ( 
.A(n_5236),
.B(n_4920),
.Y(n_5526)
);

AO21x2_ASAP7_75t_L g5527 ( 
.A1(n_5195),
.A2(n_4772),
.B(n_4769),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5187),
.Y(n_5528)
);

AO21x2_ASAP7_75t_L g5529 ( 
.A1(n_5436),
.A2(n_5454),
.B(n_5441),
.Y(n_5529)
);

OR2x2_ASAP7_75t_L g5530 ( 
.A(n_5283),
.B(n_4815),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5190),
.Y(n_5531)
);

NAND2xp5_ASAP7_75t_L g5532 ( 
.A(n_5343),
.B(n_5122),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5192),
.Y(n_5533)
);

OA21x2_ASAP7_75t_L g5534 ( 
.A1(n_5381),
.A2(n_4798),
.B(n_4794),
.Y(n_5534)
);

OAI21x1_ASAP7_75t_SL g5535 ( 
.A1(n_5285),
.A2(n_5418),
.B(n_5376),
.Y(n_5535)
);

OR2x2_ASAP7_75t_L g5536 ( 
.A(n_5207),
.B(n_4815),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5194),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5196),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_L g5539 ( 
.A(n_5383),
.B(n_5135),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5198),
.Y(n_5540)
);

AOI21xp5_ASAP7_75t_L g5541 ( 
.A1(n_5400),
.A2(n_5034),
.B(n_4849),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_5389),
.B(n_4925),
.Y(n_5542)
);

BUFx10_ASAP7_75t_L g5543 ( 
.A(n_5261),
.Y(n_5543)
);

OAI21x1_ASAP7_75t_SL g5544 ( 
.A1(n_5275),
.A2(n_4959),
.B(n_5047),
.Y(n_5544)
);

AO31x2_ASAP7_75t_L g5545 ( 
.A1(n_5468),
.A2(n_4783),
.A3(n_4851),
.B(n_4850),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5393),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_SL g5547 ( 
.A(n_5377),
.B(n_5065),
.Y(n_5547)
);

AOI22xp33_ASAP7_75t_L g5548 ( 
.A1(n_5174),
.A2(n_4876),
.B1(n_5032),
.B2(n_5017),
.Y(n_5548)
);

OAI21x1_ASAP7_75t_L g5549 ( 
.A1(n_5469),
.A2(n_5011),
.B(n_5080),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5221),
.Y(n_5550)
);

BUFx2_ASAP7_75t_L g5551 ( 
.A(n_5357),
.Y(n_5551)
);

OAI21xp5_ASAP7_75t_L g5552 ( 
.A1(n_5324),
.A2(n_4863),
.B(n_4877),
.Y(n_5552)
);

AND2x2_ASAP7_75t_L g5553 ( 
.A(n_5182),
.B(n_5007),
.Y(n_5553)
);

AOI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_5173),
.A2(n_4932),
.B(n_4712),
.Y(n_5554)
);

BUFx2_ASAP7_75t_L g5555 ( 
.A(n_5243),
.Y(n_5555)
);

INVx3_ASAP7_75t_L g5556 ( 
.A(n_5178),
.Y(n_5556)
);

INVx4_ASAP7_75t_SL g5557 ( 
.A(n_5380),
.Y(n_5557)
);

OAI21x1_ASAP7_75t_L g5558 ( 
.A1(n_5402),
.A2(n_5062),
.B(n_5058),
.Y(n_5558)
);

BUFx3_ASAP7_75t_L g5559 ( 
.A(n_5364),
.Y(n_5559)
);

AND2x4_ASAP7_75t_L g5560 ( 
.A(n_5229),
.B(n_5211),
.Y(n_5560)
);

AO31x2_ASAP7_75t_L g5561 ( 
.A1(n_5405),
.A2(n_4871),
.A3(n_4888),
.B(n_4875),
.Y(n_5561)
);

BUFx12f_ASAP7_75t_L g5562 ( 
.A(n_5408),
.Y(n_5562)
);

AOI22xp33_ASAP7_75t_L g5563 ( 
.A1(n_5160),
.A2(n_5041),
.B1(n_4932),
.B2(n_4697),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5246),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5253),
.Y(n_5565)
);

BUFx8_ASAP7_75t_L g5566 ( 
.A(n_5216),
.Y(n_5566)
);

INVx3_ASAP7_75t_L g5567 ( 
.A(n_5178),
.Y(n_5567)
);

NAND2xp5_ASAP7_75t_L g5568 ( 
.A(n_5330),
.B(n_4891),
.Y(n_5568)
);

NOR2xp33_ASAP7_75t_L g5569 ( 
.A(n_5442),
.B(n_5083),
.Y(n_5569)
);

AOI22xp33_ASAP7_75t_L g5570 ( 
.A1(n_5168),
.A2(n_5079),
.B1(n_5132),
.B2(n_5098),
.Y(n_5570)
);

AND2x2_ASAP7_75t_L g5571 ( 
.A(n_5242),
.B(n_5013),
.Y(n_5571)
);

BUFx6f_ASAP7_75t_L g5572 ( 
.A(n_5377),
.Y(n_5572)
);

OR2x2_ASAP7_75t_L g5573 ( 
.A(n_5300),
.B(n_4753),
.Y(n_5573)
);

INVx2_ASAP7_75t_SL g5574 ( 
.A(n_5219),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5254),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_5269),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5272),
.Y(n_5577)
);

NAND2x1p5_ASAP7_75t_L g5578 ( 
.A(n_5425),
.B(n_5094),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5320),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5266),
.Y(n_5580)
);

NAND2xp5_ASAP7_75t_L g5581 ( 
.A(n_5392),
.B(n_4899),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5248),
.Y(n_5582)
);

AO31x2_ASAP7_75t_L g5583 ( 
.A1(n_5333),
.A2(n_4976),
.A3(n_4990),
.B(n_4977),
.Y(n_5583)
);

BUFx8_ASAP7_75t_L g5584 ( 
.A(n_5260),
.Y(n_5584)
);

AOI21x1_ASAP7_75t_L g5585 ( 
.A1(n_5179),
.A2(n_4845),
.B(n_5084),
.Y(n_5585)
);

OA21x2_ASAP7_75t_L g5586 ( 
.A1(n_5231),
.A2(n_5067),
.B(n_4993),
.Y(n_5586)
);

HB1xp67_ASAP7_75t_L g5587 ( 
.A(n_5321),
.Y(n_5587)
);

AOI21xp5_ASAP7_75t_L g5588 ( 
.A1(n_5406),
.A2(n_4777),
.B(n_4741),
.Y(n_5588)
);

OA21x2_ASAP7_75t_L g5589 ( 
.A1(n_5304),
.A2(n_5437),
.B(n_5422),
.Y(n_5589)
);

AOI21xp5_ASAP7_75t_L g5590 ( 
.A1(n_5217),
.A2(n_4763),
.B(n_4759),
.Y(n_5590)
);

INVx2_ASAP7_75t_L g5591 ( 
.A(n_5250),
.Y(n_5591)
);

INVx2_ASAP7_75t_L g5592 ( 
.A(n_5257),
.Y(n_5592)
);

AOI21xp5_ASAP7_75t_L g5593 ( 
.A1(n_5217),
.A2(n_4773),
.B(n_4827),
.Y(n_5593)
);

BUFx3_ASAP7_75t_L g5594 ( 
.A(n_5219),
.Y(n_5594)
);

NAND2xp5_ASAP7_75t_SL g5595 ( 
.A(n_5390),
.B(n_5045),
.Y(n_5595)
);

AND2x4_ASAP7_75t_L g5596 ( 
.A(n_5229),
.B(n_4853),
.Y(n_5596)
);

OA21x2_ASAP7_75t_L g5597 ( 
.A1(n_5361),
.A2(n_4991),
.B(n_5048),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5349),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5368),
.Y(n_5599)
);

HB1xp67_ASAP7_75t_L g5600 ( 
.A(n_5197),
.Y(n_5600)
);

OR2x6_ASAP7_75t_L g5601 ( 
.A(n_5279),
.B(n_4782),
.Y(n_5601)
);

NAND3xp33_ASAP7_75t_L g5602 ( 
.A(n_5444),
.B(n_5370),
.C(n_5447),
.Y(n_5602)
);

AOI21xp5_ASAP7_75t_L g5603 ( 
.A1(n_5259),
.A2(n_5063),
.B(n_4829),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5374),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5375),
.Y(n_5605)
);

AND2x4_ASAP7_75t_L g5606 ( 
.A(n_5465),
.B(n_4853),
.Y(n_5606)
);

AOI22xp33_ASAP7_75t_L g5607 ( 
.A1(n_5166),
.A2(n_5114),
.B1(n_5140),
.B2(n_4714),
.Y(n_5607)
);

CKINVDCx5p33_ASAP7_75t_R g5608 ( 
.A(n_5464),
.Y(n_5608)
);

AND2x4_ASAP7_75t_L g5609 ( 
.A(n_5390),
.B(n_4858),
.Y(n_5609)
);

AOI21xp5_ASAP7_75t_L g5610 ( 
.A1(n_5172),
.A2(n_4965),
.B(n_4945),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5379),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5396),
.Y(n_5612)
);

INVx3_ASAP7_75t_L g5613 ( 
.A(n_5409),
.Y(n_5613)
);

AO31x2_ASAP7_75t_L g5614 ( 
.A1(n_5365),
.A2(n_5450),
.A3(n_5438),
.B(n_5295),
.Y(n_5614)
);

HB1xp67_ASAP7_75t_L g5615 ( 
.A(n_5382),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5397),
.Y(n_5616)
);

INVx11_ASAP7_75t_L g5617 ( 
.A(n_5323),
.Y(n_5617)
);

NAND2x1p5_ASAP7_75t_L g5618 ( 
.A(n_5308),
.B(n_5103),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_5399),
.Y(n_5619)
);

BUFx2_ASAP7_75t_L g5620 ( 
.A(n_5409),
.Y(n_5620)
);

INVx2_ASAP7_75t_L g5621 ( 
.A(n_5314),
.Y(n_5621)
);

BUFx6f_ASAP7_75t_L g5622 ( 
.A(n_5439),
.Y(n_5622)
);

NOR2xp33_ASAP7_75t_L g5623 ( 
.A(n_5348),
.B(n_5056),
.Y(n_5623)
);

AND2x2_ASAP7_75t_L g5624 ( 
.A(n_5407),
.B(n_4753),
.Y(n_5624)
);

OAI21x1_ASAP7_75t_L g5625 ( 
.A1(n_5200),
.A2(n_5057),
.B(n_4915),
.Y(n_5625)
);

AOI22xp33_ASAP7_75t_L g5626 ( 
.A1(n_5215),
.A2(n_4695),
.B1(n_5109),
.B2(n_5106),
.Y(n_5626)
);

AOI21xp5_ASAP7_75t_L g5627 ( 
.A1(n_5180),
.A2(n_5134),
.B(n_5117),
.Y(n_5627)
);

AO31x2_ASAP7_75t_L g5628 ( 
.A1(n_5296),
.A2(n_5055),
.A3(n_5128),
.B(n_4998),
.Y(n_5628)
);

OAI21x1_ASAP7_75t_L g5629 ( 
.A1(n_5175),
.A2(n_5119),
.B(n_5111),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_SL g5630 ( 
.A(n_5439),
.B(n_5040),
.Y(n_5630)
);

NAND2xp33_ASAP7_75t_L g5631 ( 
.A(n_5255),
.B(n_5076),
.Y(n_5631)
);

INVx3_ASAP7_75t_L g5632 ( 
.A(n_5463),
.Y(n_5632)
);

CKINVDCx14_ASAP7_75t_R g5633 ( 
.A(n_5241),
.Y(n_5633)
);

AOI21xp5_ASAP7_75t_L g5634 ( 
.A1(n_5203),
.A2(n_4751),
.B(n_4904),
.Y(n_5634)
);

INVx2_ASAP7_75t_L g5635 ( 
.A(n_5298),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5204),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5212),
.Y(n_5637)
);

INVx2_ASAP7_75t_L g5638 ( 
.A(n_5614),
.Y(n_5638)
);

OAI21x1_ASAP7_75t_L g5639 ( 
.A1(n_5507),
.A2(n_5225),
.B(n_5188),
.Y(n_5639)
);

CKINVDCx20_ASAP7_75t_R g5640 ( 
.A(n_5502),
.Y(n_5640)
);

INVx4_ASAP7_75t_SL g5641 ( 
.A(n_5477),
.Y(n_5641)
);

INVx2_ASAP7_75t_L g5642 ( 
.A(n_5614),
.Y(n_5642)
);

INVx2_ASAP7_75t_L g5643 ( 
.A(n_5615),
.Y(n_5643)
);

AND2x2_ASAP7_75t_L g5644 ( 
.A(n_5492),
.B(n_5401),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5600),
.Y(n_5645)
);

INVx2_ASAP7_75t_L g5646 ( 
.A(n_5485),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5579),
.Y(n_5647)
);

AND2x4_ASAP7_75t_L g5648 ( 
.A(n_5500),
.B(n_5338),
.Y(n_5648)
);

INVx2_ASAP7_75t_SL g5649 ( 
.A(n_5524),
.Y(n_5649)
);

AND2x2_ASAP7_75t_L g5650 ( 
.A(n_5587),
.B(n_5163),
.Y(n_5650)
);

INVx2_ASAP7_75t_L g5651 ( 
.A(n_5494),
.Y(n_5651)
);

BUFx3_ASAP7_75t_L g5652 ( 
.A(n_5511),
.Y(n_5652)
);

INVx3_ASAP7_75t_L g5653 ( 
.A(n_5606),
.Y(n_5653)
);

INVx2_ASAP7_75t_SL g5654 ( 
.A(n_5551),
.Y(n_5654)
);

OR2x2_ASAP7_75t_L g5655 ( 
.A(n_5636),
.B(n_5223),
.Y(n_5655)
);

NOR2xp33_ASAP7_75t_L g5656 ( 
.A(n_5498),
.B(n_5387),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_5496),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5555),
.B(n_5298),
.Y(n_5658)
);

AND2x2_ASAP7_75t_L g5659 ( 
.A(n_5637),
.B(n_5298),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5481),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_5512),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_5474),
.B(n_5220),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_5495),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5520),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5523),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5528),
.Y(n_5666)
);

INVx2_ASAP7_75t_L g5667 ( 
.A(n_5514),
.Y(n_5667)
);

INVx1_ASAP7_75t_L g5668 ( 
.A(n_5531),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5533),
.Y(n_5669)
);

OR2x2_ASAP7_75t_L g5670 ( 
.A(n_5476),
.B(n_5214),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5537),
.Y(n_5671)
);

NAND2x1p5_ASAP7_75t_L g5672 ( 
.A(n_5522),
.B(n_5424),
.Y(n_5672)
);

NOR2xp33_ASAP7_75t_L g5673 ( 
.A(n_5608),
.B(n_5463),
.Y(n_5673)
);

INVx3_ASAP7_75t_L g5674 ( 
.A(n_5560),
.Y(n_5674)
);

INVx2_ASAP7_75t_L g5675 ( 
.A(n_5515),
.Y(n_5675)
);

INVx3_ASAP7_75t_SL g5676 ( 
.A(n_5502),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5538),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_5540),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5550),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5564),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5565),
.Y(n_5681)
);

OA21x2_ASAP7_75t_L g5682 ( 
.A1(n_5483),
.A2(n_5159),
.B(n_5306),
.Y(n_5682)
);

INVx3_ASAP7_75t_L g5683 ( 
.A(n_5572),
.Y(n_5683)
);

CKINVDCx20_ASAP7_75t_R g5684 ( 
.A(n_5559),
.Y(n_5684)
);

OAI21xp33_ASAP7_75t_SL g5685 ( 
.A1(n_5617),
.A2(n_5279),
.B(n_5185),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5582),
.Y(n_5686)
);

AND2x2_ASAP7_75t_L g5687 ( 
.A(n_5571),
.B(n_5298),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5530),
.Y(n_5688)
);

OR2x2_ASAP7_75t_L g5689 ( 
.A(n_5472),
.B(n_5580),
.Y(n_5689)
);

AO21x2_ASAP7_75t_L g5690 ( 
.A1(n_5473),
.A2(n_5337),
.B(n_5252),
.Y(n_5690)
);

INVx3_ASAP7_75t_L g5691 ( 
.A(n_5572),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5575),
.Y(n_5692)
);

BUFx2_ASAP7_75t_L g5693 ( 
.A(n_5620),
.Y(n_5693)
);

AOI22xp33_ASAP7_75t_L g5694 ( 
.A1(n_5602),
.A2(n_5177),
.B1(n_5218),
.B2(n_5213),
.Y(n_5694)
);

INVx2_ASAP7_75t_L g5695 ( 
.A(n_5591),
.Y(n_5695)
);

AND2x2_ASAP7_75t_L g5696 ( 
.A(n_5475),
.B(n_5443),
.Y(n_5696)
);

OAI21xp33_ASAP7_75t_SL g5697 ( 
.A1(n_5508),
.A2(n_5251),
.B(n_5282),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5576),
.Y(n_5698)
);

HB1xp67_ASAP7_75t_L g5699 ( 
.A(n_5592),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_L g5700 ( 
.A(n_5624),
.B(n_5573),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_5530),
.Y(n_5701)
);

OAI21x1_ASAP7_75t_L g5702 ( 
.A1(n_5489),
.A2(n_5256),
.B(n_5240),
.Y(n_5702)
);

INVx1_ASAP7_75t_SL g5703 ( 
.A(n_5497),
.Y(n_5703)
);

AND2x2_ASAP7_75t_L g5704 ( 
.A(n_5553),
.B(n_5457),
.Y(n_5704)
);

INVx1_ASAP7_75t_SL g5705 ( 
.A(n_5594),
.Y(n_5705)
);

AND2x2_ASAP7_75t_L g5706 ( 
.A(n_5518),
.B(n_5355),
.Y(n_5706)
);

HB1xp67_ASAP7_75t_L g5707 ( 
.A(n_5621),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5577),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5546),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_5598),
.Y(n_5710)
);

INVx1_ASAP7_75t_SL g5711 ( 
.A(n_5526),
.Y(n_5711)
);

INVx4_ASAP7_75t_L g5712 ( 
.A(n_5557),
.Y(n_5712)
);

INVx2_ASAP7_75t_SL g5713 ( 
.A(n_5566),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5599),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_5633),
.B(n_5378),
.Y(n_5715)
);

AND2x2_ASAP7_75t_L g5716 ( 
.A(n_5509),
.B(n_5459),
.Y(n_5716)
);

OAI21x1_ASAP7_75t_L g5717 ( 
.A1(n_5625),
.A2(n_5373),
.B(n_5268),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5604),
.Y(n_5718)
);

HB1xp67_ASAP7_75t_SL g5719 ( 
.A(n_5584),
.Y(n_5719)
);

BUFx3_ASAP7_75t_L g5720 ( 
.A(n_5562),
.Y(n_5720)
);

OR2x6_ASAP7_75t_L g5721 ( 
.A(n_5516),
.B(n_5345),
.Y(n_5721)
);

AND2x2_ASAP7_75t_L g5722 ( 
.A(n_5605),
.B(n_5384),
.Y(n_5722)
);

OR2x6_ASAP7_75t_L g5723 ( 
.A(n_5601),
.B(n_5356),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_5611),
.B(n_5429),
.Y(n_5724)
);

HB1xp67_ASAP7_75t_L g5725 ( 
.A(n_5597),
.Y(n_5725)
);

OAI21x1_ASAP7_75t_L g5726 ( 
.A1(n_5573),
.A2(n_5414),
.B(n_5366),
.Y(n_5726)
);

INVx1_ASAP7_75t_L g5727 ( 
.A(n_5612),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_5529),
.Y(n_5728)
);

INVx2_ASAP7_75t_L g5729 ( 
.A(n_5616),
.Y(n_5729)
);

INVx3_ASAP7_75t_L g5730 ( 
.A(n_5622),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5619),
.Y(n_5731)
);

BUFx2_ASAP7_75t_SL g5732 ( 
.A(n_5622),
.Y(n_5732)
);

INVx1_ASAP7_75t_SL g5733 ( 
.A(n_5557),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5536),
.Y(n_5734)
);

OAI21xp5_ASAP7_75t_L g5735 ( 
.A1(n_5488),
.A2(n_5288),
.B(n_5227),
.Y(n_5735)
);

INVx2_ASAP7_75t_L g5736 ( 
.A(n_5536),
.Y(n_5736)
);

OAI21x1_ASAP7_75t_L g5737 ( 
.A1(n_5558),
.A2(n_5362),
.B(n_5235),
.Y(n_5737)
);

NAND2xp5_ASAP7_75t_L g5738 ( 
.A(n_5479),
.B(n_5247),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5542),
.Y(n_5739)
);

NAND2xp5_ASAP7_75t_L g5740 ( 
.A(n_5568),
.B(n_5247),
.Y(n_5740)
);

NOR2xp33_ASAP7_75t_L g5741 ( 
.A(n_5623),
.B(n_5291),
.Y(n_5741)
);

BUFx6f_ASAP7_75t_L g5742 ( 
.A(n_5574),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5635),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5504),
.Y(n_5744)
);

BUFx2_ASAP7_75t_L g5745 ( 
.A(n_5613),
.Y(n_5745)
);

INVx2_ASAP7_75t_L g5746 ( 
.A(n_5534),
.Y(n_5746)
);

HB1xp67_ASAP7_75t_L g5747 ( 
.A(n_5583),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5581),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5583),
.Y(n_5749)
);

BUFx2_ASAP7_75t_SL g5750 ( 
.A(n_5632),
.Y(n_5750)
);

BUFx2_ASAP7_75t_L g5751 ( 
.A(n_5556),
.Y(n_5751)
);

OAI21xp5_ASAP7_75t_L g5752 ( 
.A1(n_5554),
.A2(n_5263),
.B(n_5289),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_5609),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5527),
.Y(n_5754)
);

INVx2_ASAP7_75t_L g5755 ( 
.A(n_5561),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5561),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5596),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5567),
.Y(n_5758)
);

BUFx2_ASAP7_75t_L g5759 ( 
.A(n_5586),
.Y(n_5759)
);

INVx2_ASAP7_75t_L g5760 ( 
.A(n_5487),
.Y(n_5760)
);

OAI221xp5_ASAP7_75t_L g5761 ( 
.A1(n_5685),
.A2(n_5548),
.B1(n_5631),
.B2(n_5563),
.C(n_5570),
.Y(n_5761)
);

OAI21x1_ASAP7_75t_L g5762 ( 
.A1(n_5746),
.A2(n_5585),
.B(n_5513),
.Y(n_5762)
);

AOI22xp33_ASAP7_75t_L g5763 ( 
.A1(n_5690),
.A2(n_5601),
.B1(n_5544),
.B2(n_5521),
.Y(n_5763)
);

OAI22xp5_ASAP7_75t_L g5764 ( 
.A1(n_5723),
.A2(n_5501),
.B1(n_5539),
.B2(n_5482),
.Y(n_5764)
);

AOI22xp33_ASAP7_75t_L g5765 ( 
.A1(n_5694),
.A2(n_5503),
.B1(n_5626),
.B2(n_5493),
.Y(n_5765)
);

OAI22xp33_ASAP7_75t_L g5766 ( 
.A1(n_5723),
.A2(n_5654),
.B1(n_5759),
.B2(n_5721),
.Y(n_5766)
);

AOI22xp33_ASAP7_75t_L g5767 ( 
.A1(n_5752),
.A2(n_5735),
.B1(n_5697),
.B2(n_5741),
.Y(n_5767)
);

AOI22xp33_ASAP7_75t_L g5768 ( 
.A1(n_5687),
.A2(n_5757),
.B1(n_5535),
.B2(n_5725),
.Y(n_5768)
);

AND2x2_ASAP7_75t_L g5769 ( 
.A(n_5674),
.B(n_5510),
.Y(n_5769)
);

OAI22xp5_ASAP7_75t_L g5770 ( 
.A1(n_5721),
.A2(n_5499),
.B1(n_5618),
.B2(n_5532),
.Y(n_5770)
);

AOI21xp5_ASAP7_75t_L g5771 ( 
.A1(n_5649),
.A2(n_5490),
.B(n_5426),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5647),
.Y(n_5772)
);

AND2x4_ASAP7_75t_L g5773 ( 
.A(n_5653),
.B(n_5487),
.Y(n_5773)
);

BUFx2_ASAP7_75t_L g5774 ( 
.A(n_5641),
.Y(n_5774)
);

NAND2xp5_ASAP7_75t_L g5775 ( 
.A(n_5740),
.B(n_5545),
.Y(n_5775)
);

OAI22xp33_ASAP7_75t_L g5776 ( 
.A1(n_5712),
.A2(n_5589),
.B1(n_5541),
.B2(n_5578),
.Y(n_5776)
);

AOI22xp33_ASAP7_75t_SL g5777 ( 
.A1(n_5652),
.A2(n_5491),
.B1(n_5505),
.B2(n_5428),
.Y(n_5777)
);

NAND2xp5_ASAP7_75t_L g5778 ( 
.A(n_5688),
.B(n_5545),
.Y(n_5778)
);

AND2x2_ASAP7_75t_L g5779 ( 
.A(n_5674),
.B(n_5569),
.Y(n_5779)
);

OAI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_5712),
.A2(n_5595),
.B1(n_5630),
.B2(n_5307),
.Y(n_5780)
);

AOI22xp33_ASAP7_75t_L g5781 ( 
.A1(n_5650),
.A2(n_5547),
.B1(n_5634),
.B2(n_5588),
.Y(n_5781)
);

OAI221xp5_ASAP7_75t_L g5782 ( 
.A1(n_5676),
.A2(n_5552),
.B1(n_5353),
.B2(n_5607),
.C(n_5610),
.Y(n_5782)
);

BUFx3_ASAP7_75t_L g5783 ( 
.A(n_5640),
.Y(n_5783)
);

AOI21xp5_ASAP7_75t_L g5784 ( 
.A1(n_5744),
.A2(n_5525),
.B(n_5486),
.Y(n_5784)
);

INVx3_ASAP7_75t_L g5785 ( 
.A(n_5733),
.Y(n_5785)
);

OA21x2_ASAP7_75t_L g5786 ( 
.A1(n_5744),
.A2(n_5629),
.B(n_5593),
.Y(n_5786)
);

AOI22xp33_ASAP7_75t_L g5787 ( 
.A1(n_5645),
.A2(n_5331),
.B1(n_5627),
.B2(n_5448),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5647),
.Y(n_5788)
);

OAI21x1_ASAP7_75t_L g5789 ( 
.A1(n_5760),
.A2(n_5478),
.B(n_5549),
.Y(n_5789)
);

OAI22xp5_ASAP7_75t_L g5790 ( 
.A1(n_5672),
.A2(n_5346),
.B1(n_5434),
.B2(n_5394),
.Y(n_5790)
);

OAI22xp5_ASAP7_75t_L g5791 ( 
.A1(n_5750),
.A2(n_5284),
.B1(n_5590),
.B2(n_5372),
.Y(n_5791)
);

AOI22xp33_ASAP7_75t_L g5792 ( 
.A1(n_5648),
.A2(n_5739),
.B1(n_5653),
.B2(n_5644),
.Y(n_5792)
);

AOI22xp33_ASAP7_75t_L g5793 ( 
.A1(n_5648),
.A2(n_5299),
.B1(n_5358),
.B2(n_5371),
.Y(n_5793)
);

AOI221xp5_ASAP7_75t_L g5794 ( 
.A1(n_5749),
.A2(n_5419),
.B1(n_5471),
.B2(n_5398),
.C(n_5351),
.Y(n_5794)
);

BUFx6f_ASAP7_75t_L g5795 ( 
.A(n_5713),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5664),
.Y(n_5796)
);

BUFx2_ASAP7_75t_L g5797 ( 
.A(n_5641),
.Y(n_5797)
);

AND2x2_ASAP7_75t_L g5798 ( 
.A(n_5693),
.B(n_5628),
.Y(n_5798)
);

INVx1_ASAP7_75t_SL g5799 ( 
.A(n_5719),
.Y(n_5799)
);

AOI22xp33_ASAP7_75t_L g5800 ( 
.A1(n_5706),
.A2(n_5299),
.B1(n_5371),
.B2(n_5205),
.Y(n_5800)
);

AND2x2_ASAP7_75t_L g5801 ( 
.A(n_5643),
.B(n_5628),
.Y(n_5801)
);

INVx3_ASAP7_75t_L g5802 ( 
.A(n_5742),
.Y(n_5802)
);

INVx3_ASAP7_75t_L g5803 ( 
.A(n_5742),
.Y(n_5803)
);

OAI22xp33_ASAP7_75t_L g5804 ( 
.A1(n_5711),
.A2(n_5506),
.B1(n_5286),
.B2(n_5262),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5722),
.B(n_5543),
.Y(n_5805)
);

BUFx6f_ASAP7_75t_L g5806 ( 
.A(n_5720),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5699),
.Y(n_5807)
);

AOI22xp33_ASAP7_75t_L g5808 ( 
.A1(n_5748),
.A2(n_5354),
.B1(n_5262),
.B2(n_5302),
.Y(n_5808)
);

OAI22xp5_ASAP7_75t_L g5809 ( 
.A1(n_5750),
.A2(n_5412),
.B1(n_5451),
.B2(n_5385),
.Y(n_5809)
);

AOI221xp5_ASAP7_75t_L g5810 ( 
.A1(n_5747),
.A2(n_5603),
.B1(n_5446),
.B2(n_5352),
.C(n_5470),
.Y(n_5810)
);

INVx2_ASAP7_75t_L g5811 ( 
.A(n_5707),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_5638),
.A2(n_5517),
.B(n_5519),
.Y(n_5812)
);

AOI221xp5_ASAP7_75t_L g5813 ( 
.A1(n_5738),
.A2(n_5360),
.B1(n_5315),
.B2(n_5244),
.C(n_5359),
.Y(n_5813)
);

NOR2xp33_ASAP7_75t_L g5814 ( 
.A(n_5684),
.B(n_5326),
.Y(n_5814)
);

NOR2xp33_ASAP7_75t_L g5815 ( 
.A(n_5703),
.B(n_5386),
.Y(n_5815)
);

AOI22xp33_ASAP7_75t_L g5816 ( 
.A1(n_5656),
.A2(n_5302),
.B1(n_5286),
.B2(n_5411),
.Y(n_5816)
);

OAI211xp5_ASAP7_75t_L g5817 ( 
.A1(n_5715),
.A2(n_5249),
.B(n_5705),
.C(n_5745),
.Y(n_5817)
);

AOI22xp33_ASAP7_75t_L g5818 ( 
.A1(n_5696),
.A2(n_5462),
.B1(n_5440),
.B2(n_5158),
.Y(n_5818)
);

OAI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_5751),
.A2(n_5445),
.B1(n_5165),
.B2(n_5277),
.Y(n_5819)
);

INVxp67_ASAP7_75t_L g5820 ( 
.A(n_5673),
.Y(n_5820)
);

OAI22xp5_ASAP7_75t_L g5821 ( 
.A1(n_5670),
.A2(n_5189),
.B1(n_5210),
.B2(n_5301),
.Y(n_5821)
);

OAI22xp5_ASAP7_75t_L g5822 ( 
.A1(n_5689),
.A2(n_5388),
.B1(n_5417),
.B2(n_5290),
.Y(n_5822)
);

OR2x2_ASAP7_75t_L g5823 ( 
.A(n_5700),
.B(n_4858),
.Y(n_5823)
);

AOI21xp5_ASAP7_75t_L g5824 ( 
.A1(n_5726),
.A2(n_5311),
.B(n_5449),
.Y(n_5824)
);

OAI21xp33_ASAP7_75t_SL g5825 ( 
.A1(n_5658),
.A2(n_5737),
.B(n_5701),
.Y(n_5825)
);

AOI22xp33_ASAP7_75t_L g5826 ( 
.A1(n_5704),
.A2(n_5336),
.B1(n_5290),
.B2(n_5224),
.Y(n_5826)
);

AOI22xp5_ASAP7_75t_L g5827 ( 
.A1(n_5724),
.A2(n_5336),
.B1(n_5433),
.B2(n_5325),
.Y(n_5827)
);

AOI22xp33_ASAP7_75t_L g5828 ( 
.A1(n_5716),
.A2(n_5484),
.B1(n_5325),
.B2(n_5293),
.Y(n_5828)
);

AOI22xp33_ASAP7_75t_L g5829 ( 
.A1(n_5688),
.A2(n_5293),
.B1(n_5467),
.B2(n_5415),
.Y(n_5829)
);

AOI22xp33_ASAP7_75t_L g5830 ( 
.A1(n_5701),
.A2(n_5344),
.B1(n_5239),
.B2(n_5466),
.Y(n_5830)
);

AOI22xp33_ASAP7_75t_L g5831 ( 
.A1(n_5758),
.A2(n_5104),
.B1(n_5089),
.B2(n_5059),
.Y(n_5831)
);

NAND2xp5_ASAP7_75t_L g5832 ( 
.A(n_5734),
.B(n_5186),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5743),
.Y(n_5833)
);

OAI211xp5_ASAP7_75t_L g5834 ( 
.A1(n_5754),
.A2(n_4969),
.B(n_4912),
.C(n_5435),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5664),
.Y(n_5835)
);

INVx3_ASAP7_75t_L g5836 ( 
.A(n_5742),
.Y(n_5836)
);

OAI221xp5_ASAP7_75t_L g5837 ( 
.A1(n_5662),
.A2(n_5420),
.B1(n_5149),
.B2(n_5156),
.C(n_5152),
.Y(n_5837)
);

AND2x2_ASAP7_75t_L g5838 ( 
.A(n_5753),
.B(n_5480),
.Y(n_5838)
);

NAND2xp5_ASAP7_75t_L g5839 ( 
.A(n_5736),
.B(n_5186),
.Y(n_5839)
);

AOI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5659),
.A2(n_5139),
.B1(n_5136),
.B2(n_5150),
.Y(n_5840)
);

AND2x2_ASAP7_75t_L g5841 ( 
.A(n_5646),
.B(n_4812),
.Y(n_5841)
);

INVx2_ASAP7_75t_L g5842 ( 
.A(n_5743),
.Y(n_5842)
);

OAI22xp5_ASAP7_75t_L g5843 ( 
.A1(n_5655),
.A2(n_4922),
.B1(n_5116),
.B2(n_5110),
.Y(n_5843)
);

OAI21x1_ASAP7_75t_L g5844 ( 
.A1(n_5642),
.A2(n_5403),
.B(n_5226),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5710),
.Y(n_5845)
);

AOI221xp5_ASAP7_75t_L g5846 ( 
.A1(n_5660),
.A2(n_5130),
.B1(n_5015),
.B2(n_5014),
.C(n_5427),
.Y(n_5846)
);

AOI21x1_ASAP7_75t_L g5847 ( 
.A1(n_5728),
.A2(n_5232),
.B(n_5267),
.Y(n_5847)
);

OAI22xp5_ASAP7_75t_L g5848 ( 
.A1(n_5732),
.A2(n_5427),
.B1(n_4952),
.B2(n_5410),
.Y(n_5848)
);

OAI22xp33_ASAP7_75t_L g5849 ( 
.A1(n_5683),
.A2(n_4952),
.B1(n_5410),
.B2(n_5430),
.Y(n_5849)
);

OAI22xp33_ASAP7_75t_L g5850 ( 
.A1(n_5683),
.A2(n_5430),
.B1(n_5341),
.B2(n_4926),
.Y(n_5850)
);

OAI221xp5_ASAP7_75t_L g5851 ( 
.A1(n_5755),
.A2(n_5341),
.B1(n_5129),
.B2(n_5087),
.C(n_4926),
.Y(n_5851)
);

AOI22xp33_ASAP7_75t_SL g5852 ( 
.A1(n_5732),
.A2(n_5416),
.B1(n_5421),
.B2(n_5395),
.Y(n_5852)
);

AOI211xp5_ASAP7_75t_L g5853 ( 
.A1(n_5717),
.A2(n_5342),
.B(n_5209),
.C(n_5303),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5710),
.Y(n_5854)
);

OAI21x1_ASAP7_75t_L g5855 ( 
.A1(n_5756),
.A2(n_5316),
.B(n_5310),
.Y(n_5855)
);

AOI22xp33_ASAP7_75t_L g5856 ( 
.A1(n_5729),
.A2(n_5665),
.B1(n_5666),
.B2(n_5663),
.Y(n_5856)
);

OAI21x1_ASAP7_75t_L g5857 ( 
.A1(n_5639),
.A2(n_5702),
.B(n_5657),
.Y(n_5857)
);

INVx2_ASAP7_75t_SL g5858 ( 
.A(n_5691),
.Y(n_5858)
);

OAI22xp5_ASAP7_75t_L g5859 ( 
.A1(n_5691),
.A2(n_4890),
.B1(n_4812),
.B2(n_5087),
.Y(n_5859)
);

AND2x2_ASAP7_75t_L g5860 ( 
.A(n_5792),
.B(n_5730),
.Y(n_5860)
);

INVx2_ASAP7_75t_L g5861 ( 
.A(n_5807),
.Y(n_5861)
);

NAND2xp5_ASAP7_75t_L g5862 ( 
.A(n_5801),
.B(n_5668),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5811),
.Y(n_5863)
);

INVx2_ASAP7_75t_L g5864 ( 
.A(n_5833),
.Y(n_5864)
);

INVx2_ASAP7_75t_L g5865 ( 
.A(n_5842),
.Y(n_5865)
);

BUFx3_ASAP7_75t_L g5866 ( 
.A(n_5795),
.Y(n_5866)
);

AOI22xp33_ASAP7_75t_L g5867 ( 
.A1(n_5761),
.A2(n_5682),
.B1(n_5730),
.B2(n_5671),
.Y(n_5867)
);

INVx2_ASAP7_75t_L g5868 ( 
.A(n_5772),
.Y(n_5868)
);

AOI22xp33_ASAP7_75t_L g5869 ( 
.A1(n_5767),
.A2(n_5682),
.B1(n_5677),
.B2(n_5678),
.Y(n_5869)
);

INVx2_ASAP7_75t_SL g5870 ( 
.A(n_5795),
.Y(n_5870)
);

INVx2_ASAP7_75t_L g5871 ( 
.A(n_5788),
.Y(n_5871)
);

INVx1_ASAP7_75t_SL g5872 ( 
.A(n_5799),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5796),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5835),
.Y(n_5874)
);

AND2x4_ASAP7_75t_L g5875 ( 
.A(n_5774),
.B(n_5669),
.Y(n_5875)
);

AND2x2_ASAP7_75t_L g5876 ( 
.A(n_5798),
.B(n_5769),
.Y(n_5876)
);

NOR2xp33_ASAP7_75t_L g5877 ( 
.A(n_5795),
.B(n_5679),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5845),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5854),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5778),
.Y(n_5880)
);

AND2x2_ASAP7_75t_L g5881 ( 
.A(n_5779),
.B(n_5680),
.Y(n_5881)
);

AOI22xp33_ASAP7_75t_L g5882 ( 
.A1(n_5765),
.A2(n_5692),
.B1(n_5698),
.B2(n_5681),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5832),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5839),
.Y(n_5884)
);

AND2x2_ASAP7_75t_L g5885 ( 
.A(n_5785),
.B(n_5708),
.Y(n_5885)
);

INVx2_ASAP7_75t_L g5886 ( 
.A(n_5857),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5823),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5802),
.B(n_5709),
.Y(n_5888)
);

HB1xp67_ASAP7_75t_L g5889 ( 
.A(n_5775),
.Y(n_5889)
);

BUFx6f_ASAP7_75t_L g5890 ( 
.A(n_5806),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5841),
.Y(n_5891)
);

AND2x2_ASAP7_75t_L g5892 ( 
.A(n_5836),
.B(n_5714),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5856),
.Y(n_5893)
);

NOR2xp67_ASAP7_75t_L g5894 ( 
.A(n_5825),
.B(n_5651),
.Y(n_5894)
);

INVx2_ASAP7_75t_L g5895 ( 
.A(n_5786),
.Y(n_5895)
);

AND2x2_ASAP7_75t_L g5896 ( 
.A(n_5773),
.B(n_5718),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5838),
.Y(n_5897)
);

INVx3_ASAP7_75t_L g5898 ( 
.A(n_5797),
.Y(n_5898)
);

NOR2xp33_ASAP7_75t_L g5899 ( 
.A(n_5806),
.B(n_5727),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5773),
.Y(n_5900)
);

NOR2x1_ASAP7_75t_L g5901 ( 
.A(n_5766),
.B(n_5731),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5786),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5770),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_L g5904 ( 
.A(n_5784),
.B(n_5661),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_5847),
.Y(n_5905)
);

OR2x2_ASAP7_75t_L g5906 ( 
.A(n_5858),
.B(n_5667),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5762),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5768),
.B(n_5675),
.Y(n_5908)
);

INVx2_ASAP7_75t_L g5909 ( 
.A(n_5812),
.Y(n_5909)
);

INVx2_ASAP7_75t_L g5910 ( 
.A(n_5803),
.Y(n_5910)
);

NAND2xp5_ASAP7_75t_L g5911 ( 
.A(n_5781),
.B(n_5686),
.Y(n_5911)
);

AND2x4_ASAP7_75t_L g5912 ( 
.A(n_5783),
.B(n_5695),
.Y(n_5912)
);

INVxp67_ASAP7_75t_SL g5913 ( 
.A(n_5771),
.Y(n_5913)
);

AND2x2_ASAP7_75t_L g5914 ( 
.A(n_5803),
.B(n_4989),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5844),
.Y(n_5915)
);

HB1xp67_ASAP7_75t_L g5916 ( 
.A(n_5820),
.Y(n_5916)
);

AND2x4_ASAP7_75t_L g5917 ( 
.A(n_5805),
.B(n_5206),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5789),
.Y(n_5918)
);

INVx3_ASAP7_75t_L g5919 ( 
.A(n_5806),
.Y(n_5919)
);

AND2x2_ASAP7_75t_L g5920 ( 
.A(n_5764),
.B(n_5003),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_5817),
.Y(n_5921)
);

AOI22xp33_ASAP7_75t_L g5922 ( 
.A1(n_5763),
.A2(n_5274),
.B1(n_5350),
.B2(n_5347),
.Y(n_5922)
);

AND2x4_ASAP7_75t_L g5923 ( 
.A(n_5818),
.B(n_5003),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5851),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_5776),
.B(n_5129),
.Y(n_5925)
);

NAND2xp5_ASAP7_75t_L g5926 ( 
.A(n_5826),
.B(n_4890),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5859),
.Y(n_5927)
);

HB1xp67_ASAP7_75t_L g5928 ( 
.A(n_5780),
.Y(n_5928)
);

AND2x2_ASAP7_75t_L g5929 ( 
.A(n_5815),
.B(n_4694),
.Y(n_5929)
);

INVxp67_ASAP7_75t_SL g5930 ( 
.A(n_5804),
.Y(n_5930)
);

OR2x2_ASAP7_75t_L g5931 ( 
.A(n_5800),
.B(n_4694),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5777),
.B(n_5319),
.Y(n_5932)
);

INVx2_ASAP7_75t_L g5933 ( 
.A(n_5855),
.Y(n_5933)
);

NAND2xp5_ASAP7_75t_L g5934 ( 
.A(n_5921),
.B(n_5787),
.Y(n_5934)
);

AND2x2_ASAP7_75t_L g5935 ( 
.A(n_5876),
.B(n_5840),
.Y(n_5935)
);

NAND2xp5_ASAP7_75t_L g5936 ( 
.A(n_5924),
.B(n_5824),
.Y(n_5936)
);

HB1xp67_ASAP7_75t_L g5937 ( 
.A(n_5916),
.Y(n_5937)
);

BUFx2_ASAP7_75t_L g5938 ( 
.A(n_5890),
.Y(n_5938)
);

AND2x2_ASAP7_75t_L g5939 ( 
.A(n_5860),
.B(n_5814),
.Y(n_5939)
);

AND2x4_ASAP7_75t_SL g5940 ( 
.A(n_5890),
.B(n_5831),
.Y(n_5940)
);

AND2x2_ASAP7_75t_L g5941 ( 
.A(n_5898),
.B(n_5828),
.Y(n_5941)
);

AND2x2_ASAP7_75t_L g5942 ( 
.A(n_5898),
.B(n_5853),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_L g5943 ( 
.A(n_5928),
.B(n_5816),
.Y(n_5943)
);

AND2x2_ASAP7_75t_L g5944 ( 
.A(n_5870),
.B(n_5793),
.Y(n_5944)
);

INVx1_ASAP7_75t_SL g5945 ( 
.A(n_5872),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5861),
.Y(n_5946)
);

OR2x2_ASAP7_75t_L g5947 ( 
.A(n_5887),
.B(n_5821),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_5863),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5927),
.B(n_5827),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5873),
.Y(n_5950)
);

OAI22xp5_ASAP7_75t_L g5951 ( 
.A1(n_5867),
.A2(n_5782),
.B1(n_5829),
.B2(n_5791),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5874),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5868),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5871),
.Y(n_5954)
);

AND2x2_ASAP7_75t_L g5955 ( 
.A(n_5919),
.B(n_5830),
.Y(n_5955)
);

OR2x2_ASAP7_75t_L g5956 ( 
.A(n_5911),
.B(n_5822),
.Y(n_5956)
);

AND2x2_ASAP7_75t_L g5957 ( 
.A(n_5919),
.B(n_5808),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5878),
.Y(n_5958)
);

INVx1_ASAP7_75t_SL g5959 ( 
.A(n_5872),
.Y(n_5959)
);

AND2x4_ASAP7_75t_L g5960 ( 
.A(n_5866),
.B(n_5329),
.Y(n_5960)
);

INVx1_ASAP7_75t_L g5961 ( 
.A(n_5879),
.Y(n_5961)
);

AND2x4_ASAP7_75t_L g5962 ( 
.A(n_5875),
.B(n_5322),
.Y(n_5962)
);

NAND2xp5_ASAP7_75t_L g5963 ( 
.A(n_5930),
.B(n_5810),
.Y(n_5963)
);

NOR2x1_ASAP7_75t_L g5964 ( 
.A(n_5890),
.B(n_5809),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5862),
.Y(n_5965)
);

HB1xp67_ASAP7_75t_L g5966 ( 
.A(n_5904),
.Y(n_5966)
);

AND2x2_ASAP7_75t_L g5967 ( 
.A(n_5908),
.B(n_5852),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5903),
.B(n_5813),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5862),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5880),
.Y(n_5970)
);

NAND2xp5_ASAP7_75t_L g5971 ( 
.A(n_5893),
.B(n_5923),
.Y(n_5971)
);

INVx1_ASAP7_75t_L g5972 ( 
.A(n_5889),
.Y(n_5972)
);

INVxp67_ASAP7_75t_SL g5973 ( 
.A(n_5904),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5864),
.Y(n_5974)
);

AND2x2_ASAP7_75t_L g5975 ( 
.A(n_5913),
.B(n_5819),
.Y(n_5975)
);

NAND3xp33_ASAP7_75t_L g5976 ( 
.A(n_5907),
.B(n_5848),
.C(n_5794),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_L g5977 ( 
.A(n_5923),
.B(n_5882),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5881),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5911),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5883),
.Y(n_5980)
);

OR2x2_ASAP7_75t_L g5981 ( 
.A(n_5884),
.B(n_5849),
.Y(n_5981)
);

OR2x2_ASAP7_75t_L g5982 ( 
.A(n_5891),
.B(n_5850),
.Y(n_5982)
);

AND2x2_ASAP7_75t_L g5983 ( 
.A(n_5875),
.B(n_5790),
.Y(n_5983)
);

OR2x2_ASAP7_75t_L g5984 ( 
.A(n_5931),
.B(n_5834),
.Y(n_5984)
);

INVx3_ASAP7_75t_L g5985 ( 
.A(n_5912),
.Y(n_5985)
);

NOR3xp33_ASAP7_75t_L g5986 ( 
.A(n_5932),
.B(n_5837),
.C(n_5846),
.Y(n_5986)
);

AND2x2_ASAP7_75t_L g5987 ( 
.A(n_5896),
.B(n_5843),
.Y(n_5987)
);

AND2x2_ASAP7_75t_L g5988 ( 
.A(n_5929),
.B(n_5271),
.Y(n_5988)
);

INVxp67_ASAP7_75t_SL g5989 ( 
.A(n_5901),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5885),
.Y(n_5990)
);

OR2x2_ASAP7_75t_L g5991 ( 
.A(n_5926),
.B(n_5925),
.Y(n_5991)
);

OAI22xp5_ASAP7_75t_L g5992 ( 
.A1(n_5894),
.A2(n_5265),
.B1(n_5297),
.B2(n_5276),
.Y(n_5992)
);

AND2x2_ASAP7_75t_L g5993 ( 
.A(n_5901),
.B(n_5334),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5917),
.B(n_5335),
.Y(n_5994)
);

NAND2xp5_ASAP7_75t_L g5995 ( 
.A(n_5926),
.B(n_5920),
.Y(n_5995)
);

NAND2xp5_ASAP7_75t_L g5996 ( 
.A(n_5869),
.B(n_5327),
.Y(n_5996)
);

NAND3xp33_ASAP7_75t_L g5997 ( 
.A(n_5925),
.B(n_75),
.C(n_76),
.Y(n_5997)
);

AND2x2_ASAP7_75t_L g5998 ( 
.A(n_5917),
.B(n_5328),
.Y(n_5998)
);

NAND2xp5_ASAP7_75t_L g5999 ( 
.A(n_5932),
.B(n_5455),
.Y(n_5999)
);

INVxp67_ASAP7_75t_L g6000 ( 
.A(n_5877),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5865),
.Y(n_6001)
);

OR2x2_ASAP7_75t_L g6002 ( 
.A(n_5937),
.B(n_5900),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5945),
.B(n_5897),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5959),
.Y(n_6004)
);

NAND2xp5_ASAP7_75t_L g6005 ( 
.A(n_5968),
.B(n_5922),
.Y(n_6005)
);

AOI22xp5_ASAP7_75t_L g6006 ( 
.A1(n_5951),
.A2(n_5899),
.B1(n_5894),
.B2(n_5912),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5966),
.Y(n_6007)
);

OAI21xp33_ASAP7_75t_L g6008 ( 
.A1(n_5963),
.A2(n_5915),
.B(n_5902),
.Y(n_6008)
);

INVx1_ASAP7_75t_SL g6009 ( 
.A(n_5938),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5972),
.Y(n_6010)
);

AND2x2_ASAP7_75t_L g6011 ( 
.A(n_5983),
.B(n_5985),
.Y(n_6011)
);

NAND2xp5_ASAP7_75t_SL g6012 ( 
.A(n_5964),
.B(n_5895),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5973),
.Y(n_6013)
);

INVx2_ASAP7_75t_L g6014 ( 
.A(n_5985),
.Y(n_6014)
);

HB1xp67_ASAP7_75t_L g6015 ( 
.A(n_5957),
.Y(n_6015)
);

AO21x2_ASAP7_75t_L g6016 ( 
.A1(n_5989),
.A2(n_5886),
.B(n_5905),
.Y(n_6016)
);

INVx2_ASAP7_75t_L g6017 ( 
.A(n_5946),
.Y(n_6017)
);

INVx1_ASAP7_75t_SL g6018 ( 
.A(n_5940),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5970),
.Y(n_6019)
);

INVx3_ASAP7_75t_L g6020 ( 
.A(n_5960),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5980),
.Y(n_6021)
);

AND2x2_ASAP7_75t_L g6022 ( 
.A(n_5939),
.B(n_5888),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5955),
.B(n_5892),
.Y(n_6023)
);

AND2x2_ASAP7_75t_L g6024 ( 
.A(n_5944),
.B(n_5910),
.Y(n_6024)
);

OAI22xp5_ASAP7_75t_L g6025 ( 
.A1(n_5943),
.A2(n_5906),
.B1(n_5933),
.B2(n_5918),
.Y(n_6025)
);

OAI22xp5_ASAP7_75t_L g6026 ( 
.A1(n_5934),
.A2(n_5956),
.B1(n_5976),
.B2(n_6000),
.Y(n_6026)
);

AOI221xp5_ASAP7_75t_SL g6027 ( 
.A1(n_5975),
.A2(n_5909),
.B1(n_5914),
.B2(n_78),
.C(n_76),
.Y(n_6027)
);

AOI22xp33_ASAP7_75t_L g6028 ( 
.A1(n_5986),
.A2(n_5967),
.B1(n_5941),
.B2(n_5936),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_L g6029 ( 
.A(n_5979),
.B(n_5456),
.Y(n_6029)
);

AND2x2_ASAP7_75t_L g6030 ( 
.A(n_5987),
.B(n_5458),
.Y(n_6030)
);

NAND5xp2_ASAP7_75t_L g6031 ( 
.A(n_5942),
.B(n_5993),
.C(n_5971),
.D(n_5977),
.E(n_5949),
.Y(n_6031)
);

OAI221xp5_ASAP7_75t_SL g6032 ( 
.A1(n_5984),
.A2(n_5461),
.B1(n_1035),
.B2(n_1036),
.C(n_1034),
.Y(n_6032)
);

OR2x2_ASAP7_75t_L g6033 ( 
.A(n_5999),
.B(n_76),
.Y(n_6033)
);

INVxp67_ASAP7_75t_SL g6034 ( 
.A(n_5997),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5950),
.Y(n_6035)
);

BUFx3_ASAP7_75t_L g6036 ( 
.A(n_5960),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5952),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_5948),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_5958),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5961),
.Y(n_6040)
);

OAI21xp5_ASAP7_75t_L g6041 ( 
.A1(n_5992),
.A2(n_77),
.B(n_78),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5974),
.Y(n_6042)
);

AND2x2_ASAP7_75t_L g6043 ( 
.A(n_5988),
.B(n_77),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5965),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5935),
.B(n_77),
.Y(n_6045)
);

BUFx3_ASAP7_75t_L g6046 ( 
.A(n_6004),
.Y(n_6046)
);

AND2x2_ASAP7_75t_L g6047 ( 
.A(n_6011),
.B(n_5994),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_6014),
.Y(n_6048)
);

NOR4xp75_ASAP7_75t_L g6049 ( 
.A(n_6026),
.B(n_5995),
.C(n_5996),
.D(n_5998),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_6002),
.Y(n_6050)
);

INVx1_ASAP7_75t_SL g6051 ( 
.A(n_6009),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_6013),
.Y(n_6052)
);

NAND2xp5_ASAP7_75t_L g6053 ( 
.A(n_6034),
.B(n_5991),
.Y(n_6053)
);

NOR2xp67_ASAP7_75t_L g6054 ( 
.A(n_6006),
.B(n_5981),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_6009),
.Y(n_6055)
);

NAND3xp33_ASAP7_75t_L g6056 ( 
.A(n_6028),
.B(n_5947),
.C(n_5982),
.Y(n_6056)
);

AOI22xp33_ASAP7_75t_L g6057 ( 
.A1(n_6018),
.A2(n_5969),
.B1(n_5962),
.B2(n_5990),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_6007),
.Y(n_6058)
);

OR2x2_ASAP7_75t_L g6059 ( 
.A(n_6033),
.B(n_5953),
.Y(n_6059)
);

AND2x2_ASAP7_75t_L g6060 ( 
.A(n_6018),
.B(n_6022),
.Y(n_6060)
);

BUFx2_ASAP7_75t_L g6061 ( 
.A(n_6036),
.Y(n_6061)
);

AOI221xp5_ASAP7_75t_L g6062 ( 
.A1(n_6027),
.A2(n_5962),
.B1(n_6001),
.B2(n_5954),
.C(n_5953),
.Y(n_6062)
);

INVx2_ASAP7_75t_L g6063 ( 
.A(n_6003),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_6010),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_6043),
.Y(n_6065)
);

OR2x2_ASAP7_75t_L g6066 ( 
.A(n_6029),
.B(n_5954),
.Y(n_6066)
);

INVx1_ASAP7_75t_SL g6067 ( 
.A(n_6045),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_6023),
.B(n_5978),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_6024),
.B(n_6001),
.Y(n_6069)
);

NOR2xp33_ASAP7_75t_L g6070 ( 
.A(n_6031),
.B(n_79),
.Y(n_6070)
);

INVx1_ASAP7_75t_L g6071 ( 
.A(n_6019),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_6021),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_6017),
.Y(n_6073)
);

AOI33xp33_ASAP7_75t_L g6074 ( 
.A1(n_6006),
.A2(n_6044),
.A3(n_6030),
.B1(n_6037),
.B2(n_6040),
.B3(n_6039),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_6015),
.Y(n_6075)
);

NAND3xp33_ASAP7_75t_SL g6076 ( 
.A(n_6041),
.B(n_79),
.C(n_80),
.Y(n_6076)
);

INVx2_ASAP7_75t_L g6077 ( 
.A(n_6038),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_6035),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_6042),
.Y(n_6079)
);

AND2x2_ASAP7_75t_L g6080 ( 
.A(n_6020),
.B(n_79),
.Y(n_6080)
);

NAND3x1_ASAP7_75t_L g6081 ( 
.A(n_6005),
.B(n_1036),
.C(n_1033),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_6020),
.B(n_6027),
.Y(n_6082)
);

AOI22xp33_ASAP7_75t_L g6083 ( 
.A1(n_6061),
.A2(n_6008),
.B1(n_6025),
.B2(n_6012),
.Y(n_6083)
);

NAND2xp5_ASAP7_75t_L g6084 ( 
.A(n_6051),
.B(n_6008),
.Y(n_6084)
);

AND2x2_ASAP7_75t_L g6085 ( 
.A(n_6060),
.B(n_6041),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_6082),
.B(n_6016),
.Y(n_6086)
);

AND2x2_ASAP7_75t_L g6087 ( 
.A(n_6055),
.B(n_6016),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_6080),
.Y(n_6088)
);

AND2x2_ASAP7_75t_L g6089 ( 
.A(n_6046),
.B(n_80),
.Y(n_6089)
);

NAND2xp5_ASAP7_75t_L g6090 ( 
.A(n_6051),
.B(n_80),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_6050),
.Y(n_6091)
);

NOR2xp33_ASAP7_75t_L g6092 ( 
.A(n_6056),
.B(n_6032),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_6059),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_6070),
.B(n_80),
.Y(n_6094)
);

NAND2xp5_ASAP7_75t_L g6095 ( 
.A(n_6075),
.B(n_81),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_6048),
.Y(n_6096)
);

NAND2xp5_ASAP7_75t_L g6097 ( 
.A(n_6067),
.B(n_81),
.Y(n_6097)
);

INVx3_ASAP7_75t_SL g6098 ( 
.A(n_6067),
.Y(n_6098)
);

NAND2xp5_ASAP7_75t_L g6099 ( 
.A(n_6062),
.B(n_81),
.Y(n_6099)
);

NAND2xp5_ASAP7_75t_L g6100 ( 
.A(n_6062),
.B(n_81),
.Y(n_6100)
);

INVxp33_ASAP7_75t_L g6101 ( 
.A(n_6053),
.Y(n_6101)
);

HB1xp67_ASAP7_75t_L g6102 ( 
.A(n_6073),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_6052),
.Y(n_6103)
);

OR2x2_ASAP7_75t_L g6104 ( 
.A(n_6053),
.B(n_82),
.Y(n_6104)
);

HB1xp67_ASAP7_75t_L g6105 ( 
.A(n_6077),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_6079),
.Y(n_6106)
);

NAND2xp5_ASAP7_75t_L g6107 ( 
.A(n_6065),
.B(n_82),
.Y(n_6107)
);

AND2x2_ASAP7_75t_L g6108 ( 
.A(n_6069),
.B(n_6047),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_6063),
.B(n_82),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_6058),
.Y(n_6110)
);

OR2x2_ASAP7_75t_L g6111 ( 
.A(n_6076),
.B(n_82),
.Y(n_6111)
);

AND2x2_ASAP7_75t_L g6112 ( 
.A(n_6068),
.B(n_83),
.Y(n_6112)
);

NAND2xp5_ASAP7_75t_L g6113 ( 
.A(n_6064),
.B(n_83),
.Y(n_6113)
);

OR2x2_ASAP7_75t_L g6114 ( 
.A(n_6076),
.B(n_83),
.Y(n_6114)
);

INVx2_ASAP7_75t_L g6115 ( 
.A(n_6066),
.Y(n_6115)
);

INVx1_ASAP7_75t_SL g6116 ( 
.A(n_6081),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_6071),
.Y(n_6117)
);

INVx2_ASAP7_75t_SL g6118 ( 
.A(n_6072),
.Y(n_6118)
);

AND2x2_ASAP7_75t_L g6119 ( 
.A(n_6057),
.B(n_83),
.Y(n_6119)
);

AND2x2_ASAP7_75t_L g6120 ( 
.A(n_6054),
.B(n_84),
.Y(n_6120)
);

AND2x2_ASAP7_75t_L g6121 ( 
.A(n_6054),
.B(n_84),
.Y(n_6121)
);

NAND2xp5_ASAP7_75t_L g6122 ( 
.A(n_6056),
.B(n_84),
.Y(n_6122)
);

OR2x2_ASAP7_75t_L g6123 ( 
.A(n_6078),
.B(n_85),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_6090),
.Y(n_6124)
);

NAND2x2_ASAP7_75t_L g6125 ( 
.A(n_6099),
.B(n_6049),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_6089),
.Y(n_6126)
);

OAI32xp33_ASAP7_75t_L g6127 ( 
.A1(n_6101),
.A2(n_6074),
.A3(n_88),
.B1(n_85),
.B2(n_87),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_6102),
.Y(n_6128)
);

OR2x2_ASAP7_75t_L g6129 ( 
.A(n_6098),
.B(n_87),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_6105),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_6111),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_6114),
.Y(n_6132)
);

HB1xp67_ASAP7_75t_L g6133 ( 
.A(n_6096),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_6109),
.Y(n_6134)
);

INVx2_ASAP7_75t_L g6135 ( 
.A(n_6106),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_6085),
.B(n_87),
.Y(n_6136)
);

INVx1_ASAP7_75t_SL g6137 ( 
.A(n_6091),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_6119),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_6097),
.Y(n_6139)
);

NOR2xp33_ASAP7_75t_L g6140 ( 
.A(n_6116),
.B(n_87),
.Y(n_6140)
);

NAND2xp5_ASAP7_75t_L g6141 ( 
.A(n_6120),
.B(n_6121),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_6112),
.Y(n_6142)
);

OAI22xp33_ASAP7_75t_L g6143 ( 
.A1(n_6100),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_6108),
.B(n_88),
.Y(n_6144)
);

OR2x2_ASAP7_75t_L g6145 ( 
.A(n_6104),
.B(n_89),
.Y(n_6145)
);

INVxp67_ASAP7_75t_L g6146 ( 
.A(n_6084),
.Y(n_6146)
);

NAND2xp5_ASAP7_75t_L g6147 ( 
.A(n_6086),
.B(n_89),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_6087),
.Y(n_6148)
);

OAI21xp33_ASAP7_75t_SL g6149 ( 
.A1(n_6083),
.A2(n_89),
.B(n_90),
.Y(n_6149)
);

INVx2_ASAP7_75t_L g6150 ( 
.A(n_6115),
.Y(n_6150)
);

OAI22xp5_ASAP7_75t_L g6151 ( 
.A1(n_6092),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_6088),
.Y(n_6152)
);

NAND2xp5_ASAP7_75t_SL g6153 ( 
.A(n_6084),
.B(n_91),
.Y(n_6153)
);

INVx3_ASAP7_75t_L g6154 ( 
.A(n_6123),
.Y(n_6154)
);

NOR2xp33_ASAP7_75t_SL g6155 ( 
.A(n_6116),
.B(n_92),
.Y(n_6155)
);

AND2x2_ASAP7_75t_L g6156 ( 
.A(n_6093),
.B(n_92),
.Y(n_6156)
);

AOI22xp5_ASAP7_75t_L g6157 ( 
.A1(n_6122),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_6118),
.Y(n_6158)
);

AOI22xp5_ASAP7_75t_L g6159 ( 
.A1(n_6094),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_6159)
);

AND2x2_ASAP7_75t_L g6160 ( 
.A(n_6107),
.B(n_93),
.Y(n_6160)
);

NAND2xp5_ASAP7_75t_L g6161 ( 
.A(n_6095),
.B(n_94),
.Y(n_6161)
);

NAND2xp5_ASAP7_75t_L g6162 ( 
.A(n_6095),
.B(n_94),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_6107),
.Y(n_6163)
);

AOI22xp5_ASAP7_75t_L g6164 ( 
.A1(n_6149),
.A2(n_6113),
.B1(n_6103),
.B2(n_6110),
.Y(n_6164)
);

INVxp67_ASAP7_75t_L g6165 ( 
.A(n_6155),
.Y(n_6165)
);

AOI322xp5_ASAP7_75t_L g6166 ( 
.A1(n_6131),
.A2(n_6117),
.A3(n_6113),
.B1(n_97),
.B2(n_98),
.C1(n_99),
.C2(n_100),
.Y(n_6166)
);

NOR2xp33_ASAP7_75t_L g6167 ( 
.A(n_6127),
.B(n_6146),
.Y(n_6167)
);

AND2x2_ASAP7_75t_L g6168 ( 
.A(n_6144),
.B(n_95),
.Y(n_6168)
);

AND2x2_ASAP7_75t_L g6169 ( 
.A(n_6156),
.B(n_95),
.Y(n_6169)
);

O2A1O1Ixp33_ASAP7_75t_SL g6170 ( 
.A1(n_6153),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_6133),
.Y(n_6171)
);

OAI322xp33_ASAP7_75t_L g6172 ( 
.A1(n_6128),
.A2(n_96),
.A3(n_97),
.B1(n_98),
.B2(n_99),
.C1(n_100),
.C2(n_101),
.Y(n_6172)
);

INVx1_ASAP7_75t_SL g6173 ( 
.A(n_6137),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_6130),
.Y(n_6174)
);

INVx1_ASAP7_75t_SL g6175 ( 
.A(n_6135),
.Y(n_6175)
);

OAI311xp33_ASAP7_75t_L g6176 ( 
.A1(n_6148),
.A2(n_98),
.A3(n_96),
.B1(n_97),
.C1(n_99),
.Y(n_6176)
);

OR2x6_ASAP7_75t_L g6177 ( 
.A(n_6158),
.B(n_1036),
.Y(n_6177)
);

OAI21xp5_ASAP7_75t_L g6178 ( 
.A1(n_6140),
.A2(n_96),
.B(n_99),
.Y(n_6178)
);

OAI21xp5_ASAP7_75t_SL g6179 ( 
.A1(n_6147),
.A2(n_100),
.B(n_101),
.Y(n_6179)
);

NOR2xp33_ASAP7_75t_SL g6180 ( 
.A(n_6132),
.B(n_101),
.Y(n_6180)
);

INVx1_ASAP7_75t_L g6181 ( 
.A(n_6160),
.Y(n_6181)
);

OAI21xp33_ASAP7_75t_L g6182 ( 
.A1(n_6138),
.A2(n_101),
.B(n_102),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_6145),
.Y(n_6183)
);

AND2x2_ASAP7_75t_L g6184 ( 
.A(n_6142),
.B(n_102),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_6126),
.Y(n_6185)
);

XNOR2x1_ASAP7_75t_L g6186 ( 
.A(n_6151),
.B(n_102),
.Y(n_6186)
);

O2A1O1Ixp5_ASAP7_75t_SL g6187 ( 
.A1(n_6152),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_6187)
);

NAND4xp25_ASAP7_75t_SL g6188 ( 
.A(n_6141),
.B(n_105),
.C(n_103),
.D(n_104),
.Y(n_6188)
);

OAI22xp5_ASAP7_75t_L g6189 ( 
.A1(n_6125),
.A2(n_6136),
.B1(n_6134),
.B2(n_6124),
.Y(n_6189)
);

INVx2_ASAP7_75t_L g6190 ( 
.A(n_6154),
.Y(n_6190)
);

HB1xp67_ASAP7_75t_L g6191 ( 
.A(n_6154),
.Y(n_6191)
);

AOI221x1_ASAP7_75t_L g6192 ( 
.A1(n_6124),
.A2(n_106),
.B1(n_103),
.B2(n_105),
.C(n_107),
.Y(n_6192)
);

OAI21xp5_ASAP7_75t_L g6193 ( 
.A1(n_6163),
.A2(n_103),
.B(n_105),
.Y(n_6193)
);

CKINVDCx16_ASAP7_75t_R g6194 ( 
.A(n_6159),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_6161),
.Y(n_6195)
);

OAI22xp33_ASAP7_75t_L g6196 ( 
.A1(n_6157),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_6162),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_6139),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_6143),
.Y(n_6199)
);

NAND2xp5_ASAP7_75t_L g6200 ( 
.A(n_6155),
.B(n_106),
.Y(n_6200)
);

XNOR2xp5_ASAP7_75t_L g6201 ( 
.A(n_6144),
.B(n_106),
.Y(n_6201)
);

OAI21xp5_ASAP7_75t_L g6202 ( 
.A1(n_6149),
.A2(n_107),
.B(n_108),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_6144),
.B(n_108),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_6129),
.Y(n_6204)
);

NOR2xp33_ASAP7_75t_L g6205 ( 
.A(n_6149),
.B(n_109),
.Y(n_6205)
);

AOI321xp33_ASAP7_75t_L g6206 ( 
.A1(n_6127),
.A2(n_109),
.A3(n_110),
.B1(n_111),
.B2(n_112),
.C(n_113),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_6155),
.B(n_109),
.Y(n_6207)
);

NOR2xp33_ASAP7_75t_SL g6208 ( 
.A(n_6137),
.B(n_110),
.Y(n_6208)
);

A2O1A1Ixp33_ASAP7_75t_L g6209 ( 
.A1(n_6149),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_6209)
);

INVx2_ASAP7_75t_L g6210 ( 
.A(n_6150),
.Y(n_6210)
);

INVx1_ASAP7_75t_L g6211 ( 
.A(n_6129),
.Y(n_6211)
);

AND2x2_ASAP7_75t_L g6212 ( 
.A(n_6144),
.B(n_111),
.Y(n_6212)
);

OAI22xp5_ASAP7_75t_L g6213 ( 
.A1(n_6125),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_6213)
);

INVx1_ASAP7_75t_SL g6214 ( 
.A(n_6173),
.Y(n_6214)
);

OAI21xp5_ASAP7_75t_L g6215 ( 
.A1(n_6205),
.A2(n_114),
.B(n_115),
.Y(n_6215)
);

OAI21xp5_ASAP7_75t_L g6216 ( 
.A1(n_6209),
.A2(n_114),
.B(n_115),
.Y(n_6216)
);

AOI21xp5_ASAP7_75t_L g6217 ( 
.A1(n_6200),
.A2(n_115),
.B(n_116),
.Y(n_6217)
);

OAI21xp5_ASAP7_75t_SL g6218 ( 
.A1(n_6213),
.A2(n_115),
.B(n_116),
.Y(n_6218)
);

INVx2_ASAP7_75t_L g6219 ( 
.A(n_6210),
.Y(n_6219)
);

AOI22xp5_ASAP7_75t_L g6220 ( 
.A1(n_6165),
.A2(n_6199),
.B1(n_6167),
.B2(n_6208),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_L g6221 ( 
.A(n_6169),
.B(n_116),
.Y(n_6221)
);

OAI32xp33_ASAP7_75t_L g6222 ( 
.A1(n_6175),
.A2(n_118),
.A3(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_6222)
);

OAI31xp33_ASAP7_75t_L g6223 ( 
.A1(n_6176),
.A2(n_119),
.A3(n_117),
.B(n_118),
.Y(n_6223)
);

INVx3_ASAP7_75t_L g6224 ( 
.A(n_6190),
.Y(n_6224)
);

AOI22xp5_ASAP7_75t_L g6225 ( 
.A1(n_6188),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_6225)
);

NAND2xp5_ASAP7_75t_L g6226 ( 
.A(n_6168),
.B(n_120),
.Y(n_6226)
);

AOI32xp33_ASAP7_75t_L g6227 ( 
.A1(n_6171),
.A2(n_122),
.A3(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_6227)
);

A2O1A1Ixp33_ASAP7_75t_L g6228 ( 
.A1(n_6182),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_6228)
);

NAND2xp5_ASAP7_75t_L g6229 ( 
.A(n_6203),
.B(n_120),
.Y(n_6229)
);

AOI211x1_ASAP7_75t_L g6230 ( 
.A1(n_6189),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_6230)
);

AOI21xp33_ASAP7_75t_L g6231 ( 
.A1(n_6191),
.A2(n_121),
.B(n_122),
.Y(n_6231)
);

OAI21xp5_ASAP7_75t_L g6232 ( 
.A1(n_6166),
.A2(n_123),
.B(n_124),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_6207),
.Y(n_6233)
);

OAI21xp33_ASAP7_75t_L g6234 ( 
.A1(n_6180),
.A2(n_123),
.B(n_124),
.Y(n_6234)
);

NAND2xp5_ASAP7_75t_L g6235 ( 
.A(n_6212),
.B(n_124),
.Y(n_6235)
);

AOI21xp33_ASAP7_75t_SL g6236 ( 
.A1(n_6186),
.A2(n_6201),
.B(n_6194),
.Y(n_6236)
);

AOI222xp33_ASAP7_75t_L g6237 ( 
.A1(n_6174),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.C1(n_127),
.C2(n_128),
.Y(n_6237)
);

NOR3xp33_ASAP7_75t_L g6238 ( 
.A(n_6172),
.B(n_125),
.C(n_126),
.Y(n_6238)
);

OAI31xp33_ASAP7_75t_L g6239 ( 
.A1(n_6179),
.A2(n_127),
.A3(n_125),
.B(n_126),
.Y(n_6239)
);

INVx1_ASAP7_75t_L g6240 ( 
.A(n_6177),
.Y(n_6240)
);

AOI222xp33_ASAP7_75t_L g6241 ( 
.A1(n_6204),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.C1(n_129),
.C2(n_130),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_6177),
.Y(n_6242)
);

OAI21xp5_ASAP7_75t_L g6243 ( 
.A1(n_6164),
.A2(n_128),
.B(n_129),
.Y(n_6243)
);

AOI21xp33_ASAP7_75t_SL g6244 ( 
.A1(n_6196),
.A2(n_129),
.B(n_130),
.Y(n_6244)
);

OAI21xp5_ASAP7_75t_L g6245 ( 
.A1(n_6211),
.A2(n_130),
.B(n_131),
.Y(n_6245)
);

INVx1_ASAP7_75t_SL g6246 ( 
.A(n_6184),
.Y(n_6246)
);

INVxp67_ASAP7_75t_L g6247 ( 
.A(n_6202),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_6183),
.Y(n_6248)
);

OAI21xp33_ASAP7_75t_L g6249 ( 
.A1(n_6181),
.A2(n_130),
.B(n_131),
.Y(n_6249)
);

HB1xp67_ASAP7_75t_L g6250 ( 
.A(n_6185),
.Y(n_6250)
);

OAI22xp33_ASAP7_75t_L g6251 ( 
.A1(n_6192),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_6251)
);

AOI31xp33_ASAP7_75t_L g6252 ( 
.A1(n_6178),
.A2(n_134),
.A3(n_132),
.B(n_133),
.Y(n_6252)
);

AND2x2_ASAP7_75t_L g6253 ( 
.A(n_6195),
.B(n_132),
.Y(n_6253)
);

OAI21xp5_ASAP7_75t_L g6254 ( 
.A1(n_6215),
.A2(n_6193),
.B(n_6187),
.Y(n_6254)
);

OA22x2_ASAP7_75t_L g6255 ( 
.A1(n_6220),
.A2(n_6197),
.B1(n_6198),
.B2(n_6206),
.Y(n_6255)
);

AOI221xp5_ASAP7_75t_L g6256 ( 
.A1(n_6251),
.A2(n_6170),
.B1(n_134),
.B2(n_132),
.C(n_133),
.Y(n_6256)
);

INVx1_ASAP7_75t_L g6257 ( 
.A(n_6224),
.Y(n_6257)
);

AOI21xp5_ASAP7_75t_L g6258 ( 
.A1(n_6223),
.A2(n_133),
.B(n_134),
.Y(n_6258)
);

AOI322xp5_ASAP7_75t_L g6259 ( 
.A1(n_6214),
.A2(n_135),
.A3(n_136),
.B1(n_137),
.B2(n_138),
.C1(n_139),
.C2(n_140),
.Y(n_6259)
);

A2O1A1Ixp33_ASAP7_75t_L g6260 ( 
.A1(n_6227),
.A2(n_6239),
.B(n_6234),
.C(n_6249),
.Y(n_6260)
);

AND5x1_ASAP7_75t_L g6261 ( 
.A(n_6217),
.B(n_137),
.C(n_135),
.D(n_136),
.E(n_138),
.Y(n_6261)
);

OAI21xp33_ASAP7_75t_L g6262 ( 
.A1(n_6218),
.A2(n_136),
.B(n_138),
.Y(n_6262)
);

OAI21xp5_ASAP7_75t_L g6263 ( 
.A1(n_6247),
.A2(n_136),
.B(n_139),
.Y(n_6263)
);

AOI21xp5_ASAP7_75t_L g6264 ( 
.A1(n_6221),
.A2(n_139),
.B(n_140),
.Y(n_6264)
);

OAI21xp33_ASAP7_75t_SL g6265 ( 
.A1(n_6243),
.A2(n_6246),
.B(n_6219),
.Y(n_6265)
);

OAI21xp5_ASAP7_75t_L g6266 ( 
.A1(n_6236),
.A2(n_139),
.B(n_140),
.Y(n_6266)
);

NAND2xp5_ASAP7_75t_L g6267 ( 
.A(n_6238),
.B(n_141),
.Y(n_6267)
);

AOI21xp5_ASAP7_75t_L g6268 ( 
.A1(n_6226),
.A2(n_141),
.B(n_142),
.Y(n_6268)
);

OAI221xp5_ASAP7_75t_SL g6269 ( 
.A1(n_6240),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_6269)
);

OAI321xp33_ASAP7_75t_L g6270 ( 
.A1(n_6248),
.A2(n_142),
.A3(n_143),
.B1(n_144),
.B2(n_145),
.C(n_146),
.Y(n_6270)
);

AOI222xp33_ASAP7_75t_L g6271 ( 
.A1(n_6224),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.C1(n_145),
.C2(n_146),
.Y(n_6271)
);

AOI221xp5_ASAP7_75t_L g6272 ( 
.A1(n_6230),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.C(n_147),
.Y(n_6272)
);

NOR3xp33_ASAP7_75t_L g6273 ( 
.A(n_6232),
.B(n_145),
.C(n_147),
.Y(n_6273)
);

AOI211xp5_ASAP7_75t_L g6274 ( 
.A1(n_6244),
.A2(n_6231),
.B(n_6245),
.C(n_6222),
.Y(n_6274)
);

NOR3xp33_ASAP7_75t_L g6275 ( 
.A(n_6216),
.B(n_6252),
.C(n_6228),
.Y(n_6275)
);

AOI211x1_ASAP7_75t_SL g6276 ( 
.A1(n_6242),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_6276)
);

NOR2xp33_ASAP7_75t_L g6277 ( 
.A(n_6229),
.B(n_147),
.Y(n_6277)
);

OAI21xp33_ASAP7_75t_L g6278 ( 
.A1(n_6253),
.A2(n_148),
.B(n_149),
.Y(n_6278)
);

AOI22xp33_ASAP7_75t_SL g6279 ( 
.A1(n_6250),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_6279)
);

OAI21xp33_ASAP7_75t_L g6280 ( 
.A1(n_6233),
.A2(n_150),
.B(n_151),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_6225),
.B(n_153),
.Y(n_6281)
);

AOI22xp5_ASAP7_75t_L g6282 ( 
.A1(n_6235),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_6282)
);

NAND2xp5_ASAP7_75t_L g6283 ( 
.A(n_6241),
.B(n_154),
.Y(n_6283)
);

AOI21xp33_ASAP7_75t_L g6284 ( 
.A1(n_6237),
.A2(n_156),
.B(n_157),
.Y(n_6284)
);

NAND3xp33_ASAP7_75t_L g6285 ( 
.A(n_6241),
.B(n_156),
.C(n_157),
.Y(n_6285)
);

OAI221xp5_ASAP7_75t_L g6286 ( 
.A1(n_6223),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.C(n_159),
.Y(n_6286)
);

AOI221x1_ASAP7_75t_L g6287 ( 
.A1(n_6236),
.A2(n_159),
.B1(n_156),
.B2(n_158),
.C(n_160),
.Y(n_6287)
);

AND2x2_ASAP7_75t_L g6288 ( 
.A(n_6214),
.B(n_158),
.Y(n_6288)
);

O2A1O1Ixp33_ASAP7_75t_L g6289 ( 
.A1(n_6231),
.A2(n_161),
.B(n_158),
.C(n_160),
.Y(n_6289)
);

NOR3xp33_ASAP7_75t_L g6290 ( 
.A(n_6232),
.B(n_160),
.C(n_161),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_6224),
.Y(n_6291)
);

NAND2xp5_ASAP7_75t_L g6292 ( 
.A(n_6214),
.B(n_160),
.Y(n_6292)
);

INVx2_ASAP7_75t_L g6293 ( 
.A(n_6224),
.Y(n_6293)
);

AO22x1_ASAP7_75t_L g6294 ( 
.A1(n_6238),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_6294)
);

AOI211xp5_ASAP7_75t_L g6295 ( 
.A1(n_6236),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_6295)
);

NAND2xp5_ASAP7_75t_L g6296 ( 
.A(n_6294),
.B(n_6258),
.Y(n_6296)
);

AOI21xp5_ASAP7_75t_L g6297 ( 
.A1(n_6286),
.A2(n_162),
.B(n_163),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_6288),
.Y(n_6298)
);

O2A1O1Ixp33_ASAP7_75t_L g6299 ( 
.A1(n_6284),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_6299)
);

OAI21xp33_ASAP7_75t_L g6300 ( 
.A1(n_6267),
.A2(n_164),
.B(n_165),
.Y(n_6300)
);

AOI221xp5_ASAP7_75t_L g6301 ( 
.A1(n_6289),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.C(n_167),
.Y(n_6301)
);

AOI322xp5_ASAP7_75t_L g6302 ( 
.A1(n_6265),
.A2(n_165),
.A3(n_166),
.B1(n_167),
.B2(n_168),
.C1(n_169),
.C2(n_170),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_6277),
.B(n_166),
.Y(n_6303)
);

NAND2xp5_ASAP7_75t_L g6304 ( 
.A(n_6259),
.B(n_6276),
.Y(n_6304)
);

OAI21xp5_ASAP7_75t_SL g6305 ( 
.A1(n_6256),
.A2(n_166),
.B(n_167),
.Y(n_6305)
);

NOR4xp25_ASAP7_75t_L g6306 ( 
.A(n_6257),
.B(n_169),
.C(n_167),
.D(n_168),
.Y(n_6306)
);

AOI21xp5_ASAP7_75t_L g6307 ( 
.A1(n_6281),
.A2(n_168),
.B(n_169),
.Y(n_6307)
);

NOR2xp33_ASAP7_75t_SL g6308 ( 
.A(n_6293),
.B(n_168),
.Y(n_6308)
);

OR2x2_ASAP7_75t_L g6309 ( 
.A(n_6292),
.B(n_170),
.Y(n_6309)
);

AOI221xp5_ASAP7_75t_L g6310 ( 
.A1(n_6272),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.C(n_173),
.Y(n_6310)
);

A2O1A1Ixp33_ASAP7_75t_L g6311 ( 
.A1(n_6262),
.A2(n_6280),
.B(n_6285),
.C(n_6278),
.Y(n_6311)
);

OAI222xp33_ASAP7_75t_L g6312 ( 
.A1(n_6255),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.C1(n_173),
.C2(n_174),
.Y(n_6312)
);

AOI221xp5_ASAP7_75t_L g6313 ( 
.A1(n_6270),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.C(n_174),
.Y(n_6313)
);

AOI221xp5_ASAP7_75t_L g6314 ( 
.A1(n_6273),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.C(n_175),
.Y(n_6314)
);

O2A1O1Ixp33_ASAP7_75t_L g6315 ( 
.A1(n_6269),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_6315)
);

AOI22xp5_ASAP7_75t_L g6316 ( 
.A1(n_6290),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_6316)
);

INVx1_ASAP7_75t_SL g6317 ( 
.A(n_6291),
.Y(n_6317)
);

OAI32xp33_ASAP7_75t_L g6318 ( 
.A1(n_6283),
.A2(n_175),
.A3(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_6318)
);

AOI21xp5_ASAP7_75t_L g6319 ( 
.A1(n_6260),
.A2(n_176),
.B(n_177),
.Y(n_6319)
);

NAND2xp5_ASAP7_75t_SL g6320 ( 
.A(n_6295),
.B(n_177),
.Y(n_6320)
);

AOI22xp33_ASAP7_75t_L g6321 ( 
.A1(n_6275),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_6321)
);

NAND2xp5_ASAP7_75t_L g6322 ( 
.A(n_6279),
.B(n_178),
.Y(n_6322)
);

AOI22xp33_ASAP7_75t_L g6323 ( 
.A1(n_6266),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_6323)
);

INVxp67_ASAP7_75t_SL g6324 ( 
.A(n_6271),
.Y(n_6324)
);

OAI22xp5_ASAP7_75t_SL g6325 ( 
.A1(n_6274),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_6325)
);

AOI22xp5_ASAP7_75t_L g6326 ( 
.A1(n_6282),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_6326)
);

AOI22xp5_ASAP7_75t_L g6327 ( 
.A1(n_6264),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_6327)
);

AOI22xp33_ASAP7_75t_L g6328 ( 
.A1(n_6268),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_6328)
);

AOI21xp5_ASAP7_75t_L g6329 ( 
.A1(n_6263),
.A2(n_182),
.B(n_183),
.Y(n_6329)
);

INVx1_ASAP7_75t_L g6330 ( 
.A(n_6287),
.Y(n_6330)
);

AOI21xp5_ASAP7_75t_L g6331 ( 
.A1(n_6254),
.A2(n_182),
.B(n_183),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_6261),
.B(n_184),
.Y(n_6332)
);

OAI221xp5_ASAP7_75t_L g6333 ( 
.A1(n_6286),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_6333)
);

AO21x1_ASAP7_75t_L g6334 ( 
.A1(n_6283),
.A2(n_184),
.B(n_185),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_6332),
.Y(n_6335)
);

XOR2xp5_ASAP7_75t_L g6336 ( 
.A(n_6325),
.B(n_185),
.Y(n_6336)
);

OAI21xp5_ASAP7_75t_L g6337 ( 
.A1(n_6319),
.A2(n_186),
.B(n_187),
.Y(n_6337)
);

BUFx2_ASAP7_75t_L g6338 ( 
.A(n_6330),
.Y(n_6338)
);

AOI22xp5_ASAP7_75t_L g6339 ( 
.A1(n_6324),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_6339)
);

AOI22xp5_ASAP7_75t_L g6340 ( 
.A1(n_6317),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6309),
.Y(n_6341)
);

OAI22xp5_ASAP7_75t_L g6342 ( 
.A1(n_6322),
.A2(n_6304),
.B1(n_6321),
.B2(n_6296),
.Y(n_6342)
);

AOI32xp33_ASAP7_75t_L g6343 ( 
.A1(n_6313),
.A2(n_189),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_6343)
);

OAI311xp33_ASAP7_75t_L g6344 ( 
.A1(n_6305),
.A2(n_189),
.A3(n_190),
.B1(n_191),
.C1(n_192),
.Y(n_6344)
);

AOI221xp5_ASAP7_75t_L g6345 ( 
.A1(n_6306),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_6345)
);

INVx1_ASAP7_75t_L g6346 ( 
.A(n_6334),
.Y(n_6346)
);

O2A1O1Ixp33_ASAP7_75t_L g6347 ( 
.A1(n_6312),
.A2(n_6320),
.B(n_6311),
.C(n_6318),
.Y(n_6347)
);

OAI22xp5_ASAP7_75t_L g6348 ( 
.A1(n_6328),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_6348)
);

AOI211xp5_ASAP7_75t_L g6349 ( 
.A1(n_6333),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_6349)
);

XNOR2xp5_ASAP7_75t_L g6350 ( 
.A(n_6303),
.B(n_193),
.Y(n_6350)
);

AOI21xp5_ASAP7_75t_L g6351 ( 
.A1(n_6315),
.A2(n_194),
.B(n_195),
.Y(n_6351)
);

NAND2xp33_ASAP7_75t_SL g6352 ( 
.A(n_6298),
.B(n_195),
.Y(n_6352)
);

AOI21xp5_ASAP7_75t_L g6353 ( 
.A1(n_6297),
.A2(n_196),
.B(n_197),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_SL g6354 ( 
.A(n_6302),
.B(n_196),
.Y(n_6354)
);

O2A1O1Ixp33_ASAP7_75t_L g6355 ( 
.A1(n_6299),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_6355)
);

O2A1O1Ixp5_ASAP7_75t_L g6356 ( 
.A1(n_6331),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_6356)
);

INVx2_ASAP7_75t_SL g6357 ( 
.A(n_6327),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_6308),
.Y(n_6358)
);

OAI22xp5_ASAP7_75t_L g6359 ( 
.A1(n_6323),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_6359)
);

AOI21xp33_ASAP7_75t_L g6360 ( 
.A1(n_6300),
.A2(n_199),
.B(n_200),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_6316),
.Y(n_6361)
);

OAI211xp5_ASAP7_75t_L g6362 ( 
.A1(n_6310),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_6362)
);

NOR2xp33_ASAP7_75t_L g6363 ( 
.A(n_6307),
.B(n_199),
.Y(n_6363)
);

AOI221xp5_ASAP7_75t_L g6364 ( 
.A1(n_6301),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_6364)
);

AOI221xp5_ASAP7_75t_L g6365 ( 
.A1(n_6314),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_6326),
.Y(n_6366)
);

INVx2_ASAP7_75t_L g6367 ( 
.A(n_6329),
.Y(n_6367)
);

AOI221xp5_ASAP7_75t_L g6368 ( 
.A1(n_6360),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.C(n_205),
.Y(n_6368)
);

HB1xp67_ASAP7_75t_L g6369 ( 
.A(n_6338),
.Y(n_6369)
);

NAND4xp25_ASAP7_75t_L g6370 ( 
.A(n_6339),
.B(n_206),
.C(n_202),
.D(n_205),
.Y(n_6370)
);

OAI22xp5_ASAP7_75t_L g6371 ( 
.A1(n_6336),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_6371)
);

OAI21xp33_ASAP7_75t_L g6372 ( 
.A1(n_6335),
.A2(n_206),
.B(n_207),
.Y(n_6372)
);

CKINVDCx20_ASAP7_75t_R g6373 ( 
.A(n_6350),
.Y(n_6373)
);

AND2x2_ASAP7_75t_L g6374 ( 
.A(n_6363),
.B(n_206),
.Y(n_6374)
);

OAI221xp5_ASAP7_75t_L g6375 ( 
.A1(n_6343),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.C(n_210),
.Y(n_6375)
);

OAI21xp5_ASAP7_75t_L g6376 ( 
.A1(n_6351),
.A2(n_6356),
.B(n_6353),
.Y(n_6376)
);

AND2x4_ASAP7_75t_L g6377 ( 
.A(n_6358),
.B(n_207),
.Y(n_6377)
);

NOR2x1_ASAP7_75t_L g6378 ( 
.A(n_6354),
.B(n_208),
.Y(n_6378)
);

NAND2xp5_ASAP7_75t_L g6379 ( 
.A(n_6345),
.B(n_208),
.Y(n_6379)
);

OAI31xp33_ASAP7_75t_L g6380 ( 
.A1(n_6362),
.A2(n_210),
.A3(n_208),
.B(n_209),
.Y(n_6380)
);

OAI21xp5_ASAP7_75t_L g6381 ( 
.A1(n_6355),
.A2(n_209),
.B(n_210),
.Y(n_6381)
);

NAND3xp33_ASAP7_75t_L g6382 ( 
.A(n_6364),
.B(n_209),
.C(n_211),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_6367),
.Y(n_6383)
);

AOI22xp5_ASAP7_75t_L g6384 ( 
.A1(n_6342),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_6384)
);

NAND4xp25_ASAP7_75t_SL g6385 ( 
.A(n_6347),
.B(n_214),
.C(n_212),
.D(n_213),
.Y(n_6385)
);

AND3x4_ASAP7_75t_L g6386 ( 
.A(n_6344),
.B(n_212),
.C(n_213),
.Y(n_6386)
);

AOI22xp5_ASAP7_75t_L g6387 ( 
.A1(n_6357),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_6387)
);

OAI22xp33_ASAP7_75t_L g6388 ( 
.A1(n_6340),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_6388)
);

AOI211xp5_ASAP7_75t_L g6389 ( 
.A1(n_6359),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_6389)
);

NAND2xp5_ASAP7_75t_L g6390 ( 
.A(n_6377),
.B(n_6346),
.Y(n_6390)
);

AOI22xp5_ASAP7_75t_L g6391 ( 
.A1(n_6386),
.A2(n_6361),
.B1(n_6366),
.B2(n_6352),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_6383),
.Y(n_6392)
);

AOI221xp5_ASAP7_75t_L g6393 ( 
.A1(n_6385),
.A2(n_6348),
.B1(n_6365),
.B2(n_6337),
.C(n_6349),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_6369),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_6378),
.Y(n_6395)
);

OAI31xp33_ASAP7_75t_L g6396 ( 
.A1(n_6388),
.A2(n_6341),
.A3(n_217),
.B(n_215),
.Y(n_6396)
);

NOR2x1_ASAP7_75t_L g6397 ( 
.A(n_6382),
.B(n_215),
.Y(n_6397)
);

AOI22xp33_ASAP7_75t_SL g6398 ( 
.A1(n_6371),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_6398)
);

NOR4xp25_ASAP7_75t_L g6399 ( 
.A(n_6372),
.B(n_6375),
.C(n_6379),
.D(n_6370),
.Y(n_6399)
);

OR2x2_ASAP7_75t_L g6400 ( 
.A(n_6381),
.B(n_216),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_6387),
.Y(n_6401)
);

OR2x2_ASAP7_75t_L g6402 ( 
.A(n_6384),
.B(n_217),
.Y(n_6402)
);

INVxp67_ASAP7_75t_L g6403 ( 
.A(n_6374),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_L g6404 ( 
.A(n_6380),
.B(n_218),
.Y(n_6404)
);

AND2x2_ASAP7_75t_L g6405 ( 
.A(n_6376),
.B(n_218),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6373),
.Y(n_6406)
);

INVx2_ASAP7_75t_SL g6407 ( 
.A(n_6389),
.Y(n_6407)
);

NOR2x1_ASAP7_75t_L g6408 ( 
.A(n_6368),
.B(n_218),
.Y(n_6408)
);

NOR2x1_ASAP7_75t_L g6409 ( 
.A(n_6385),
.B(n_219),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6377),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_6404),
.Y(n_6411)
);

NAND4xp75_ASAP7_75t_L g6412 ( 
.A(n_6397),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_6392),
.Y(n_6413)
);

AO22x2_ASAP7_75t_L g6414 ( 
.A1(n_6394),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_6409),
.Y(n_6415)
);

XNOR2xp5_ASAP7_75t_L g6416 ( 
.A(n_6391),
.B(n_219),
.Y(n_6416)
);

XOR2xp5_ASAP7_75t_L g6417 ( 
.A(n_6406),
.B(n_220),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_6410),
.Y(n_6418)
);

INVx2_ASAP7_75t_L g6419 ( 
.A(n_6390),
.Y(n_6419)
);

AO22x2_ASAP7_75t_L g6420 ( 
.A1(n_6405),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_6420)
);

XNOR2xp5_ASAP7_75t_L g6421 ( 
.A(n_6399),
.B(n_222),
.Y(n_6421)
);

INVx2_ASAP7_75t_L g6422 ( 
.A(n_6407),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_6408),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6400),
.Y(n_6424)
);

NOR2xp67_ASAP7_75t_L g6425 ( 
.A(n_6403),
.B(n_222),
.Y(n_6425)
);

INVx2_ASAP7_75t_L g6426 ( 
.A(n_6402),
.Y(n_6426)
);

OR2x2_ASAP7_75t_L g6427 ( 
.A(n_6401),
.B(n_223),
.Y(n_6427)
);

AOI221xp5_ASAP7_75t_L g6428 ( 
.A1(n_6413),
.A2(n_6393),
.B1(n_6398),
.B2(n_6396),
.C(n_6395),
.Y(n_6428)
);

AOI22xp5_ASAP7_75t_L g6429 ( 
.A1(n_6421),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_6429)
);

NOR2x1_ASAP7_75t_L g6430 ( 
.A(n_6427),
.B(n_223),
.Y(n_6430)
);

NOR3xp33_ASAP7_75t_L g6431 ( 
.A(n_6419),
.B(n_224),
.C(n_225),
.Y(n_6431)
);

AND2x2_ASAP7_75t_L g6432 ( 
.A(n_6418),
.B(n_224),
.Y(n_6432)
);

AND2x4_ASAP7_75t_L g6433 ( 
.A(n_6422),
.B(n_224),
.Y(n_6433)
);

AND2x4_ASAP7_75t_L g6434 ( 
.A(n_6426),
.B(n_225),
.Y(n_6434)
);

AOI221xp5_ASAP7_75t_L g6435 ( 
.A1(n_6414),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.C(n_229),
.Y(n_6435)
);

OAI211xp5_ASAP7_75t_SL g6436 ( 
.A1(n_6411),
.A2(n_226),
.B(n_227),
.C(n_228),
.Y(n_6436)
);

XNOR2x1_ASAP7_75t_L g6437 ( 
.A(n_6430),
.B(n_6416),
.Y(n_6437)
);

INVxp67_ASAP7_75t_L g6438 ( 
.A(n_6432),
.Y(n_6438)
);

AND2x2_ASAP7_75t_SL g6439 ( 
.A(n_6431),
.B(n_6415),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6433),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6434),
.Y(n_6441)
);

INVx3_ASAP7_75t_L g6442 ( 
.A(n_6428),
.Y(n_6442)
);

NOR2xp67_ASAP7_75t_L g6443 ( 
.A(n_6429),
.B(n_6423),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_L g6444 ( 
.A(n_6435),
.B(n_6425),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6442),
.Y(n_6445)
);

OAI21xp5_ASAP7_75t_L g6446 ( 
.A1(n_6438),
.A2(n_6417),
.B(n_6424),
.Y(n_6446)
);

OAI22xp33_ASAP7_75t_SL g6447 ( 
.A1(n_6440),
.A2(n_6436),
.B1(n_6420),
.B2(n_6412),
.Y(n_6447)
);

INVx2_ASAP7_75t_L g6448 ( 
.A(n_6439),
.Y(n_6448)
);

INVxp33_ASAP7_75t_SL g6449 ( 
.A(n_6444),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6445),
.Y(n_6450)
);

AO22x2_ASAP7_75t_L g6451 ( 
.A1(n_6450),
.A2(n_6437),
.B1(n_6441),
.B2(n_6448),
.Y(n_6451)
);

OAI22xp5_ASAP7_75t_SL g6452 ( 
.A1(n_6451),
.A2(n_6449),
.B1(n_6446),
.B2(n_6447),
.Y(n_6452)
);

CKINVDCx20_ASAP7_75t_R g6453 ( 
.A(n_6451),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_6452),
.Y(n_6454)
);

AOI21xp33_ASAP7_75t_SL g6455 ( 
.A1(n_6454),
.A2(n_6453),
.B(n_6443),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6455),
.Y(n_6456)
);

AOI22xp5_ASAP7_75t_L g6457 ( 
.A1(n_6456),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_6457)
);

OR2x2_ASAP7_75t_L g6458 ( 
.A(n_6457),
.B(n_1037),
.Y(n_6458)
);

AOI221xp5_ASAP7_75t_L g6459 ( 
.A1(n_6458),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_6459)
);

AOI211xp5_ASAP7_75t_L g6460 ( 
.A1(n_6459),
.A2(n_231),
.B(n_232),
.C(n_233),
.Y(n_6460)
);


endmodule