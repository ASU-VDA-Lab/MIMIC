module real_aes_15541_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_844, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_844;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g797 ( .A(n_0), .B(n_798), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_1), .A2(n_4), .B1(n_133), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_2), .A2(n_43), .B1(n_140), .B2(n_176), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_3), .A2(n_24), .B1(n_176), .B2(n_218), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_5), .A2(n_15), .B1(n_130), .B2(n_207), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_6), .A2(n_62), .B1(n_190), .B2(n_220), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_7), .A2(n_16), .B1(n_140), .B2(n_161), .Y(n_576) );
INVx1_ASAP7_75t_L g798 ( .A(n_8), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_9), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_10), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_11), .A2(n_17), .B1(n_189), .B2(n_192), .Y(n_188) );
OR2x2_ASAP7_75t_L g790 ( .A(n_12), .B(n_39), .Y(n_790) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_14), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_18), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_19), .A2(n_101), .B1(n_130), .B2(n_133), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_38), .B1(n_165), .B2(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_21), .B(n_131), .Y(n_162) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_22), .A2(n_58), .B(n_149), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_23), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_25), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_26), .B(n_137), .Y(n_496) );
INVx4_ASAP7_75t_R g544 ( .A(n_27), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_28), .A2(n_48), .B1(n_178), .B2(n_179), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_29), .A2(n_55), .B1(n_130), .B2(n_179), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_30), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_31), .B(n_165), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_32), .Y(n_241) );
INVx1_ASAP7_75t_L g475 ( .A(n_33), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_34), .B(n_176), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_SL g487 ( .A1(n_35), .A2(n_136), .B(n_140), .C(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_36), .A2(n_56), .B1(n_140), .B2(n_179), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_37), .A2(n_98), .B1(n_836), .B2(n_840), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_40), .A2(n_89), .B1(n_140), .B2(n_217), .Y(n_216) );
XOR2x2_ASAP7_75t_L g778 ( .A(n_41), .B(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_42), .A2(n_46), .B1(n_140), .B2(n_161), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_44), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_45), .A2(n_60), .B1(n_130), .B2(n_139), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_47), .A2(n_74), .B1(n_780), .B2(n_781), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_47), .Y(n_781) );
INVx1_ASAP7_75t_L g499 ( .A(n_49), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_50), .B(n_140), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_51), .Y(n_516) );
INVx2_ASAP7_75t_L g796 ( .A(n_52), .Y(n_796) );
BUFx3_ASAP7_75t_L g789 ( .A(n_53), .Y(n_789) );
INVx1_ASAP7_75t_L g817 ( .A(n_53), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_54), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_57), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_59), .A2(n_90), .B1(n_140), .B2(n_179), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_61), .A2(n_69), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_61), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_63), .A2(n_78), .B1(n_139), .B2(n_178), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_64), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_65), .A2(n_80), .B1(n_140), .B2(n_161), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_66), .A2(n_100), .B1(n_130), .B2(n_192), .Y(n_238) );
AND2x4_ASAP7_75t_L g126 ( .A(n_67), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g149 ( .A(n_68), .Y(n_149) );
INVx1_ASAP7_75t_L g806 ( .A(n_69), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_70), .A2(n_92), .B1(n_178), .B2(n_179), .Y(n_471) );
AO22x1_ASAP7_75t_L g533 ( .A1(n_71), .A2(n_79), .B1(n_204), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
AND2x2_ASAP7_75t_L g491 ( .A(n_73), .B(n_171), .Y(n_491) );
INVx1_ASAP7_75t_L g780 ( .A(n_74), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_75), .A2(n_778), .B1(n_782), .B2(n_783), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_75), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_76), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_77), .B(n_220), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_81), .B(n_176), .Y(n_517) );
INVx2_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_83), .B(n_171), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_84), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_85), .A2(n_99), .B1(n_179), .B2(n_220), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_86), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_87), .B(n_147), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_88), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_91), .B(n_171), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_93), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_94), .B(n_171), .Y(n_513) );
INVx1_ASAP7_75t_L g112 ( .A(n_95), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_95), .B(n_816), .Y(n_815) );
NAND2xp33_ASAP7_75t_L g167 ( .A(n_96), .B(n_131), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_97), .A2(n_195), .B(n_220), .C(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g546 ( .A(n_98), .B(n_547), .Y(n_546) );
XNOR2xp5_ASAP7_75t_L g819 ( .A(n_98), .B(n_820), .Y(n_819) );
NAND2xp33_ASAP7_75t_L g521 ( .A(n_102), .B(n_166), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_784), .B(n_799), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_777), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_113), .B1(n_453), .B2(n_454), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_110), .Y(n_453) );
BUFx8_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g792 ( .A(n_111), .B(n_788), .Y(n_792) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
XOR2xp5_ASAP7_75t_L g804 ( .A(n_114), .B(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_356), .Y(n_114) );
NAND4xp25_ASAP7_75t_L g115 ( .A(n_116), .B(n_280), .C(n_311), .D(n_340), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_247), .Y(n_116) );
OAI322xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_183), .A3(n_212), .B1(n_225), .B2(n_233), .C1(n_242), .C2(n_244), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_119), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_153), .Y(n_119) );
AND2x2_ASAP7_75t_L g277 ( .A(n_120), .B(n_278), .Y(n_277) );
INVx4_ASAP7_75t_L g313 ( .A(n_120), .Y(n_313) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g288 ( .A(n_121), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g291 ( .A(n_121), .B(n_185), .Y(n_291) );
AND2x2_ASAP7_75t_L g308 ( .A(n_121), .B(n_201), .Y(n_308) );
AND2x2_ASAP7_75t_L g406 ( .A(n_121), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g229 ( .A(n_122), .Y(n_229) );
AND2x4_ASAP7_75t_L g412 ( .A(n_122), .B(n_407), .Y(n_412) );
AO31x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .A3(n_144), .B(n_150), .Y(n_122) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_123), .A2(n_196), .A3(n_237), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_124), .A2(n_539), .B(n_542), .Y(n_538) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_125), .A2(n_174), .A3(n_180), .B(n_181), .Y(n_173) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_125), .A2(n_187), .A3(n_196), .B(n_198), .Y(n_186) );
AO31x2_ASAP7_75t_L g201 ( .A1(n_125), .A2(n_202), .A3(n_209), .B(n_210), .Y(n_201) );
AO31x2_ASAP7_75t_L g574 ( .A1(n_125), .A2(n_152), .A3(n_575), .B(n_578), .Y(n_574) );
BUFx10_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
BUFx10_ASAP7_75t_L g466 ( .A(n_126), .Y(n_466) );
INVx1_ASAP7_75t_L g490 ( .A(n_126), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_135), .B1(n_138), .B2(n_141), .Y(n_128) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_131), .Y(n_534) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g134 ( .A(n_132), .Y(n_134) );
INVx3_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVx1_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
INVx1_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
INVx1_ASAP7_75t_L g208 ( .A(n_132), .Y(n_208) );
INVx2_ASAP7_75t_L g218 ( .A(n_132), .Y(n_218) );
INVx1_ASAP7_75t_L g220 ( .A(n_132), .Y(n_220) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_134), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_135), .A2(n_164), .B(n_167), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_135), .A2(n_141), .B1(n_175), .B2(n_177), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_135), .A2(n_188), .B1(n_193), .B2(n_194), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_135), .A2(n_141), .B1(n_203), .B2(n_206), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_135), .A2(n_216), .B1(n_219), .B2(n_221), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_135), .A2(n_194), .B1(n_238), .B2(n_239), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_135), .A2(n_141), .B1(n_257), .B2(n_258), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_135), .A2(n_463), .B1(n_464), .B2(n_465), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_135), .A2(n_221), .B1(n_471), .B2(n_472), .Y(n_470) );
OAI22x1_ASAP7_75t_L g575 ( .A1(n_135), .A2(n_221), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
O2A1O1Ixp5_ASAP7_75t_L g159 ( .A1(n_136), .A2(n_160), .B(n_161), .C(n_162), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_136), .A2(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_136), .B(n_533), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_136), .A2(n_529), .B(n_533), .C(n_536), .Y(n_590) );
BUFx8_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
INVx1_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
INVx1_ASAP7_75t_L g486 ( .A(n_137), .Y(n_486) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx4_ASAP7_75t_L g161 ( .A(n_140), .Y(n_161) );
INVx1_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g465 ( .A(n_142), .Y(n_465) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g519 ( .A(n_143), .Y(n_519) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_144), .A2(n_222), .A3(n_256), .B(n_259), .Y(n_255) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_144), .A2(n_538), .B(n_546), .Y(n_537) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_146), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_146), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g152 ( .A(n_147), .Y(n_152) );
INVx2_ASAP7_75t_L g197 ( .A(n_147), .Y(n_197) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_147), .A2(n_490), .B(n_531), .Y(n_536) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_152), .B(n_260), .Y(n_259) );
AND2x4_ASAP7_75t_L g417 ( .A(n_153), .B(n_318), .Y(n_417) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g246 ( .A(n_154), .Y(n_246) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_154), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_172), .Y(n_154) );
AND2x2_ASAP7_75t_L g234 ( .A(n_155), .B(n_173), .Y(n_234) );
INVx1_ASAP7_75t_L g275 ( .A(n_155), .Y(n_275) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_170), .Y(n_155) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_156), .A2(n_158), .B(n_170), .Y(n_270) );
INVx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_157), .B(n_182), .Y(n_181) );
BUFx3_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_157), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_157), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g503 ( .A(n_157), .B(n_466), .Y(n_503) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_163), .B(n_168), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_161), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_166), .A2(n_208), .B1(n_544), .B2(n_545), .Y(n_543) );
INVx2_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_SL g222 ( .A(n_169), .Y(n_222) );
INVx2_ASAP7_75t_L g180 ( .A(n_171), .Y(n_180) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_171), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g266 ( .A(n_172), .Y(n_266) );
AND2x2_ASAP7_75t_L g330 ( .A(n_172), .B(n_269), .Y(n_330) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g284 ( .A(n_173), .Y(n_284) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_173), .Y(n_337) );
OR2x2_ASAP7_75t_L g408 ( .A(n_173), .B(n_214), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_176), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g473 ( .A(n_179), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_179), .B(n_498), .Y(n_497) );
AO31x2_ASAP7_75t_L g461 ( .A1(n_180), .A2(n_462), .A3(n_466), .B(n_467), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g286 ( .A(n_183), .B(n_287), .C(n_290), .D(n_292), .Y(n_286) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g424 ( .A(n_184), .B(n_412), .Y(n_424) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_185), .B(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g278 ( .A(n_185), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g298 ( .A(n_185), .Y(n_298) );
INVx1_ASAP7_75t_L g315 ( .A(n_185), .Y(n_315) );
INVx1_ASAP7_75t_L g323 ( .A(n_185), .Y(n_323) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_185), .Y(n_437) );
INVx4_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_186), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g355 ( .A(n_186), .B(n_255), .Y(n_355) );
AND2x2_ASAP7_75t_L g363 ( .A(n_186), .B(n_201), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_186), .B(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g428 ( .A(n_186), .Y(n_428) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_191), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g221 ( .A(n_195), .Y(n_221) );
AO31x2_ASAP7_75t_L g469 ( .A1(n_196), .A2(n_222), .A3(n_470), .B(n_474), .Y(n_469) );
AOI21x1_ASAP7_75t_L g478 ( .A1(n_196), .A2(n_479), .B(n_491), .Y(n_478) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_197), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_197), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g547 ( .A(n_197), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_197), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g232 ( .A(n_201), .Y(n_232) );
OR2x2_ASAP7_75t_L g293 ( .A(n_201), .B(n_255), .Y(n_293) );
INVx2_ASAP7_75t_L g300 ( .A(n_201), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_201), .B(n_253), .Y(n_324) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_201), .Y(n_411) );
OAI21xp33_ASAP7_75t_SL g495 ( .A1(n_204), .A2(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_209), .A2(n_215), .A3(n_222), .B(n_223), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_212), .B(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g235 ( .A(n_214), .B(n_236), .Y(n_235) );
BUFx2_ASAP7_75t_L g245 ( .A(n_214), .Y(n_245) );
INVx2_ASAP7_75t_L g263 ( .A(n_214), .Y(n_263) );
AND2x4_ASAP7_75t_L g295 ( .A(n_214), .B(n_267), .Y(n_295) );
OR2x2_ASAP7_75t_L g375 ( .A(n_214), .B(n_275), .Y(n_375) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_218), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_221), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_230), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_227), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g292 ( .A(n_227), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_227), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_228), .B(n_298), .Y(n_306) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g251 ( .A(n_229), .Y(n_251) );
OR2x2_ASAP7_75t_L g344 ( .A(n_229), .B(n_254), .Y(n_344) );
INVx1_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g243 ( .A(n_231), .Y(n_243) );
INVx1_ASAP7_75t_L g279 ( .A(n_232), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
OAI322xp33_ASAP7_75t_L g247 ( .A1(n_234), .A2(n_248), .A3(n_261), .B1(n_264), .B2(n_271), .C1(n_272), .C2(n_276), .Y(n_247) );
AND2x4_ASAP7_75t_L g294 ( .A(n_234), .B(n_295), .Y(n_294) );
AOI211xp5_ASAP7_75t_SL g325 ( .A1(n_234), .A2(n_326), .B(n_327), .C(n_331), .Y(n_325) );
AND2x2_ASAP7_75t_L g345 ( .A(n_234), .B(n_235), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_234), .B(n_262), .Y(n_351) );
AND2x4_ASAP7_75t_SL g273 ( .A(n_235), .B(n_274), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g364 ( .A(n_235), .B(n_291), .C(n_319), .Y(n_364) );
AND2x2_ASAP7_75t_L g395 ( .A(n_235), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g262 ( .A(n_236), .B(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g267 ( .A(n_236), .Y(n_267) );
BUFx2_ASAP7_75t_L g335 ( .A(n_236), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_245), .B(n_269), .Y(n_268) );
NAND2x1_ASAP7_75t_L g309 ( .A(n_245), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_246), .B(n_262), .Y(n_393) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g336 ( .A(n_251), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
AND2x4_ASAP7_75t_L g299 ( .A(n_255), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g386 ( .A(n_255), .Y(n_386) );
INVx2_ASAP7_75t_L g407 ( .A(n_255), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_261), .A2(n_420), .B1(n_422), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g331 ( .A(n_262), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g285 ( .A(n_263), .B(n_269), .Y(n_285) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g304 ( .A(n_265), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x4_ASAP7_75t_L g274 ( .A(n_266), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g396 ( .A(n_266), .Y(n_396) );
INVx2_ASAP7_75t_L g282 ( .A(n_267), .Y(n_282) );
AND2x2_ASAP7_75t_L g310 ( .A(n_267), .B(n_269), .Y(n_310) );
INVx3_ASAP7_75t_L g318 ( .A(n_267), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_267), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g303 ( .A(n_268), .Y(n_303) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
OAI222xp33_ASAP7_75t_L g442 ( .A1(n_272), .A2(n_432), .B1(n_443), .B2(n_446), .C1(n_448), .C2(n_450), .Y(n_442) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g383 ( .A(n_274), .Y(n_383) );
AND2x2_ASAP7_75t_L g447 ( .A(n_274), .B(n_317), .Y(n_447) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_277), .B(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_286), .B1(n_294), .B2(n_296), .C(n_301), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g369 ( .A(n_282), .Y(n_369) );
INVx2_ASAP7_75t_L g431 ( .A(n_283), .Y(n_431) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g332 ( .A(n_284), .Y(n_332) );
AND2x2_ASAP7_75t_L g368 ( .A(n_284), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g334 ( .A(n_285), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g360 ( .A(n_285), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g449 ( .A(n_285), .Y(n_449) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g398 ( .A(n_289), .Y(n_398) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g421 ( .A(n_291), .B(n_299), .Y(n_421) );
AND2x2_ASAP7_75t_L g444 ( .A(n_291), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g305 ( .A(n_293), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g440 ( .A(n_293), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_294), .A2(n_348), .B1(n_382), .B2(n_384), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g409 ( .A1(n_294), .A2(n_410), .B(n_413), .Y(n_409) );
INVxp67_ASAP7_75t_L g326 ( .A(n_295), .Y(n_326) );
INVx2_ASAP7_75t_SL g430 ( .A(n_295), .Y(n_430) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OR2x2_ASAP7_75t_L g343 ( .A(n_297), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g441 ( .A(n_297), .B(n_440), .Y(n_441) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g314 ( .A(n_299), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_299), .B(n_323), .Y(n_339) );
INVx2_ASAP7_75t_L g366 ( .A(n_299), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B1(n_307), .B2(n_309), .Y(n_301) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_303), .A2(n_377), .B1(n_390), .B2(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g399 ( .A(n_308), .B(n_400), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B(n_320), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g380 ( .A(n_313), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_313), .B(n_363), .Y(n_391) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_317), .B(n_330), .Y(n_422) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_318), .A2(n_436), .B(n_438), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_325), .B(n_333), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g379 ( .A(n_324), .Y(n_379) );
INVx1_ASAP7_75t_L g445 ( .A(n_324), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g418 ( .A(n_328), .Y(n_418) );
OR2x2_ASAP7_75t_L g429 ( .A(n_329), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .C(n_338), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_334), .A2(n_395), .B1(n_397), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_336), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g374 ( .A(n_337), .Y(n_374) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_339), .B(n_343), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_339), .A2(n_402), .B1(n_405), .B2(n_408), .C(n_409), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B(n_346), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g350 ( .A(n_344), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_351), .B1(n_352), .B2(n_844), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g433 ( .A(n_355), .B(n_411), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_387), .C(n_414), .D(n_434), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_370), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_364), .B2(n_365), .C(n_367), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_360), .A2(n_417), .B1(n_439), .B2(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g413 ( .A(n_362), .Y(n_413) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g397 ( .A(n_363), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_363), .B(n_406), .Y(n_405) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_363), .B(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_365), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g372 ( .A(n_369), .B(n_373), .Y(n_372) );
OAI21xp33_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_376), .B(n_381), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2x1_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g400 ( .A(n_386), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_415), .B(n_419), .C(n_425), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_401), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_389), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g448 ( .A(n_396), .B(n_449), .Y(n_448) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx3_ASAP7_75t_L g452 ( .A(n_412), .Y(n_452) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp33_ASAP7_75t_R g425 ( .A1(n_426), .A2(n_429), .B1(n_431), .B2(n_432), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g439 ( .A(n_428), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_442), .Y(n_434) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_669), .Y(n_454) );
NOR2xp67_ASAP7_75t_L g455 ( .A(n_456), .B(n_611), .Y(n_455) );
NAND3xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_548), .C(n_593), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_504), .B(n_525), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_458), .A2(n_549), .B1(n_568), .B2(n_580), .Y(n_548) );
AOI22x1_ASAP7_75t_L g673 ( .A1(n_458), .A2(n_674), .B1(n_678), .B2(n_679), .Y(n_673) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_476), .Y(n_459) );
OR2x2_ASAP7_75t_L g634 ( .A(n_460), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_469), .Y(n_460) );
OR2x2_ASAP7_75t_L g509 ( .A(n_461), .B(n_469), .Y(n_509) );
AND2x2_ASAP7_75t_L g552 ( .A(n_461), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g560 ( .A(n_461), .Y(n_560) );
BUFx2_ASAP7_75t_L g610 ( .A(n_461), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_465), .A2(n_501), .B(n_502), .Y(n_500) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_465), .A2(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
AND2x2_ASAP7_75t_L g555 ( .A(n_469), .B(n_492), .Y(n_555) );
INVx1_ASAP7_75t_L g562 ( .A(n_469), .Y(n_562) );
INVx1_ASAP7_75t_L g567 ( .A(n_469), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_469), .B(n_560), .Y(n_629) );
INVx1_ASAP7_75t_L g650 ( .A(n_469), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_469), .B(n_553), .Y(n_720) );
INVx1_ASAP7_75t_L g613 ( .A(n_476), .Y(n_613) );
OR2x2_ASAP7_75t_L g665 ( .A(n_476), .B(n_629), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_492), .Y(n_476) );
AND2x2_ASAP7_75t_L g510 ( .A(n_477), .B(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g558 ( .A(n_477), .B(n_559), .Y(n_558) );
INVxp67_ASAP7_75t_L g564 ( .A(n_477), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_477), .B(n_507), .Y(n_641) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g553 ( .A(n_478), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_487), .B(n_490), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B(n_485), .Y(n_480) );
BUFx4f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_486), .B(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g507 ( .A(n_492), .Y(n_507) );
INVx1_ASAP7_75t_L g607 ( .A(n_492), .Y(n_607) );
AND2x2_ASAP7_75t_L g609 ( .A(n_492), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g627 ( .A(n_492), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g649 ( .A(n_492), .B(n_650), .Y(n_649) );
NAND2x1p5_ASAP7_75t_SL g660 ( .A(n_492), .B(n_636), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_492), .B(n_567), .Y(n_750) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_500), .B(n_503), .Y(n_494) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_505), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_688) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_506), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_506), .B(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g767 ( .A(n_506), .B(n_625), .Y(n_767) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g566 ( .A(n_507), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_507), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g655 ( .A(n_507), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g606 ( .A(n_508), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g696 ( .A(n_509), .Y(n_696) );
OR2x2_ASAP7_75t_L g770 ( .A(n_509), .B(n_697), .Y(n_770) );
INVx1_ASAP7_75t_L g601 ( .A(n_510), .Y(n_601) );
INVx3_ASAP7_75t_L g605 ( .A(n_511), .Y(n_605) );
BUFx2_ASAP7_75t_L g616 ( .A(n_511), .Y(n_616) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g586 ( .A(n_512), .B(n_537), .Y(n_586) );
INVx2_ASAP7_75t_L g632 ( .A(n_512), .Y(n_632) );
INVx1_ASAP7_75t_L g664 ( .A(n_512), .Y(n_664) );
AND2x2_ASAP7_75t_L g677 ( .A(n_512), .B(n_574), .Y(n_677) );
AND2x2_ASAP7_75t_L g699 ( .A(n_512), .B(n_598), .Y(n_699) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_520), .B(n_523), .Y(n_514) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g690 ( .A(n_526), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_526), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g715 ( .A(n_526), .B(n_583), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_526), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
INVx2_ASAP7_75t_L g572 ( .A(n_527), .Y(n_572) );
AND2x2_ASAP7_75t_L g599 ( .A(n_527), .B(n_600), .Y(n_599) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_532), .B(n_535), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g573 ( .A(n_537), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g592 ( .A(n_537), .Y(n_592) );
INVx2_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
OR2x2_ASAP7_75t_L g620 ( .A(n_537), .B(n_574), .Y(n_620) );
AND2x2_ASAP7_75t_L g631 ( .A(n_537), .B(n_632), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B1(n_556), .B2(n_561), .C(n_563), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI32xp33_ASAP7_75t_L g661 ( .A1(n_551), .A2(n_565), .A3(n_662), .B1(n_665), .B2(n_666), .Y(n_661) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g651 ( .A(n_552), .Y(n_651) );
AND2x2_ASAP7_75t_L g687 ( .A(n_552), .B(n_566), .Y(n_687) );
INVx1_ASAP7_75t_L g751 ( .A(n_552), .Y(n_751) );
OR2x2_ASAP7_75t_L g625 ( .A(n_553), .B(n_560), .Y(n_625) );
INVx2_ASAP7_75t_L g636 ( .A(n_553), .Y(n_636) );
BUFx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g775 ( .A(n_555), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVxp67_ASAP7_75t_L g762 ( .A(n_558), .Y(n_762) );
INVx1_ASAP7_75t_L g776 ( .A(n_558), .Y(n_776) );
OR2x2_ASAP7_75t_L g656 ( .A(n_559), .B(n_636), .Y(n_656) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_561), .B(n_656), .Y(n_678) );
INVx1_ASAP7_75t_L g709 ( .A(n_561), .Y(n_709) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g743 ( .A(n_562), .Y(n_743) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2x1_ASAP7_75t_L g712 ( .A(n_564), .B(n_713), .Y(n_712) );
OAI21xp5_ASAP7_75t_SL g734 ( .A1(n_565), .A2(n_735), .B(n_740), .Y(n_734) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
AND2x2_ASAP7_75t_L g644 ( .A(n_570), .B(n_586), .Y(n_644) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_570), .Y(n_774) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g676 ( .A(n_571), .Y(n_676) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g658 ( .A(n_572), .B(n_632), .Y(n_658) );
AND2x2_ASAP7_75t_L g729 ( .A(n_572), .B(n_600), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_573), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g657 ( .A(n_573), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g736 ( .A(n_573), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g585 ( .A(n_574), .Y(n_585) );
INVx2_ASAP7_75t_L g598 ( .A(n_574), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_574), .B(n_589), .Y(n_646) );
AND2x2_ASAP7_75t_L g706 ( .A(n_574), .B(n_600), .Y(n_706) );
NAND2xp33_ASAP7_75t_SL g580 ( .A(n_581), .B(n_587), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g681 ( .A(n_584), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_584), .B(n_664), .Y(n_756) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g588 ( .A(n_585), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g717 ( .A(n_585), .B(n_632), .Y(n_717) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
OR2x2_ASAP7_75t_L g662 ( .A(n_588), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g619 ( .A(n_589), .Y(n_619) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g645 ( .A(n_592), .B(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_606), .B1(n_608), .B2(n_609), .Y(n_593) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_601), .B(n_602), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g608 ( .A(n_596), .B(n_605), .Y(n_608) );
BUFx2_ASAP7_75t_L g626 ( .A(n_596), .Y(n_626) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g637 ( .A(n_597), .Y(n_637) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g652 ( .A(n_599), .B(n_616), .Y(n_652) );
INVx2_ASAP7_75t_L g668 ( .A(n_599), .Y(n_668) );
AND2x2_ASAP7_75t_L g710 ( .A(n_599), .B(n_632), .Y(n_710) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g685 ( .A(n_605), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g732 ( .A(n_606), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g763 ( .A(n_607), .Y(n_763) );
INVx2_ASAP7_75t_L g702 ( .A(n_610), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_621), .C(n_638), .D(n_653), .Y(n_611) );
NAND2xp33_ASAP7_75t_SL g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_614), .A2(n_692), .B1(n_708), .B2(n_710), .C(n_711), .Y(n_707) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g689 ( .A(n_618), .Y(n_689) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g682 ( .A(n_619), .Y(n_682) );
INVx2_ASAP7_75t_L g754 ( .A(n_620), .Y(n_754) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_626), .B1(n_627), .B2(n_630), .C1(n_633), .C2(n_637), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g708 ( .A(n_624), .B(n_709), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_624), .A2(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g747 ( .A(n_625), .B(n_691), .Y(n_747) );
OAI21xp33_ASAP7_75t_SL g721 ( .A1(n_626), .A2(n_647), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g640 ( .A(n_629), .B(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_629), .Y(n_692) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g691 ( .A(n_632), .Y(n_691) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g697 ( .A(n_636), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_642), .B1(n_647), .B2(n_652), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_644), .A2(n_654), .B1(n_657), .B2(n_659), .C(n_661), .Y(n_653) );
INVx3_ASAP7_75t_R g768 ( .A(n_645), .Y(n_768) );
INVx1_ASAP7_75t_L g686 ( .A(n_646), .Y(n_686) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_649), .Y(n_703) );
INVx1_ASAP7_75t_L g713 ( .A(n_649), .Y(n_713) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_658), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g731 ( .A(n_658), .Y(n_731) );
AND2x2_ASAP7_75t_L g759 ( .A(n_658), .B(n_706), .Y(n_759) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g753 ( .A(n_663), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_725), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_707), .C(n_721), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_683), .C(n_693), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_674), .A2(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g724 ( .A(n_676), .Y(n_724) );
AND2x2_ASAP7_75t_L g765 ( .A(n_676), .B(n_754), .Y(n_765) );
NAND2x1_ASAP7_75t_L g723 ( .A(n_677), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g745 ( .A(n_682), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g737 ( .A(n_691), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_698), .B1(n_700), .B2(n_704), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g733 ( .A(n_697), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_699), .B(n_729), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g772 ( .A(n_705), .Y(n_772) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI22xp33_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_714), .B1(n_716), .B2(n_718), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_752), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B(n_732), .C(n_734), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g741 ( .A1(n_728), .A2(n_742), .B(n_744), .Y(n_741) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
O2A1O1Ixp5_ASAP7_75t_SL g752 ( .A1(n_732), .A2(n_753), .B(n_755), .C(n_757), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_736), .A2(n_741), .B1(n_746), .B2(n_748), .Y(n_740) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_764), .C(n_771), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_768), .B2(n_769), .Y(n_764) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI21xp5_ASAP7_75t_SL g771 ( .A1(n_772), .A2(n_773), .B(n_775), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g783 ( .A(n_778), .Y(n_783) );
BUFx4f_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx3_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_791), .Y(n_786) );
BUFx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g818 ( .A(n_790), .Y(n_818) );
OR2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
AND2x2_ASAP7_75t_L g836 ( .A(n_792), .B(n_837), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_793), .B(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_794), .B(n_797), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_795), .B(n_833), .Y(n_832) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_796), .B(n_826), .Y(n_842) );
INVx2_ASAP7_75t_SL g834 ( .A(n_797), .Y(n_834) );
OAI21xp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_828), .B(n_835), .Y(n_799) );
OAI22xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B1(n_808), .B2(n_823), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_819), .B(n_821), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx4_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_812), .B(n_822), .Y(n_821) );
BUFx12f_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx4_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx3_ASAP7_75t_L g826 ( .A(n_814), .Y(n_826) );
CKINVDCx8_ASAP7_75t_R g839 ( .A(n_814), .Y(n_839) );
AND2x6_ASAP7_75t_SL g814 ( .A(n_815), .B(n_818), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_819), .A2(n_824), .B(n_827), .Y(n_823) );
INVxp67_ASAP7_75t_L g827 ( .A(n_821), .Y(n_827) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
BUFx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
INVx4_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
BUFx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OR2x4_ASAP7_75t_L g841 ( .A(n_833), .B(n_842), .Y(n_841) );
BUFx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx3_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
endmodule