module fake_jpeg_10102_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_47),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_23),
.B(n_22),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_23),
.A3(n_32),
.B1(n_19),
.B2(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_22),
.B(n_34),
.C(n_17),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_16),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_63),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_34),
.B1(n_19),
.B2(n_21),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_57),
.B1(n_39),
.B2(n_23),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_62),
.Y(n_70)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_34),
.B1(n_19),
.B2(n_17),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_56),
.B1(n_52),
.B2(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_16),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_65),
.B(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_68),
.B(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_75),
.Y(n_117)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_21),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_86),
.B(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_51),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_42),
.B(n_14),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_60),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_37),
.B1(n_18),
.B2(n_33),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_90),
.B1(n_96),
.B2(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_16),
.B1(n_18),
.B2(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_58),
.B1(n_54),
.B2(n_60),
.Y(n_111)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_29),
.B(n_39),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_111),
.B1(n_113),
.B2(n_123),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_104),
.B(n_110),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_14),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_67),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_65),
.B(n_92),
.C(n_85),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_42),
.B1(n_60),
.B2(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_67),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_20),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_84),
.B(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_135),
.Y(n_173)
);

CKINVDCx6p67_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_79),
.B(n_93),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_132),
.B(n_105),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_78),
.B(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_83),
.B1(n_77),
.B2(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_137),
.B1(n_139),
.B2(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_98),
.B1(n_66),
.B2(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_140),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_96),
.B1(n_86),
.B2(n_87),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_65),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_107),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_146),
.C(n_20),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_72),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_73),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_149),
.B(n_115),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_92),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_75),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_104),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_15),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_156),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_75),
.B1(n_89),
.B2(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_94),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_29),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_28),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_158),
.A2(n_160),
.B(n_167),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_137),
.B1(n_139),
.B2(n_136),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_163),
.B1(n_166),
.B2(n_175),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_122),
.B1(n_106),
.B2(n_125),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_123),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_184),
.C(n_138),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_106),
.B1(n_120),
.B2(n_99),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_101),
.B(n_99),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_127),
.A2(n_135),
.B1(n_134),
.B2(n_147),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_181),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_102),
.A3(n_24),
.B1(n_27),
.B2(n_28),
.C1(n_26),
.C2(n_25),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_128),
.C(n_145),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_24),
.B(n_20),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_180),
.A2(n_186),
.B(n_189),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_0),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_190),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_82),
.B(n_102),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_199),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_204),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_142),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_200),
.C(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_157),
.B1(n_152),
.B2(n_149),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_206),
.B1(n_162),
.B2(n_167),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_128),
.B1(n_157),
.B2(n_141),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_208),
.B(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_160),
.C(n_171),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_12),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_12),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_214),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_12),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_11),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_185),
.B1(n_161),
.B2(n_159),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_235),
.B1(n_237),
.B2(n_199),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_26),
.Y(n_256)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_158),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_231),
.C(n_238),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_170),
.B1(n_188),
.B2(n_164),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_162),
.B(n_187),
.C(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_213),
.B1(n_216),
.B2(n_205),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_201),
.A2(n_170),
.B1(n_188),
.B2(n_168),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_233),
.B1(n_220),
.B2(n_224),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_186),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_201),
.A2(n_168),
.B1(n_172),
.B2(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_186),
.B1(n_178),
.B2(n_180),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_114),
.B1(n_82),
.B2(n_28),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_216),
.C(n_196),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_1),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_241),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_256),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_203),
.B(n_194),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_218),
.B(n_230),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_203),
.B1(n_197),
.B2(n_195),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_206),
.C(n_192),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_251),
.C(n_253),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_114),
.C(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_114),
.B1(n_26),
.B2(n_25),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_229),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_25),
.C(n_2),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_256),
.C(n_247),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_6),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_267),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_263),
.B(n_235),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_228),
.B(n_240),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_236),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_237),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_233),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_282),
.B(n_10),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_221),
.C(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_249),
.B1(n_251),
.B2(n_238),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_280),
.B1(n_10),
.B2(n_2),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_253),
.B1(n_242),
.B2(n_9),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_285),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_242),
.B1(n_6),
.B2(n_9),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_14),
.B(n_13),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_10),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_286),
.C(n_265),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_265),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_6),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_261),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_293),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_268),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_290),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_295),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_296),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_1),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_1),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_2),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_284),
.C(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_282),
.C(n_3),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_296),
.C(n_293),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_4),
.B(n_5),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_306),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_3),
.B(n_4),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_299),
.C(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_305),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_309),
.B(n_300),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_311),
.B(n_4),
.CI(n_274),
.CON(n_312),
.SN(n_312)
);


endmodule