module real_aes_8551_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_852;
wire n_766;
wire n_974;
wire n_919;
wire n_1089;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_666;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_816;
wire n_400;
wire n_539;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_994;
wire n_495;
wire n_1078;
wire n_892;
wire n_370;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_1053;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_1025;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_973;
wire n_504;
wire n_671;
wire n_960;
wire n_1084;
wire n_1081;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_913;
wire n_490;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_598;
wire n_404;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_1056;
wire n_749;
wire n_385;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_507;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1102;
wire n_1076;
wire n_463;
wire n_661;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_0), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_1), .A2(n_281), .B1(n_621), .B2(n_769), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_2), .A2(n_157), .B1(n_529), .B2(n_537), .Y(n_1042) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_3), .Y(n_618) );
INVx1_ASAP7_75t_L g1037 ( .A(n_4), .Y(n_1037) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_5), .A2(n_337), .B1(n_480), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_6), .A2(n_130), .B1(n_529), .B2(n_793), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_7), .Y(n_435) );
AOI222xp33_ASAP7_75t_L g513 ( .A1(n_8), .A2(n_183), .B1(n_285), .B2(n_419), .C1(n_514), .C2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_9), .A2(n_100), .B1(n_528), .B2(n_709), .Y(n_1022) );
AO22x2_ASAP7_75t_L g393 ( .A1(n_10), .A2(n_215), .B1(n_394), .B2(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g1067 ( .A(n_10), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_11), .A2(n_147), .B1(n_451), .B2(n_493), .Y(n_788) );
AOI222xp33_ASAP7_75t_L g889 ( .A1(n_12), .A2(n_313), .B1(n_324), .B2(n_418), .C1(n_425), .C2(n_758), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_13), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_14), .A2(n_208), .B1(n_528), .B2(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g746 ( .A(n_15), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_16), .A2(n_51), .B1(n_780), .B2(n_1050), .Y(n_1049) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_17), .A2(n_190), .B1(n_644), .B2(n_863), .C(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g728 ( .A(n_18), .Y(n_728) );
INVx1_ASAP7_75t_L g734 ( .A(n_19), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_20), .A2(n_235), .B1(n_591), .B2(n_592), .Y(n_1007) );
XOR2xp5_ASAP7_75t_L g1070 ( .A(n_21), .B(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g950 ( .A(n_22), .Y(n_950) );
AOI22xp5_ASAP7_75t_SL g699 ( .A1(n_23), .A2(n_186), .B1(n_610), .B2(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_24), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_25), .A2(n_349), .B1(n_821), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_26), .A2(n_91), .B1(n_418), .B2(n_425), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_27), .A2(n_200), .B1(n_591), .B2(n_592), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_28), .A2(n_304), .B1(n_489), .B2(n_660), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1038 ( .A1(n_29), .A2(n_187), .B1(n_427), .B2(n_536), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_30), .A2(n_111), .B1(n_479), .B2(n_481), .C(n_483), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_31), .A2(n_151), .B1(n_616), .B2(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_32), .A2(n_309), .B1(n_780), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_33), .A2(n_113), .B1(n_643), .B2(n_770), .Y(n_944) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_34), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_35), .A2(n_134), .B1(n_646), .B2(n_1025), .Y(n_1024) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_36), .A2(n_119), .B1(n_394), .B2(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_37), .A2(n_256), .B1(n_451), .B2(n_542), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g797 ( .A1(n_38), .A2(n_184), .B1(n_284), .B2(n_427), .C1(n_675), .C2(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_39), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_40), .B(n_1021), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_41), .A2(n_75), .B1(n_491), .B2(n_542), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_42), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_43), .A2(n_194), .B1(n_503), .B2(n_506), .C(n_509), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_44), .B(n_574), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_45), .Y(n_973) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_46), .A2(n_126), .B1(n_675), .B2(n_765), .Y(n_1082) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_47), .A2(n_307), .B1(n_444), .B2(n_685), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_48), .A2(n_97), .B1(n_542), .B2(n_550), .Y(n_819) );
AOI222xp33_ASAP7_75t_L g631 ( .A1(n_49), .A2(n_78), .B1(n_133), .B2(n_632), .C1(n_633), .C2(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g722 ( .A(n_50), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_52), .A2(n_142), .B1(n_643), .B2(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g681 ( .A(n_53), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_54), .B(n_633), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_55), .A2(n_268), .B1(n_666), .B2(n_863), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_56), .A2(n_221), .B1(n_471), .B2(n_542), .Y(n_1048) );
AO22x1_ASAP7_75t_L g952 ( .A1(n_57), .A2(n_953), .B1(n_982), .B2(n_983), .Y(n_952) );
INVx1_ASAP7_75t_L g982 ( .A(n_57), .Y(n_982) );
AOI222xp33_ASAP7_75t_L g871 ( .A1(n_58), .A2(n_173), .B1(n_334), .B2(n_412), .C1(n_714), .C2(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_59), .A2(n_93), .B1(n_455), .B2(n_835), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_60), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_61), .A2(n_301), .B1(n_471), .B2(n_489), .Y(n_947) );
INVx1_ASAP7_75t_L g499 ( .A(n_62), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_63), .A2(n_179), .B1(n_528), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_64), .A2(n_84), .B1(n_625), .B2(n_626), .Y(n_837) );
INVx1_ASAP7_75t_L g552 ( .A(n_65), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_66), .B(n_625), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_67), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_68), .A2(n_364), .B1(n_479), .B2(n_1030), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_69), .A2(n_158), .B1(n_1025), .B2(n_1087), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_70), .A2(n_218), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_71), .A2(n_283), .B1(n_550), .B2(n_1092), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_72), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_73), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_74), .A2(n_327), .B1(n_860), .B2(n_863), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_76), .A2(n_360), .B1(n_653), .B2(n_675), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_77), .Y(n_940) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_79), .A2(n_245), .B1(n_481), .B2(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_80), .Y(n_903) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_81), .A2(n_368), .B(n_376), .C(n_1069), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_82), .A2(n_201), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_83), .A2(n_265), .B1(n_529), .B2(n_765), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_85), .A2(n_191), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_86), .A2(n_109), .B1(n_489), .B2(n_491), .C(n_494), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_87), .Y(n_852) );
AO22x2_ASAP7_75t_L g401 ( .A1(n_88), .A2(n_248), .B1(n_394), .B2(n_395), .Y(n_401) );
INVx1_ASAP7_75t_L g1064 ( .A(n_88), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_89), .A2(n_105), .B1(n_491), .B2(n_657), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_90), .A2(n_226), .B1(n_481), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_92), .A2(n_209), .B1(n_709), .B2(n_710), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_94), .A2(n_269), .B1(n_469), .B2(n_471), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_95), .A2(n_127), .B1(n_503), .B2(n_626), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_96), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_98), .A2(n_259), .B1(n_536), .B2(n_537), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_99), .A2(n_180), .B1(n_624), .B2(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_101), .A2(n_848), .B1(n_873), .B2(n_874), .Y(n_847) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_101), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_102), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_103), .A2(n_357), .B1(n_419), .B2(n_793), .Y(n_792) );
AOI222xp33_ASAP7_75t_L g822 ( .A1(n_104), .A2(n_115), .B1(n_174), .B2(n_425), .C1(n_514), .C2(n_823), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_106), .A2(n_988), .B1(n_1008), .B2(n_1009), .Y(n_987) );
INVx1_ASAP7_75t_L g1008 ( .A(n_106), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_107), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_108), .A2(n_250), .B1(n_551), .B2(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g510 ( .A(n_110), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_112), .Y(n_900) );
INVx1_ASAP7_75t_L g712 ( .A(n_114), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_116), .A2(n_263), .B1(n_444), .B2(n_447), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_117), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_118), .A2(n_254), .B1(n_473), .B2(n_548), .Y(n_698) );
INVx1_ASAP7_75t_L g1068 ( .A(n_119), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_120), .A2(n_288), .B1(n_479), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_121), .A2(n_262), .B1(n_462), .B2(n_465), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_122), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_123), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_124), .Y(n_914) );
AO22x1_ASAP7_75t_L g824 ( .A1(n_125), .A2(n_825), .B1(n_826), .B2(n_840), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_125), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_128), .A2(n_145), .B1(n_456), .B2(n_821), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_129), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_131), .A2(n_338), .B1(n_469), .B2(n_480), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_132), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_135), .A2(n_139), .B1(n_444), .B2(n_447), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g907 ( .A(n_136), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_137), .A2(n_477), .B1(n_516), .B2(n_517), .Y(n_476) );
INVx1_ASAP7_75t_L g516 ( .A(n_137), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_138), .Y(n_968) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_140), .A2(n_267), .B1(n_610), .B2(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g495 ( .A(n_141), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_143), .A2(n_335), .B1(n_450), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_144), .A2(n_155), .B1(n_610), .B2(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_146), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_148), .A2(n_198), .B1(n_675), .B2(n_793), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_149), .A2(n_291), .B1(n_657), .B2(n_770), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_150), .A2(n_239), .B1(n_450), .B2(n_455), .Y(n_449) );
AND2x6_ASAP7_75t_L g370 ( .A(n_152), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g1061 ( .A(n_152), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_153), .A2(n_272), .B1(n_648), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_154), .A2(n_318), .B1(n_419), .B2(n_427), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_156), .A2(n_251), .B1(n_574), .B2(n_742), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_159), .A2(n_323), .B1(n_610), .B2(n_725), .Y(n_724) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_160), .A2(n_231), .B1(n_247), .B2(n_412), .C1(n_419), .C2(n_574), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_161), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_162), .A2(n_300), .B1(n_643), .B2(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g689 ( .A(n_163), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_164), .A2(n_330), .B1(n_465), .B2(n_730), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_165), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_166), .A2(n_347), .B1(n_545), .B2(n_821), .Y(n_1046) );
INVx1_ASAP7_75t_L g981 ( .A(n_167), .Y(n_981) );
INVx1_ASAP7_75t_L g745 ( .A(n_168), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_169), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_170), .A2(n_305), .B1(n_465), .B2(n_644), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_171), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_172), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_175), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_176), .A2(n_340), .B1(n_447), .B2(n_949), .Y(n_948) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_177), .A2(n_238), .B1(n_394), .B2(n_398), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_177), .B(n_1066), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_178), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_181), .A2(n_356), .B1(n_659), .B2(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g1016 ( .A(n_182), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_185), .Y(n_760) );
AOI222xp33_ASAP7_75t_L g839 ( .A1(n_188), .A2(n_317), .B1(n_329), .B2(n_514), .C1(n_515), .C2(n_536), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_189), .A2(n_241), .B1(n_585), .B2(n_657), .Y(n_656) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_192), .B(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_193), .A2(n_294), .B1(n_532), .B2(n_651), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_195), .Y(n_799) );
OA22x2_ASAP7_75t_L g717 ( .A1(n_196), .A2(n_718), .B1(n_719), .B2(n_749), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_196), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_197), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_199), .A2(n_282), .B1(n_583), .B2(n_643), .C(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_202), .A2(n_203), .B1(n_550), .B2(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g683 ( .A(n_204), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_205), .A2(n_289), .B1(n_532), .B2(n_534), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_206), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_207), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_210), .A2(n_253), .B1(n_480), .B2(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_211), .B(n_651), .Y(n_1019) );
INVx1_ASAP7_75t_L g920 ( .A(n_212), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_213), .A2(n_280), .B1(n_481), .B2(n_816), .Y(n_815) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_214), .A2(n_237), .B1(n_527), .B2(n_528), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_216), .A2(n_303), .B1(n_529), .B2(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_217), .A2(n_271), .B1(n_545), .B2(n_646), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_219), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_220), .A2(n_273), .B1(n_551), .B2(n_685), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_222), .A2(n_355), .B1(n_456), .B2(n_548), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_223), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g1078 ( .A(n_224), .Y(n_1078) );
INVx1_ASAP7_75t_L g678 ( .A(n_225), .Y(n_678) );
INVx1_ASAP7_75t_L g512 ( .A(n_227), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_228), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_229), .A2(n_322), .B1(n_419), .B2(n_793), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_230), .A2(n_249), .B1(n_456), .B2(n_821), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_232), .A2(n_366), .B1(n_624), .B2(n_626), .C(n_627), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_233), .A2(n_339), .B1(n_350), .B2(n_412), .C1(n_515), .C2(n_536), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_234), .A2(n_363), .B1(n_506), .B2(n_624), .Y(n_1083) );
INVx2_ASAP7_75t_L g375 ( .A(n_236), .Y(n_375) );
INVx1_ASAP7_75t_L g1103 ( .A(n_240), .Y(n_1103) );
XNOR2xp5_ASAP7_75t_L g1104 ( .A(n_240), .B(n_1073), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_242), .A2(n_383), .B1(n_384), .B2(n_474), .Y(n_382) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_242), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_243), .A2(n_286), .B1(n_427), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_244), .A2(n_352), .B1(n_583), .B2(n_589), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_246), .Y(n_569) );
INVx1_ASAP7_75t_L g941 ( .A(n_252), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_255), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_257), .A2(n_559), .B1(n_593), .B2(n_594), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_257), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_258), .Y(n_404) );
INVx1_ASAP7_75t_L g723 ( .A(n_260), .Y(n_723) );
XOR2x2_ASAP7_75t_L g1012 ( .A(n_261), .B(n_1013), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_264), .Y(n_628) );
OA22x2_ASAP7_75t_L g752 ( .A1(n_266), .A2(n_753), .B1(n_754), .B2(n_781), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_266), .Y(n_753) );
INVx1_ASAP7_75t_L g394 ( .A(n_270), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_270), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_274), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_275), .A2(n_331), .B1(n_462), .B2(n_501), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_276), .Y(n_901) );
INVx1_ASAP7_75t_L g487 ( .A(n_277), .Y(n_487) );
INVx1_ASAP7_75t_L g748 ( .A(n_278), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_279), .B(n_534), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1076 ( .A(n_287), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_290), .Y(n_619) );
INVx1_ASAP7_75t_L g737 ( .A(n_292), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_293), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_295), .Y(n_856) );
INVx1_ASAP7_75t_L g978 ( .A(n_296), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_297), .A2(n_320), .B1(n_589), .B2(n_780), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_298), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_299), .B(n_503), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_302), .A2(n_361), .B1(n_508), .B2(n_625), .Y(n_791) );
INVx1_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_308), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_310), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g371 ( .A(n_311), .Y(n_371) );
INVx1_ASAP7_75t_L g715 ( .A(n_312), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_314), .A2(n_321), .B1(n_548), .B2(n_551), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g936 ( .A(n_315), .Y(n_936) );
INVx1_ASAP7_75t_L g686 ( .A(n_316), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_319), .Y(n_613) );
AO22x2_ASAP7_75t_L g597 ( .A1(n_325), .A2(n_598), .B1(n_635), .B2(n_636), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_325), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_326), .Y(n_759) );
INVx1_ASAP7_75t_L g484 ( .A(n_328), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g1088 ( .A1(n_332), .A2(n_348), .B1(n_668), .B2(n_1089), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_333), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_336), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_341), .Y(n_919) );
INVx1_ASAP7_75t_L g671 ( .A(n_342), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_343), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_344), .B(n_515), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_345), .A2(n_359), .B1(n_585), .B2(n_949), .Y(n_1045) );
XOR2x2_ASAP7_75t_L g639 ( .A(n_346), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_351), .B(n_673), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_353), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_354), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_358), .Y(n_972) );
INVx1_ASAP7_75t_L g731 ( .A(n_362), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_365), .Y(n_934) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_372), .Y(n_369) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_371), .Y(n_1060) );
OA21x2_ASAP7_75t_L g1101 ( .A1(n_372), .A2(n_1059), .B(n_1102), .Y(n_1101) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_803), .B1(n_1054), .B2(n_1055), .C(n_1056), .Y(n_376) );
INVx1_ASAP7_75t_L g1054 ( .A(n_377), .Y(n_1054) );
XOR2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_693), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_557), .B2(n_692), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_475), .B1(n_555), .B2(n_556), .Y(n_380) );
INVx1_ASAP7_75t_L g555 ( .A(n_381), .Y(n_555) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_441), .Y(n_384) );
NOR3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_409), .C(n_430), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_404), .B2(n_405), .Y(n_386) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g563 ( .A(n_389), .Y(n_563) );
INVx1_ASAP7_75t_SL g957 ( .A(n_389), .Y(n_957) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_390), .Y(n_867) );
BUFx3_ASAP7_75t_L g918 ( .A(n_390), .Y(n_918) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_399), .Y(n_390) );
INVx2_ASAP7_75t_L g470 ( .A(n_391), .Y(n_470) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
AND2x2_ASAP7_75t_L g408 ( .A(n_392), .B(n_397), .Y(n_408) );
AND2x2_ASAP7_75t_L g446 ( .A(n_392), .B(n_423), .Y(n_446) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g413 ( .A(n_393), .B(n_397), .Y(n_413) );
AND2x2_ASAP7_75t_L g424 ( .A(n_393), .B(n_403), .Y(n_424) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_396), .Y(n_398) );
INVx2_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
INVx1_ASAP7_75t_L g458 ( .A(n_397), .Y(n_458) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_400), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g448 ( .A(n_400), .B(n_446), .Y(n_448) );
AND2x4_ASAP7_75t_L g505 ( .A(n_400), .B(n_470), .Y(n_505) );
AND2x6_ASAP7_75t_L g508 ( .A(n_400), .B(n_408), .Y(n_508) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_401), .Y(n_422) );
INVx1_ASAP7_75t_L g440 ( .A(n_401), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_401), .B(n_403), .Y(n_459) );
AND2x2_ASAP7_75t_L g414 ( .A(n_402), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g454 ( .A(n_403), .B(n_440), .Y(n_454) );
OA211x2_ASAP7_75t_L g670 ( .A1(n_405), .A2(n_671), .B(n_672), .C(n_674), .Y(n_670) );
OA211x2_ASAP7_75t_L g881 ( .A1(n_405), .A2(n_882), .B(n_883), .C(n_884), .Y(n_881) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g566 ( .A(n_406), .Y(n_566) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g736 ( .A(n_407), .Y(n_736) );
AND2x2_ASAP7_75t_L g453 ( .A(n_408), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g473 ( .A(n_408), .B(n_414), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_408), .B(n_454), .Y(n_486) );
OAI21xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_416), .B(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g632 ( .A(n_410), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_410), .A2(n_712), .B(n_713), .Y(n_711) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI222xp33_ASAP7_75t_L g740 ( .A1(n_411), .A2(n_741), .B1(n_745), .B2(n_746), .C1(n_747), .C2(n_748), .Y(n_740) );
INVx4_ASAP7_75t_L g758 ( .A(n_411), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g911 ( .A1(n_411), .A2(n_912), .B1(n_913), .B2(n_914), .C(n_915), .Y(n_911) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_412), .Y(n_514) );
INVx2_ASAP7_75t_L g524 ( .A(n_412), .Y(n_524) );
BUFx3_ASAP7_75t_L g798 ( .A(n_412), .Y(n_798) );
AND2x6_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g437 ( .A(n_413), .Y(n_437) );
AND2x4_ASAP7_75t_L g529 ( .A(n_413), .B(n_439), .Y(n_529) );
AND2x2_ASAP7_75t_L g445 ( .A(n_414), .B(n_446), .Y(n_445) );
AND2x6_ASAP7_75t_L g469 ( .A(n_414), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g962 ( .A(n_418), .Y(n_962) );
INVx2_ASAP7_75t_SL g995 ( .A(n_418), .Y(n_995) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx4f_ASAP7_75t_SL g536 ( .A(n_420), .Y(n_536) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_420), .Y(n_633) );
BUFx2_ASAP7_75t_L g714 ( .A(n_420), .Y(n_714) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_420), .Y(n_744) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g429 ( .A(n_422), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_423), .Y(n_434) );
AND2x4_ASAP7_75t_L g428 ( .A(n_424), .B(n_429), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_424), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g537 ( .A(n_424), .B(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx4f_ASAP7_75t_SL g515 ( .A(n_427), .Y(n_515) );
BUFx12f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_428), .Y(n_527) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_428), .Y(n_574) );
INVx1_ASAP7_75t_L g1079 ( .A(n_428), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_432), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_575) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g511 ( .A(n_433), .Y(n_511) );
INVx4_ASAP7_75t_L g909 ( .A(n_433), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_433), .A2(n_630), .B1(n_999), .B2(n_1000), .Y(n_998) );
AND2x2_ASAP7_75t_L g545 ( .A(n_434), .B(n_467), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_436), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_436), .Y(n_579) );
BUFx2_ASAP7_75t_L g630 ( .A(n_436), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_436), .A2(n_907), .B1(n_908), .B2(n_910), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_436), .A2(n_511), .B1(n_940), .B2(n_941), .Y(n_939) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_460), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
BUFx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
INVx2_ASAP7_75t_L g602 ( .A(n_445), .Y(n_602) );
BUFx2_ASAP7_75t_SL g643 ( .A(n_445), .Y(n_643) );
AND2x2_ASAP7_75t_L g464 ( .A(n_446), .B(n_454), .Y(n_464) );
AND2x4_ASAP7_75t_L g466 ( .A(n_446), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_446), .B(n_454), .Y(n_498) );
BUFx2_ASAP7_75t_L g605 ( .A(n_447), .Y(n_605) );
INVxp67_ASAP7_75t_L g857 ( .A(n_447), .Y(n_857) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g482 ( .A(n_448), .Y(n_482) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_448), .Y(n_646) );
BUFx3_ASAP7_75t_L g780 ( .A(n_448), .Y(n_780) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g591 ( .A(n_451), .Y(n_591) );
INVx5_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g669 ( .A(n_452), .Y(n_669) );
INVx4_ASAP7_75t_L g701 ( .A(n_452), .Y(n_701) );
INVx1_ASAP7_75t_L g773 ( .A(n_452), .Y(n_773) );
INVx2_ASAP7_75t_L g821 ( .A(n_452), .Y(n_821) );
INVx3_ASAP7_75t_L g835 ( .A(n_452), .Y(n_835) );
INVx8_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g592 ( .A(n_456), .Y(n_592) );
BUFx2_ASAP7_75t_L g610 ( .A(n_456), .Y(n_610) );
BUFx2_ASAP7_75t_L g648 ( .A(n_456), .Y(n_648) );
BUFx4f_ASAP7_75t_SL g975 ( .A(n_456), .Y(n_975) );
INVx6_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_457), .A2(n_484), .B1(n_485), .B2(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g898 ( .A(n_457), .Y(n_898) );
INVx1_ASAP7_75t_SL g1089 ( .A(n_457), .Y(n_1089) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g538 ( .A(n_458), .Y(n_538) );
INVx1_ASAP7_75t_L g467 ( .A(n_459), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_468), .Y(n_460) );
BUFx4f_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g548 ( .A(n_464), .Y(n_548) );
BUFx3_ASAP7_75t_L g585 ( .A(n_464), .Y(n_585) );
BUFx3_ASAP7_75t_L g770 ( .A(n_464), .Y(n_770) );
BUFx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_SL g501 ( .A(n_466), .Y(n_501) );
BUFx3_ASAP7_75t_L g551 ( .A(n_466), .Y(n_551) );
BUFx3_ASAP7_75t_L g622 ( .A(n_466), .Y(n_622) );
BUFx3_ASAP7_75t_L g657 ( .A(n_466), .Y(n_657) );
INVx1_ASAP7_75t_L g817 ( .A(n_466), .Y(n_817) );
BUFx3_ASAP7_75t_L g863 ( .A(n_466), .Y(n_863) );
BUFx2_ASAP7_75t_L g949 ( .A(n_466), .Y(n_949) );
INVx11_ASAP7_75t_L g490 ( .A(n_469), .Y(n_490) );
INVx11_ASAP7_75t_L g543 ( .A(n_469), .Y(n_543) );
INVx1_ASAP7_75t_L g687 ( .A(n_471), .Y(n_687) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g660 ( .A(n_472), .Y(n_660) );
INVx2_ASAP7_75t_L g730 ( .A(n_472), .Y(n_730) );
INVx6_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g493 ( .A(n_473), .Y(n_493) );
BUFx3_ASAP7_75t_L g550 ( .A(n_473), .Y(n_550) );
BUFx3_ASAP7_75t_L g616 ( .A(n_473), .Y(n_616) );
INVx1_ASAP7_75t_L g556 ( .A(n_475), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_518), .B1(n_553), .B2(n_554), .Y(n_475) );
INVx1_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
INVx1_ASAP7_75t_L g517 ( .A(n_477), .Y(n_517) );
AND4x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .C(n_502), .D(n_513), .Y(n_477) );
INVx1_ASAP7_75t_SL g855 ( .A(n_479), .Y(n_855) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g589 ( .A(n_480), .Y(n_589) );
INVx3_ASAP7_75t_L g721 ( .A(n_480), .Y(n_721) );
BUFx3_ASAP7_75t_L g777 ( .A(n_480), .Y(n_777) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_485), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_485), .A2(n_972), .B1(n_973), .B2(n_974), .Y(n_971) );
BUFx2_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
INVx4_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g659 ( .A(n_490), .Y(n_659) );
INVx2_ASAP7_75t_L g704 ( .A(n_490), .Y(n_704) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_490), .Y(n_833) );
INVx5_ASAP7_75t_SL g862 ( .A(n_490), .Y(n_862) );
INVx2_ASAP7_75t_SL g888 ( .A(n_490), .Y(n_888) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_499), .B2(n_500), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_496), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g679 ( .A(n_497), .Y(n_679) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_500), .A2(n_645), .B1(n_903), .B2(n_904), .Y(n_902) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g673 ( .A(n_503), .Y(n_673) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g532 ( .A(n_504), .Y(n_532) );
INVx5_ASAP7_75t_L g625 ( .A(n_504), .Y(n_625) );
INVx2_ASAP7_75t_L g1021 ( .A(n_504), .Y(n_1021) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_SL g651 ( .A(n_507), .Y(n_651) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
BUFx4f_ASAP7_75t_L g534 ( .A(n_508), .Y(n_534) );
BUFx2_ASAP7_75t_L g626 ( .A(n_508), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_511), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
INVx2_ASAP7_75t_SL g568 ( .A(n_514), .Y(n_568) );
INVx1_ASAP7_75t_L g747 ( .A(n_515), .Y(n_747) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
AO22x2_ASAP7_75t_L g783 ( .A1(n_520), .A2(n_553), .B1(n_784), .B2(n_785), .Y(n_783) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_552), .Y(n_520) );
NAND2x1_ASAP7_75t_L g521 ( .A(n_522), .B(n_539), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_530), .Y(n_522) );
OAI21xp5_ASAP7_75t_SL g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
BUFx3_ASAP7_75t_L g634 ( .A(n_527), .Y(n_634) );
BUFx2_ASAP7_75t_L g872 ( .A(n_527), .Y(n_872) );
INVx2_ASAP7_75t_L g913 ( .A(n_527), .Y(n_913) );
BUFx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g675 ( .A(n_529), .Y(n_675) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_529), .Y(n_710) );
BUFx2_ASAP7_75t_SL g823 ( .A(n_529), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .C(n_535), .Y(n_530) );
INVx1_ASAP7_75t_L g570 ( .A(n_536), .Y(n_570) );
INVx1_ASAP7_75t_L g654 ( .A(n_537), .Y(n_654) );
BUFx2_ASAP7_75t_L g709 ( .A(n_537), .Y(n_709) );
BUFx2_ASAP7_75t_L g765 ( .A(n_537), .Y(n_765) );
BUFx3_ASAP7_75t_L g793 ( .A(n_537), .Y(n_793) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .Y(n_540) );
INVx4_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_543), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
INVx3_ASAP7_75t_L g685 ( .A(n_543), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_543), .A2(n_728), .B1(n_729), .B2(n_731), .C(n_732), .Y(n_727) );
INVx4_ASAP7_75t_L g980 ( .A(n_543), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g1031 ( .A(n_548), .Y(n_1031) );
INVx1_ASAP7_75t_L g692 ( .A(n_557), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_595), .B1(n_690), .B2(n_691), .Y(n_557) );
INVx1_ASAP7_75t_L g690 ( .A(n_558), .Y(n_690) );
INVx2_ASAP7_75t_L g594 ( .A(n_559), .Y(n_594) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_580), .Y(n_559) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .C(n_575), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_563), .A2(n_734), .B1(n_735), .B2(n_737), .C(n_738), .Y(n_733) );
OAI221xp5_ASAP7_75t_SL g866 ( .A1(n_565), .A2(n_867), .B1(n_868), .B2(n_869), .C(n_870), .Y(n_866) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_571), .C(n_572), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_568), .A2(n_994), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_993) );
OAI222xp33_ASAP7_75t_L g1075 ( .A1(n_568), .A2(n_1076), .B1(n_1077), .B2(n_1078), .C1(n_1079), .C2(n_1080), .Y(n_1075) );
OAI222xp33_ASAP7_75t_L g756 ( .A1(n_570), .A2(n_757), .B1(n_759), .B2(n_760), .C1(n_761), .C2(n_762), .Y(n_756) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g761 ( .A(n_574), .Y(n_761) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g969 ( .A(n_579), .Y(n_969) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_587), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_585), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g691 ( .A(n_595), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_637), .B2(n_638), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g636 ( .A(n_598), .Y(n_636) );
AND4x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_611), .C(n_623), .D(n_631), .Y(n_598) );
NOR2xp33_ASAP7_75t_SL g599 ( .A(n_600), .B(n_606), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_600) );
INVx3_ASAP7_75t_L g1050 ( .A(n_602), .Y(n_1050) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
XOR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_662), .Y(n_638) );
NAND4xp75_ASAP7_75t_L g640 ( .A(n_641), .B(n_649), .C(n_655), .D(n_661), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_647), .Y(n_641) );
INVx4_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_L g666 ( .A(n_645), .Y(n_666) );
OAI221xp5_ASAP7_75t_SL g720 ( .A1(n_645), .A2(n_721), .B1(n_722), .B2(n_723), .C(n_724), .Y(n_720) );
INVx4_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g739 ( .A(n_654), .Y(n_739) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVxp67_ASAP7_75t_L g680 ( .A(n_657), .Y(n_680) );
XOR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_689), .Y(n_662) );
NAND4xp75_ASAP7_75t_L g663 ( .A(n_664), .B(n_670), .C(n_676), .D(n_688), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_682), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_679), .A2(n_729), .B1(n_851), .B2(n_852), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_679), .A2(n_687), .B1(n_900), .B2(n_901), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_686), .B2(n_687), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_716), .B2(n_802), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
XOR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_715), .Y(n_695) );
NOR4xp75_ASAP7_75t_L g696 ( .A(n_697), .B(n_702), .C(n_706), .D(n_711), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_698), .B(n_699), .Y(n_697) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g726 ( .A(n_701), .Y(n_726) );
NAND2x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g802 ( .A(n_716), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_750), .B1(n_800), .B2(n_801), .Y(n_716) );
INVx1_ASAP7_75t_L g800 ( .A(n_717), .Y(n_800) );
INVx1_ASAP7_75t_L g749 ( .A(n_719), .Y(n_749) );
OR4x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_727), .C(n_733), .D(n_740), .Y(n_719) );
INVx2_ASAP7_75t_L g1087 ( .A(n_721), .Y(n_1087) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_729), .A2(n_978), .B1(n_979), .B2(n_981), .Y(n_977) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_735), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_735), .A2(n_918), .B1(n_933), .B2(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g959 ( .A(n_736), .Y(n_959) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx4_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g1077 ( .A(n_744), .Y(n_1077) );
INVx1_ASAP7_75t_L g801 ( .A(n_750), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_782), .B2(n_783), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g781 ( .A(n_754), .Y(n_781) );
NAND3x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_767), .C(n_774), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_763), .Y(n_755) );
OAI21xp5_ASAP7_75t_SL g1015 ( .A1(n_757), .A2(n_1016), .B(n_1017), .Y(n_1015) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
BUFx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
XOR2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_799), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g786 ( .A(n_787), .B(n_790), .C(n_794), .D(n_797), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
AND2x2_ASAP7_75t_SL g790 ( .A(n_791), .B(n_792), .Y(n_790) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx3_ASAP7_75t_L g937 ( .A(n_798), .Y(n_937) );
INVx1_ASAP7_75t_L g1055 ( .A(n_803), .Y(n_1055) );
AOI22xp5_ASAP7_75t_SL g803 ( .A1(n_804), .A2(n_927), .B1(n_1052), .B2(n_1053), .Y(n_803) );
INVx1_ASAP7_75t_L g1052 ( .A(n_804), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_844), .B1(n_925), .B2(n_926), .Y(n_804) );
INVx1_ASAP7_75t_L g925 ( .A(n_805), .Y(n_925) );
OAI22xp5_ASAP7_75t_SL g805 ( .A1(n_806), .A2(n_824), .B1(n_841), .B2(n_843), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_808), .Y(n_842) );
XOR2x2_ASAP7_75t_L g891 ( .A(n_808), .B(n_892), .Y(n_891) );
NAND4xp75_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .C(n_818), .D(n_822), .Y(n_809) );
AND2x2_ASAP7_75t_SL g810 ( .A(n_811), .B(n_812), .Y(n_810) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx1_ASAP7_75t_L g843 ( .A(n_824), .Y(n_843) );
INVx1_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
NAND4xp75_ASAP7_75t_SL g826 ( .A(n_827), .B(n_830), .C(n_836), .D(n_839), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_834), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_SL g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVxp67_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g926 ( .A(n_844), .Y(n_926) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_875), .B1(n_923), .B2(n_924), .Y(n_845) );
INVx1_ASAP7_75t_L g924 ( .A(n_846), .Y(n_924) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_SL g874 ( .A(n_848), .Y(n_874) );
AND4x1_ASAP7_75t_L g848 ( .A(n_849), .B(n_858), .C(n_865), .D(n_871), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_853), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_856), .B2(n_857), .Y(n_853) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_864), .Y(n_858) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_867), .A2(n_959), .B1(n_991), .B2(n_992), .Y(n_990) );
INVx1_ASAP7_75t_L g923 ( .A(n_875), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_891), .B1(n_921), .B2(n_922), .Y(n_875) );
INVx3_ASAP7_75t_SL g922 ( .A(n_876), .Y(n_922) );
XOR2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_890), .Y(n_876) );
NAND4xp75_ASAP7_75t_L g877 ( .A(n_878), .B(n_881), .C(n_885), .D(n_889), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g1026 ( .A(n_888), .Y(n_1026) );
INVx1_ASAP7_75t_L g921 ( .A(n_891), .Y(n_921) );
XOR2xp5_ASAP7_75t_SL g892 ( .A(n_893), .B(n_920), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_894), .B(n_905), .Y(n_893) );
NOR3xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_899), .C(n_902), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
NOR3xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_911), .C(n_916), .Y(n_905) );
INVx3_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
INVx2_ASAP7_75t_L g967 ( .A(n_909), .Y(n_967) );
INVx1_ASAP7_75t_L g1053 ( .A(n_927), .Y(n_1053) );
XOR2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_985), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_951), .B1(n_952), .B2(n_984), .Y(n_928) );
INVx2_ASAP7_75t_SL g984 ( .A(n_929), .Y(n_984) );
XOR2x2_ASAP7_75t_L g929 ( .A(n_930), .B(n_950), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_942), .Y(n_930) );
NOR3xp33_ASAP7_75t_L g931 ( .A(n_932), .B(n_935), .C(n_939), .Y(n_931) );
OAI21xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B(n_938), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_937), .A2(n_961), .B1(n_962), .B2(n_963), .C(n_964), .Y(n_960) );
OAI21xp5_ASAP7_75t_SL g1036 ( .A1(n_937), .A2(n_1037), .B(n_1038), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g983 ( .A(n_953), .Y(n_983) );
AND3x1_ASAP7_75t_L g953 ( .A(n_954), .B(n_970), .C(n_976), .Y(n_953) );
NOR3xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_960), .C(n_965), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_957), .B1(n_958), .B2(n_959), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_965) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .B1(n_1010), .B2(n_1011), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g1009 ( .A(n_988), .Y(n_1009) );
AND2x2_ASAP7_75t_L g988 ( .A(n_989), .B(n_1001), .Y(n_988) );
NOR3xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_993), .C(n_998), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1005), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1004), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1007), .Y(n_1005) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
XNOR2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1033), .Y(n_1011) );
NAND3x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1023), .C(n_1028), .Y(n_1013) );
NOR2x1_ASAP7_75t_SL g1014 ( .A(n_1015), .B(n_1018), .Y(n_1014) );
NAND3xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .C(n_1022), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1027), .Y(n_1023) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1032), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
XOR2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1051), .Y(n_1033) );
NAND2xp5_ASAP7_75t_SL g1034 ( .A(n_1035), .B(n_1043), .Y(n_1034) );
NOR2xp33_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1039), .Y(n_1035) );
NAND3xp33_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1041), .C(n_1042), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1047), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1046), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1049), .Y(n_1047) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_1057), .Y(n_1056) );
NOR2x1_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1062), .Y(n_1057) );
OR2x2_ASAP7_75t_SL g1107 ( .A(n_1058), .B(n_1063), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1061), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_1059), .Y(n_1095) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1060), .B(n_1098), .Y(n_1102) );
CKINVDCx16_ASAP7_75t_R g1098 ( .A(n_1061), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g1062 ( .A(n_1063), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1068), .Y(n_1066) );
OAI322xp33_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1094), .A3(n_1096), .B1(n_1099), .B2(n_1103), .C1(n_1104), .C2(n_1105), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_1072), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1084), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1081), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1090), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1093), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_1101), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_1106), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g1106 ( .A(n_1107), .Y(n_1106) );
endmodule