module fake_jpeg_28433_n_274 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_21),
.B1(n_39),
.B2(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_45),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_28),
.C(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_50),
.B(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_69),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_17),
.B(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_76),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_21),
.B(n_35),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_73),
.Y(n_115)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_32),
.B1(n_36),
.B2(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_59),
.B1(n_35),
.B2(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_35),
.B1(n_37),
.B2(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_107),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_109),
.B1(n_139),
.B2(n_99),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_65),
.B1(n_62),
.B2(n_49),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_73),
.B(n_59),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_128),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_113),
.B1(n_123),
.B2(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_36),
.B1(n_29),
.B2(n_26),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_24),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_23),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_46),
.B1(n_22),
.B2(n_4),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_136),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_70),
.B(n_59),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_86),
.C(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_15),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_22),
.B(n_7),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_100),
.B1(n_98),
.B2(n_71),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_100),
.B1(n_71),
.B2(n_95),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_5),
.B(n_7),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_11),
.B(n_13),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_95),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_156),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_86),
.B(n_85),
.C(n_74),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_158),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_105),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_149),
.A2(n_159),
.B(n_132),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_105),
.B1(n_8),
.B2(n_9),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_140),
.B1(n_130),
.B2(n_109),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_110),
.B(n_16),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_85),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_161),
.B(n_162),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_110),
.B(n_8),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_10),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_10),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_135),
.B(n_117),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_11),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_13),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_14),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_130),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_144),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_177),
.B1(n_190),
.B2(n_192),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_141),
.B(n_144),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_130),
.B1(n_132),
.B2(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_135),
.Y(n_182)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_129),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_189),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_158),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_118),
.B1(n_120),
.B2(n_107),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_145),
.A2(n_120),
.B1(n_107),
.B2(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_152),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_117),
.C(n_114),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_150),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_205),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_210),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_184),
.A3(n_179),
.B1(n_177),
.B2(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_149),
.C(n_148),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_187),
.C(n_171),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_145),
.B1(n_144),
.B2(n_155),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_180),
.B1(n_190),
.B2(n_159),
.Y(n_224)
);

OA21x2_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_160),
.B(n_149),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_151),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_141),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_217),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_183),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_141),
.B1(n_146),
.B2(n_159),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_188),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_186),
.B(n_180),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_229),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_232),
.B1(n_197),
.B2(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_206),
.C(n_199),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_203),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_213),
.A2(n_165),
.B(n_187),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_233),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_192),
.B1(n_194),
.B2(n_193),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_215),
.C(n_174),
.Y(n_253)
);

BUFx12_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_212),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_204),
.B1(n_205),
.B2(n_197),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_224),
.B1(n_232),
.B2(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_226),
.C(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_222),
.C(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_253),
.C(n_239),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_219),
.B1(n_221),
.B2(n_223),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_247),
.B1(n_216),
.B2(n_209),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_220),
.C(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_244),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_173),
.C(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_161),
.C(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_236),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_260),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_257),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_234),
.B(n_246),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_258),
.A2(n_238),
.B(n_215),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_242),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_255),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_209),
.A3(n_208),
.B1(n_238),
.B2(n_191),
.C1(n_174),
.C2(n_178),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_208),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.C(n_263),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_151),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_269),
.B(n_170),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_268),
.B(n_154),
.C(n_143),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_270),
.C(n_170),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_122),
.B(n_127),
.Y(n_274)
);


endmodule