module fake_jpeg_16262_n_266 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_266);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_55),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_34),
.B1(n_23),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_56),
.B1(n_58),
.B2(n_32),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_22),
.B(n_20),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_67),
.B(n_2),
.Y(n_87)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_21),
.B1(n_23),
.B2(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_62),
.B1(n_52),
.B2(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_23),
.B1(n_21),
.B2(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_35),
.B1(n_26),
.B2(n_28),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_35),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_74),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_79),
.B(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_29),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_77),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_18),
.B(n_28),
.C(n_17),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_17),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_32),
.B(n_17),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_38),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_38),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_106),
.Y(n_109)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_100),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_107),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_57),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_125),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_46),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_127),
.B(n_79),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_33),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_32),
.B(n_4),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_3),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_114),
.C(n_112),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_96),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_102),
.B1(n_93),
.B2(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_146),
.B1(n_118),
.B2(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_96),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_160),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_147),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_101),
.C(n_80),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_155),
.C(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_153),
.B1(n_122),
.B2(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_152),
.B(n_156),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_95),
.A3(n_81),
.B1(n_80),
.B2(n_103),
.C1(n_76),
.C2(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_116),
.Y(n_153)
);

CKINVDCx11_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_76),
.C(n_106),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_97),
.B(n_83),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_98),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_110),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_113),
.B(n_123),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_184),
.B(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_129),
.B1(n_109),
.B2(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_177),
.B1(n_182),
.B2(n_108),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_139),
.B1(n_162),
.B2(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_112),
.C(n_141),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_130),
.B1(n_105),
.B2(n_84),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_180),
.A2(n_156),
.B1(n_130),
.B2(n_84),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_150),
.B(n_149),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_110),
.B(n_122),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_136),
.B(n_144),
.C(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_194),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_189),
.B1(n_198),
.B2(n_206),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_178),
.B1(n_184),
.B2(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_192),
.C(n_197),
.Y(n_211)
);

XOR2x2_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_183),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_195),
.B(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_138),
.C(n_137),
.Y(n_192)
);

OA21x2_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_15),
.B(n_16),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_183),
.B(n_16),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_172),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_137),
.B(n_78),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_25),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_3),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_86),
.C(n_33),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_175),
.C(n_185),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_108),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_169),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_25),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_181),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_200),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_5),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_199),
.B(n_202),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_165),
.B1(n_171),
.B2(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_163),
.B(n_12),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_196),
.B1(n_202),
.B2(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_227),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_196),
.B1(n_188),
.B2(n_31),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_10),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_8),
.B(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_8),
.Y(n_242)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_218),
.B1(n_214),
.B2(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_230),
.A2(n_211),
.B(n_24),
.C(n_8),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_10),
.B(n_11),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_6),
.C(n_7),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_245),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_6),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_242),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_243),
.Y(n_248)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_241),
.B(n_231),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_223),
.C(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_10),
.A3(n_11),
.B1(n_229),
.B2(n_231),
.C1(n_243),
.C2(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_255),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_245),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_252),
.B1(n_238),
.B2(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_256),
.C(n_260),
.Y(n_263)
);

OAI32xp33_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_264),
.A3(n_11),
.B1(n_238),
.B2(n_262),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_238),
.Y(n_266)
);


endmodule