module fake_jpeg_1887_n_276 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_276);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.C(n_32),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_82),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_0),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_62),
.Y(n_127)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_19),
.B(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_74),
.Y(n_109)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_27),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_85),
.B(n_111),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_50),
.B1(n_53),
.B2(n_78),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_61),
.B1(n_57),
.B2(n_81),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_25),
.B1(n_43),
.B2(n_38),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_125),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_44),
.B(n_31),
.C(n_38),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_43),
.B1(n_35),
.B2(n_30),
.Y(n_107)
);

OR2x4_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_44),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_35),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_2),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_71),
.B(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_86),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_27),
.B1(n_31),
.B2(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_14),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_144),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_134),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_75),
.B1(n_56),
.B2(n_77),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_132),
.B1(n_127),
.B2(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_3),
.C(n_7),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_7),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_99),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_8),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

BUFx4f_ASAP7_75t_SL g146 ( 
.A(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_148),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_10),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_158),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_155),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_160),
.B1(n_104),
.B2(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_156),
.B(n_157),
.Y(n_186)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_98),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_94),
.B(n_90),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_91),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_92),
.C(n_107),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_137),
.C(n_149),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_181),
.B1(n_134),
.B2(n_154),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_88),
.B1(n_119),
.B2(n_101),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_173),
.B1(n_184),
.B2(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_88),
.B1(n_119),
.B2(n_100),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_97),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_163),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_122),
.A3(n_127),
.B1(n_128),
.B2(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_91),
.B1(n_113),
.B2(n_123),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_137),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_136),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_193),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_203),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_207),
.B1(n_208),
.B2(n_146),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_136),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_202),
.C(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_152),
.B(n_149),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_144),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_205),
.C(n_142),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_198),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_173),
.B1(n_172),
.B2(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_168),
.B1(n_150),
.B2(n_157),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_152),
.Y(n_202)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_152),
.B1(n_147),
.B2(n_113),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_165),
.A2(n_187),
.B1(n_163),
.B2(n_167),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_220),
.B1(n_189),
.B2(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_168),
.B1(n_176),
.B2(n_170),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_219),
.B1(n_146),
.B2(n_140),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_183),
.B(n_169),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_226),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_179),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.C(n_188),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_188),
.A2(n_169),
.B(n_145),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_231),
.C(n_236),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_211),
.C(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_233),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_235),
.B1(n_239),
.B2(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_205),
.C(n_202),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_193),
.B1(n_206),
.B2(n_204),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_148),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_219),
.B1(n_218),
.B2(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_247),
.B1(n_250),
.B2(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

BUFx12_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_224),
.B1(n_221),
.B2(n_222),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_259),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_231),
.B1(n_237),
.B2(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_253),
.B(n_255),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_237),
.B(n_221),
.Y(n_254)
);

OAI31xp33_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_241),
.A3(n_247),
.B(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_229),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_236),
.C(n_222),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_248),
.B(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_248),
.C(n_242),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_252),
.B(n_257),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_268),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_245),
.B(n_258),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_141),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_258),
.B1(n_245),
.B2(n_235),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_226),
.B1(n_156),
.B2(n_123),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_271),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_270),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_265),
.B1(n_269),
.B2(n_190),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_273),
.Y(n_276)
);


endmodule