module fake_aes_9288_n_680 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_680);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_680;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_76), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_16), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_9), .Y(n_84) );
INVxp33_ASAP7_75t_L g85 ( .A(n_6), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_1), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_40), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_74), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_28), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_4), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_50), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_43), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_33), .Y(n_97) );
BUFx2_ASAP7_75t_SL g98 ( .A(n_41), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
BUFx2_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_34), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_4), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_2), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_35), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_10), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_65), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_30), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_8), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_6), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_58), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_39), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_27), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_56), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_59), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_37), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
INVx4_ASAP7_75t_R g121 ( .A(n_61), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_52), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_66), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_95), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_95), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_117), .B(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
BUFx8_ASAP7_75t_L g128 ( .A(n_117), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_95), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_100), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_95), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_93), .B(n_0), .Y(n_136) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_87), .A2(n_29), .B(n_77), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_100), .B(n_1), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_80), .B(n_2), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_85), .B(n_3), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_112), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_80), .B(n_120), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_81), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_120), .B(n_3), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_108), .B(n_5), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
BUFx8_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
AND3x2_ASAP7_75t_L g153 ( .A(n_103), .B(n_5), .C(n_7), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_94), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_118), .B(n_8), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_91), .Y(n_158) );
BUFx8_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_97), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_144), .B(n_122), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
AND3x1_ASAP7_75t_L g167 ( .A(n_136), .B(n_97), .C(n_122), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_131), .A2(n_161), .B1(n_128), .B2(n_159), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_128), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_131), .B(n_110), .Y(n_171) );
INVx6_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_151), .B(n_159), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_128), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_144), .B(n_119), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_161), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
OAI221xp5_ASAP7_75t_L g179 ( .A1(n_139), .A2(n_106), .B1(n_102), .B2(n_86), .C(n_110), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_158), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_128), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_151), .B(n_91), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_160), .B(n_119), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_151), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_127), .B(n_109), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_139), .A2(n_98), .B1(n_82), .B2(n_104), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_127), .B(n_123), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_159), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_132), .B(n_116), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_132), .B(n_116), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_145), .Y(n_200) );
NAND3x1_ASAP7_75t_L g201 ( .A(n_149), .B(n_83), .C(n_115), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_146), .B(n_107), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_142), .B(n_105), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_140), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_146), .B(n_101), .Y(n_208) );
OR2x6_ASAP7_75t_L g209 ( .A(n_191), .B(n_126), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_194), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_200), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_177), .Y(n_212) );
INVx6_ASAP7_75t_L g213 ( .A(n_200), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_204), .B(n_142), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_194), .Y(n_215) );
INVx5_ASAP7_75t_L g216 ( .A(n_200), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_164), .B(n_126), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_171), .B(n_156), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_196), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_168), .A2(n_156), .B1(n_141), .B2(n_154), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_172), .B(n_154), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_162), .Y(n_222) );
NOR2x1p5_ASAP7_75t_L g223 ( .A(n_169), .B(n_141), .Y(n_223) );
BUFx4f_ASAP7_75t_L g224 ( .A(n_191), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_164), .B(n_153), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_163), .B(n_145), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_162), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_187), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_165), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_195), .B(n_160), .Y(n_233) );
INVxp67_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_188), .B(n_145), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_172), .A2(n_148), .B1(n_155), .B2(n_152), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_166), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_183), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_165), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_197), .B(n_148), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_205), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_186), .B(n_148), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_167), .A2(n_148), .B1(n_155), .B2(n_152), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_203), .A2(n_157), .B1(n_155), .B2(n_152), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_192), .Y(n_250) );
AOI22xp5_ASAP7_75t_SL g251 ( .A1(n_183), .A2(n_92), .B1(n_101), .B2(n_98), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_172), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_172), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_164), .B(n_153), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_187), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_169), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_193), .B(n_92), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_180), .Y(n_258) );
BUFx4f_ASAP7_75t_SL g259 ( .A(n_173), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_190), .B(n_157), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_176), .B(n_137), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_176), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_170), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_186), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_203), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_216), .B(n_186), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_266), .A2(n_174), .B1(n_201), .B2(n_179), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_223), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_217), .A2(n_176), .B1(n_190), .B2(n_202), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_217), .A2(n_190), .B1(n_202), .B2(n_157), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_264), .Y(n_272) );
NAND3xp33_ASAP7_75t_SL g273 ( .A(n_240), .B(n_174), .C(n_181), .Y(n_273) );
BUFx4f_ASAP7_75t_L g274 ( .A(n_225), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_263), .A2(n_192), .B(n_99), .C(n_111), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_223), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_217), .A2(n_202), .B1(n_150), .B2(n_134), .Y(n_278) );
CKINVDCx11_ASAP7_75t_R g279 ( .A(n_209), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_212), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_261), .A2(n_185), .B(n_208), .Y(n_281) );
BUFx12f_ASAP7_75t_L g282 ( .A(n_240), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_224), .B(n_135), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_216), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_227), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
INVx5_ASAP7_75t_L g287 ( .A(n_210), .Y(n_287) );
OAI22x1_ASAP7_75t_L g288 ( .A1(n_234), .A2(n_201), .B1(n_88), .B2(n_114), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_217), .A2(n_189), .B1(n_134), .B2(n_150), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_263), .A2(n_150), .B1(n_134), .B2(n_143), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_209), .A2(n_135), .B1(n_138), .B2(n_113), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_244), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_210), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_214), .B(n_138), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_209), .A2(n_138), .B1(n_135), .B2(n_143), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_214), .B(n_138), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_261), .A2(n_137), .B(n_198), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_218), .B(n_135), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_209), .B(n_137), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_209), .B(n_9), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_220), .B(n_10), .Y(n_303) );
INVx4_ASAP7_75t_L g304 ( .A(n_216), .Y(n_304) );
OR2x6_ASAP7_75t_L g305 ( .A(n_225), .B(n_143), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_258), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_229), .Y(n_308) );
CKINVDCx16_ASAP7_75t_R g309 ( .A(n_251), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_216), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_216), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
AO31x2_ASAP7_75t_L g313 ( .A1(n_260), .A2(n_129), .A3(n_130), .B(n_124), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_258), .Y(n_314) );
BUFx2_ASAP7_75t_SL g315 ( .A(n_256), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_225), .B(n_143), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
INVx5_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_271), .A2(n_249), .B1(n_262), .B2(n_224), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_277), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_302), .A2(n_279), .B1(n_280), .B2(n_303), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_271), .B(n_249), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_315), .B(n_233), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_277), .Y(n_326) );
OAI211xp5_ASAP7_75t_L g327 ( .A1(n_268), .A2(n_279), .B(n_247), .C(n_303), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_294), .B(n_247), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_309), .A2(n_251), .B1(n_224), .B2(n_259), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
OAI22xp5_ASAP7_75t_SL g331 ( .A1(n_302), .A2(n_225), .B1(n_254), .B2(n_265), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_274), .B(n_237), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_306), .B(n_265), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_296), .A2(n_237), .B1(n_221), .B2(n_254), .C(n_238), .Y(n_336) );
AOI21xp33_ASAP7_75t_L g337 ( .A1(n_270), .A2(n_254), .B(n_262), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_273), .B(n_254), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_285), .Y(n_340) );
BUFx12f_ASAP7_75t_L g341 ( .A(n_282), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_298), .B(n_226), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_311), .B(n_232), .Y(n_344) );
INVx3_ASAP7_75t_SL g345 ( .A(n_305), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_310), .B(n_232), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_291), .Y(n_347) );
OR2x6_ASAP7_75t_L g348 ( .A(n_283), .B(n_261), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_274), .A2(n_226), .B1(n_232), .B2(n_235), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_286), .Y(n_350) );
NAND3xp33_ASAP7_75t_SL g351 ( .A(n_283), .B(n_257), .C(n_215), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_299), .A2(n_242), .B(n_219), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_352), .A2(n_292), .B(n_281), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_332), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_323), .A2(n_288), .B1(n_300), .B2(n_290), .C(n_293), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_332), .B(n_272), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_341), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_325), .A2(n_282), .B1(n_215), .B2(n_297), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_324), .B(n_289), .Y(n_360) );
AO21x2_ASAP7_75t_L g361 ( .A1(n_352), .A2(n_301), .B(n_275), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_331), .A2(n_320), .B1(n_329), .B2(n_334), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_348), .A2(n_261), .B(n_301), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_331), .A2(n_276), .B1(n_269), .B2(n_267), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_333), .A2(n_316), .B1(n_305), .B2(n_310), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_322), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_334), .A2(n_267), .B1(n_301), .B2(n_278), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_337), .A2(n_278), .B1(n_275), .B2(n_239), .C(n_252), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_328), .B(n_291), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_340), .B(n_308), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_327), .A2(n_239), .B1(n_253), .B2(n_252), .C(n_219), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_318), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_345), .A2(n_316), .B1(n_305), .B2(n_230), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_347), .B(n_326), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_348), .A2(n_316), .B1(n_308), .B2(n_292), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_326), .B(n_335), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_338), .A2(n_226), .B1(n_314), .B2(n_312), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_379), .B(n_335), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_355), .B(n_348), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_366), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_366), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_355), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_362), .A2(n_356), .B1(n_377), .B2(n_359), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_377), .A2(n_351), .B1(n_346), .B2(n_336), .Y(n_387) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_363), .A2(n_348), .B1(n_318), .B2(n_342), .C1(n_330), .C2(n_339), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_366), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_369), .B(n_348), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_369), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_346), .B1(n_345), .B2(n_343), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_371), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_346), .B1(n_345), .B2(n_344), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_379), .B(n_371), .C(n_378), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_368), .B(n_143), .C(n_318), .Y(n_397) );
OAI33xp33_ASAP7_75t_L g398 ( .A1(n_378), .A2(n_124), .A3(n_129), .B1(n_125), .B2(n_130), .B3(n_317), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_370), .A2(n_318), .B1(n_330), .B2(n_339), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_361), .A2(n_124), .B(n_130), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_376), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_358), .B(n_341), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_360), .A2(n_349), .B1(n_330), .B2(n_339), .C(n_342), .Y(n_403) );
AOI33xp33_ASAP7_75t_L g404 ( .A1(n_357), .A2(n_129), .A3(n_125), .B1(n_253), .B2(n_346), .B3(n_344), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_374), .B(n_318), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_360), .A2(n_344), .B1(n_342), .B2(n_307), .C(n_350), .Y(n_407) );
OAI31xp33_ASAP7_75t_L g408 ( .A1(n_365), .A2(n_344), .A3(n_321), .B(n_319), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_357), .B(n_321), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_373), .A2(n_321), .B1(n_318), .B2(n_319), .C(n_286), .Y(n_411) );
OAI33xp33_ASAP7_75t_L g412 ( .A1(n_370), .A2(n_372), .A3(n_375), .B1(n_125), .B2(n_14), .B3(n_15), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_405), .B(n_361), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_394), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_380), .B1(n_372), .B2(n_374), .C(n_350), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g418 ( .A1(n_396), .A2(n_374), .A3(n_350), .B(n_255), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_412), .B(n_354), .C(n_198), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_361), .B1(n_354), .B2(n_226), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_401), .B(n_313), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
AND2x4_ASAP7_75t_SL g424 ( .A(n_406), .B(n_295), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_409), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_405), .B(n_313), .Y(n_426) );
INVx4_ASAP7_75t_L g427 ( .A(n_406), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_405), .B(n_313), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_384), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_390), .B(n_313), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_399), .A2(n_295), .B(n_287), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_390), .B(n_11), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_390), .B(n_11), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_410), .B(n_12), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_410), .B(n_13), .Y(n_437) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_397), .A2(n_246), .B(n_248), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_412), .A2(n_198), .B1(n_175), .B2(n_182), .C(n_207), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_385), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_384), .B(n_14), .Y(n_441) );
INVx5_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_399), .B(n_207), .C(n_206), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_381), .B(n_16), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_389), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_396), .A2(n_175), .B1(n_182), .B2(n_206), .C(n_207), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_381), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_401), .B(n_17), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_409), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_389), .B(n_17), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_385), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_389), .B(n_18), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_18), .Y(n_454) );
OAI211xp5_ASAP7_75t_L g455 ( .A1(n_408), .A2(n_287), .B(n_133), .C(n_255), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_408), .B(n_235), .C(n_232), .D(n_241), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_448), .B(n_402), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_440), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_440), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_452), .B(n_391), .Y(n_460) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_443), .B(n_445), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_452), .B(n_415), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_415), .B(n_391), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_417), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_445), .B(n_393), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_436), .B(n_382), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_436), .B(n_382), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_428), .Y(n_469) );
INVx3_ASAP7_75t_SL g470 ( .A(n_442), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_427), .B(n_393), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g472 ( .A(n_437), .B(n_395), .C(n_392), .D(n_407), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_425), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_427), .B(n_409), .Y(n_474) );
NAND4xp75_ASAP7_75t_L g475 ( .A(n_437), .B(n_407), .C(n_393), .D(n_388), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_427), .B(n_403), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_434), .B(n_404), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_434), .B(n_400), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_435), .B(n_403), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_416), .A2(n_411), .B1(n_397), .B2(n_398), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_454), .Y(n_482) );
NOR3xp33_ASAP7_75t_SL g483 ( .A(n_455), .B(n_388), .C(n_411), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_454), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_435), .B(n_400), .Y(n_485) );
OR2x6_ASAP7_75t_L g486 ( .A(n_427), .B(n_400), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_441), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_449), .A2(n_398), .A3(n_400), .B1(n_133), .B2(n_121), .B3(n_25), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_429), .B(n_287), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_441), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_429), .B(n_295), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_429), .B(n_295), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_449), .B(n_287), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_442), .B(n_20), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_442), .B(n_21), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_451), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_453), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_432), .B(n_23), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_432), .B(n_207), .Y(n_501) );
AOI31xp67_ASAP7_75t_SL g502 ( .A1(n_421), .A2(n_24), .A3(n_26), .B(n_31), .Y(n_502) );
OR2x4_ASAP7_75t_L g503 ( .A(n_421), .B(n_175), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_431), .B(n_32), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_426), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_426), .B(n_430), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_430), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_414), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_446), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_416), .B(n_235), .C(n_241), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_443), .A2(n_230), .B(n_210), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_442), .B(n_36), .Y(n_512) );
INVx3_ASAP7_75t_SL g513 ( .A(n_442), .Y(n_513) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_485), .A2(n_447), .B(n_433), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_458), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_506), .B(n_422), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_495), .B(n_442), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_506), .B(n_422), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_470), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_509), .Y(n_521) );
AOI211xp5_ASAP7_75t_L g522 ( .A1(n_513), .A2(n_418), .B(n_433), .C(n_439), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_473), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_461), .A2(n_439), .B(n_418), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_505), .B(n_422), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_463), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_472), .A2(n_419), .B1(n_442), .B2(n_420), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_457), .B(n_450), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_475), .A2(n_472), .B1(n_477), .B2(n_480), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_507), .B(n_413), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_466), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_474), .B(n_425), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_462), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_464), .B(n_413), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_467), .B(n_450), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_468), .B(n_444), .Y(n_538) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_486), .B(n_438), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_465), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_469), .B(n_444), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_499), .B(n_424), .Y(n_542) );
NOR2xp67_ASAP7_75t_SL g543 ( .A(n_504), .B(n_456), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_478), .Y(n_544) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_463), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_483), .B(n_447), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_460), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_482), .B(n_444), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_484), .B(n_423), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_487), .A2(n_456), .B1(n_423), .B2(n_414), .C(n_206), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_460), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_479), .B(n_423), .Y(n_553) );
OAI21xp33_ASAP7_75t_L g554 ( .A1(n_476), .A2(n_414), .B(n_424), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_474), .B(n_424), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_490), .B(n_438), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_486), .B(n_38), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_508), .Y(n_558) );
XNOR2x2_ASAP7_75t_SL g559 ( .A(n_503), .B(n_438), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_492), .B(n_438), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_497), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_498), .B(n_42), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_500), .B(n_45), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_494), .Y(n_565) );
XOR2x2_ASAP7_75t_L g566 ( .A(n_496), .B(n_46), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_489), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_486), .B(n_206), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_488), .B(n_235), .C(n_241), .Y(n_569) );
XNOR2x2_ASAP7_75t_L g570 ( .A(n_512), .B(n_49), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_553), .B(n_481), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_525), .Y(n_572) );
NAND2xp33_ASAP7_75t_SL g573 ( .A(n_543), .B(n_502), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_537), .B(n_493), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_516), .B(n_491), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_528), .B(n_510), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_535), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_534), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_555), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_518), .B(n_133), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_546), .A2(n_511), .B(n_133), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_531), .B(n_51), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_533), .B(n_206), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_515), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_519), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_540), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_545), .B(n_133), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_526), .B(n_133), .Y(n_589) );
XNOR2x1_ASAP7_75t_L g590 ( .A(n_566), .B(n_53), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_565), .B(n_54), .Y(n_591) );
NOR2x1p5_ASAP7_75t_L g592 ( .A(n_557), .B(n_207), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_560), .B(n_182), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_548), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_532), .B(n_182), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_532), .B(n_182), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_547), .B(n_175), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_567), .B(n_55), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_552), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_561), .B(n_175), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_538), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_564), .B(n_57), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_520), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_549), .Y(n_606) );
NOR2xp67_ASAP7_75t_L g607 ( .A(n_524), .B(n_60), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_536), .B(n_64), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_551), .A2(n_210), .B1(n_241), .B2(n_211), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_551), .A2(n_522), .B1(n_529), .B2(n_524), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_550), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_550), .Y(n_613) );
NAND2xp33_ASAP7_75t_SL g614 ( .A(n_557), .B(n_210), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_568), .B(n_211), .C(n_248), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g616 ( .A(n_559), .B(n_67), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_534), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_527), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_523), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_523), .B(n_68), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_554), .B(n_69), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_558), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_559), .A2(n_250), .B(n_246), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_541), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_536), .B(n_70), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_539), .B(n_73), .Y(n_626) );
INVx2_ASAP7_75t_SL g627 ( .A(n_517), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_541), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_556), .B(n_78), .Y(n_629) );
XOR2xp5_ASAP7_75t_L g630 ( .A(n_570), .B(n_250), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_517), .B(n_228), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_556), .B(n_226), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_562), .B(n_226), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_563), .A2(n_226), .B1(n_245), .B2(n_222), .C1(n_228), .C2(n_231), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_542), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_514), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_569), .A2(n_514), .B1(n_236), .B2(n_222), .C(n_231), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_531), .B(n_236), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_546), .A2(n_243), .B(n_245), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_525), .Y(n_640) );
XOR2xp5_ASAP7_75t_L g641 ( .A(n_590), .B(n_599), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_571), .B(n_636), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_624), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_605), .A2(n_578), .B1(n_617), .B2(n_579), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_611), .A2(n_583), .B(n_580), .C(n_619), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_573), .A2(n_571), .B1(n_583), .B2(n_576), .Y(n_646) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_592), .B(n_607), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_573), .A2(n_635), .B1(n_603), .B2(n_638), .Y(n_648) );
NOR2xp33_ASAP7_75t_R g649 ( .A(n_614), .B(n_616), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_630), .A2(n_594), .B(n_638), .C(n_619), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_617), .A2(n_590), .B1(n_612), .B2(n_610), .C(n_606), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_613), .B(n_628), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_627), .A2(n_575), .B1(n_626), .B2(n_618), .Y(n_653) );
AND4x1_ASAP7_75t_L g654 ( .A(n_621), .B(n_591), .C(n_637), .D(n_615), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_640), .A2(n_577), .B1(n_572), .B2(n_595), .C(n_586), .Y(n_655) );
OR3x1_ASAP7_75t_L g656 ( .A(n_621), .B(n_591), .C(n_601), .Y(n_656) );
AO22x2_ASAP7_75t_L g657 ( .A1(n_644), .A2(n_587), .B1(n_585), .B2(n_600), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g658 ( .A(n_641), .B(n_574), .Y(n_658) );
AOI221x1_ASAP7_75t_L g659 ( .A1(n_653), .A2(n_588), .B1(n_608), .B2(n_625), .C(n_623), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g660 ( .A(n_649), .B(n_626), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_646), .A2(n_648), .B(n_645), .C(n_650), .Y(n_661) );
AOI322xp5_ASAP7_75t_L g662 ( .A1(n_642), .A2(n_574), .A3(n_581), .B1(n_596), .B2(n_597), .C1(n_622), .C2(n_620), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_651), .A2(n_582), .B(n_634), .C(n_584), .Y(n_663) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_643), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g665 ( .A1(n_655), .A2(n_581), .A3(n_597), .B1(n_596), .B2(n_622), .C1(n_593), .C2(n_589), .Y(n_665) );
NAND3xp33_ASAP7_75t_SL g666 ( .A(n_661), .B(n_654), .C(n_656), .Y(n_666) );
NOR4xp25_ASAP7_75t_L g667 ( .A(n_663), .B(n_652), .C(n_604), .D(n_602), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_657), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_660), .A2(n_647), .B1(n_632), .B2(n_633), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_664), .A2(n_609), .B1(n_593), .B2(n_589), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_666), .B(n_598), .C(n_629), .Y(n_671) );
XOR2xp5_ASAP7_75t_L g672 ( .A(n_670), .B(n_658), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_667), .A2(n_665), .B1(n_662), .B2(n_664), .C(n_659), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_673), .A2(n_668), .B1(n_669), .B2(n_631), .C(n_639), .Y(n_674) );
NAND3x1_ASAP7_75t_L g675 ( .A(n_672), .B(n_602), .C(n_213), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_675), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_676), .A2(n_671), .B(n_199), .C(n_243), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_678), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_679), .A2(n_677), .B(n_199), .Y(n_680) );
endmodule