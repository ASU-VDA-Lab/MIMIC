module fake_netlist_5_1044_n_4411 (n_137, n_924, n_676, n_294, n_431, n_318, n_380, n_419, n_977, n_653, n_611, n_444, n_642, n_469, n_615, n_851, n_82, n_194, n_316, n_785, n_389, n_843, n_855, n_549, n_684, n_850, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_865, n_61, n_913, n_678, n_664, n_376, n_697, n_503, n_967, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_928, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_916, n_452, n_885, n_397, n_493, n_111, n_525, n_880, n_703, n_698, n_980, n_483, n_544, n_683, n_1007, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_998, n_116, n_841, n_956, n_22, n_467, n_564, n_802, n_423, n_840, n_284, n_46, n_245, n_21, n_501, n_823, n_725, n_983, n_139, n_38, n_105, n_280, n_744, n_1021, n_590, n_629, n_672, n_4, n_873, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_898, n_254, n_690, n_33, n_1013, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_1022, n_526, n_915, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_859, n_864, n_951, n_821, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_909, n_625, n_854, n_949, n_621, n_753, n_997, n_100, n_455, n_674, n_1008, n_932, n_417, n_946, n_612, n_1001, n_212, n_385, n_498, n_516, n_933, n_788, n_507, n_119, n_497, n_689, n_738, n_912, n_606, n_559, n_275, n_640, n_968, n_252, n_624, n_825, n_26, n_295, n_133, n_1010, n_330, n_877, n_508, n_739, n_506, n_2, n_737, n_610, n_972, n_692, n_986, n_755, n_6, n_509, n_568, n_936, n_39, n_147, n_373, n_820, n_757, n_947, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_999, n_668, n_733, n_991, n_375, n_301, n_828, n_779, n_576, n_941, n_929, n_981, n_68, n_804, n_93, n_867, n_186, n_537, n_134, n_902, n_191, n_587, n_945, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_878, n_524, n_943, n_399, n_341, n_204, n_394, n_250, n_579, n_992, n_938, n_741, n_548, n_543, n_260, n_812, n_842, n_298, n_650, n_984, n_320, n_694, n_518, n_505, n_286, n_883, n_122, n_282, n_752, n_331, n_10, n_905, n_906, n_24, n_406, n_519, n_470, n_908, n_782, n_919, n_325, n_449, n_132, n_862, n_90, n_900, n_724, n_856, n_546, n_1016, n_101, n_760, n_658, n_281, n_918, n_240, n_942, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_959, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_940, n_896, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_920, n_894, n_271, n_934, n_1017, n_94, n_831, n_826, n_335, n_123, n_886, n_978, n_964, n_654, n_370, n_167, n_976, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_833, n_297, n_156, n_5, n_853, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_988, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_1009, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_961, n_995, n_955, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_882, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_897, n_215, n_350, n_196, n_798, n_662, n_459, n_1020, n_646, n_211, n_218, n_400, n_930, n_181, n_436, n_962, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_994, n_926, n_287, n_344, n_848, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_958, n_849, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_922, n_145, n_48, n_521, n_614, n_663, n_845, n_50, n_337, n_430, n_313, n_631, n_673, n_837, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_974, n_395, n_164, n_432, n_553, n_727, n_839, n_901, n_311, n_813, n_957, n_830, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_888, n_296, n_613, n_871, n_241, n_637, n_357, n_875, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_829, n_144, n_858, n_114, n_96, n_923, n_772, n_691, n_881, n_717, n_165, n_468, n_499, n_939, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_866, n_969, n_236, n_388, n_761, n_1012, n_1, n_1019, n_249, n_903, n_1006, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_889, n_80, n_973, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_836, n_990, n_84, n_462, n_975, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_907, n_722, n_458, n_288, n_770, n_188, n_190, n_844, n_201, n_263, n_471, n_609, n_852, n_989, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_834, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_892, n_893, n_1015, n_1000, n_891, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_979, n_1002, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_846, n_874, n_465, n_838, n_76, n_358, n_362, n_876, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_953, n_601, n_279, n_917, n_1014, n_966, n_70, n_987, n_253, n_261, n_174, n_289, n_745, n_963, n_954, n_627, n_767, n_172, n_206, n_217, n_993, n_440, n_726, n_478, n_793, n_545, n_982, n_441, n_860, n_450, n_648, n_312, n_476, n_818, n_429, n_861, n_534, n_948, n_884, n_899, n_345, n_210, n_944, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_970, n_911, n_557, n_182, n_143, n_83, n_1005, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_832, n_180, n_857, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_937, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_879, n_16, n_720, n_0, n_58, n_623, n_405, n_824, n_18, n_359, n_863, n_910, n_971, n_490, n_805, n_117, n_326, n_794, n_768, n_921, n_996, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_847, n_815, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_822, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_895, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_887, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_870, n_931, n_159, n_334, n_599, n_766, n_811, n_952, n_541, n_807, n_391, n_701, n_434, n_1023, n_645, n_539, n_835, n_175, n_538, n_666, n_262, n_803, n_868, n_238, n_639, n_799, n_914, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_965, n_927, n_20, n_536, n_531, n_935, n_1004, n_121, n_242, n_817, n_872, n_360, n_36, n_594, n_764, n_200, n_890, n_162, n_960, n_64, n_759, n_1018, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_1011, n_904, n_985, n_869, n_324, n_810, n_634, n_416, n_199, n_827, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_925, n_424, n_1003, n_7, n_706, n_746, n_256, n_305, n_533, n_950, n_747, n_52, n_278, n_784, n_110, n_4411);

input n_137;
input n_924;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_977;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_851;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_843;
input n_855;
input n_549;
input n_684;
input n_850;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_865;
input n_61;
input n_913;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_967;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_928;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_916;
input n_452;
input n_885;
input n_397;
input n_493;
input n_111;
input n_525;
input n_880;
input n_703;
input n_698;
input n_980;
input n_483;
input n_544;
input n_683;
input n_1007;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_998;
input n_116;
input n_841;
input n_956;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_840;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_823;
input n_725;
input n_983;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_1021;
input n_590;
input n_629;
input n_672;
input n_4;
input n_873;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_898;
input n_254;
input n_690;
input n_33;
input n_1013;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_1022;
input n_526;
input n_915;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_859;
input n_864;
input n_951;
input n_821;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_909;
input n_625;
input n_854;
input n_949;
input n_621;
input n_753;
input n_997;
input n_100;
input n_455;
input n_674;
input n_1008;
input n_932;
input n_417;
input n_946;
input n_612;
input n_1001;
input n_212;
input n_385;
input n_498;
input n_516;
input n_933;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_912;
input n_606;
input n_559;
input n_275;
input n_640;
input n_968;
input n_252;
input n_624;
input n_825;
input n_26;
input n_295;
input n_133;
input n_1010;
input n_330;
input n_877;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_972;
input n_692;
input n_986;
input n_755;
input n_6;
input n_509;
input n_568;
input n_936;
input n_39;
input n_147;
input n_373;
input n_820;
input n_757;
input n_947;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_999;
input n_668;
input n_733;
input n_991;
input n_375;
input n_301;
input n_828;
input n_779;
input n_576;
input n_941;
input n_929;
input n_981;
input n_68;
input n_804;
input n_93;
input n_867;
input n_186;
input n_537;
input n_134;
input n_902;
input n_191;
input n_587;
input n_945;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_878;
input n_524;
input n_943;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_992;
input n_938;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_842;
input n_298;
input n_650;
input n_984;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_883;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_905;
input n_906;
input n_24;
input n_406;
input n_519;
input n_470;
input n_908;
input n_782;
input n_919;
input n_325;
input n_449;
input n_132;
input n_862;
input n_90;
input n_900;
input n_724;
input n_856;
input n_546;
input n_1016;
input n_101;
input n_760;
input n_658;
input n_281;
input n_918;
input n_240;
input n_942;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_959;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_940;
input n_896;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_920;
input n_894;
input n_271;
input n_934;
input n_1017;
input n_94;
input n_831;
input n_826;
input n_335;
input n_123;
input n_886;
input n_978;
input n_964;
input n_654;
input n_370;
input n_167;
input n_976;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_833;
input n_297;
input n_156;
input n_5;
input n_853;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_988;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_1009;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_961;
input n_995;
input n_955;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_882;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_1020;
input n_646;
input n_211;
input n_218;
input n_400;
input n_930;
input n_181;
input n_436;
input n_962;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_994;
input n_926;
input n_287;
input n_344;
input n_848;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_958;
input n_849;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_922;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_845;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_837;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_974;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_839;
input n_901;
input n_311;
input n_813;
input n_957;
input n_830;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_888;
input n_296;
input n_613;
input n_871;
input n_241;
input n_637;
input n_357;
input n_875;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_829;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_772;
input n_691;
input n_881;
input n_717;
input n_165;
input n_468;
input n_499;
input n_939;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_866;
input n_969;
input n_236;
input n_388;
input n_761;
input n_1012;
input n_1;
input n_1019;
input n_249;
input n_903;
input n_1006;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_889;
input n_80;
input n_973;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_836;
input n_990;
input n_84;
input n_462;
input n_975;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_907;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_844;
input n_201;
input n_263;
input n_471;
input n_609;
input n_852;
input n_989;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_834;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_892;
input n_893;
input n_1015;
input n_1000;
input n_891;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_979;
input n_1002;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_846;
input n_874;
input n_465;
input n_838;
input n_76;
input n_358;
input n_362;
input n_876;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_953;
input n_601;
input n_279;
input n_917;
input n_1014;
input n_966;
input n_70;
input n_987;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_963;
input n_954;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_993;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_982;
input n_441;
input n_860;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_861;
input n_534;
input n_948;
input n_884;
input n_899;
input n_345;
input n_210;
input n_944;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_970;
input n_911;
input n_557;
input n_182;
input n_143;
input n_83;
input n_1005;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_832;
input n_180;
input n_857;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_937;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_879;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_824;
input n_18;
input n_359;
input n_863;
input n_910;
input n_971;
input n_490;
input n_805;
input n_117;
input n_326;
input n_794;
input n_768;
input n_921;
input n_996;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_847;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_822;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_895;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_887;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_870;
input n_931;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_952;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_1023;
input n_645;
input n_539;
input n_835;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_868;
input n_238;
input n_639;
input n_799;
input n_914;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_965;
input n_927;
input n_20;
input n_536;
input n_531;
input n_935;
input n_1004;
input n_121;
input n_242;
input n_817;
input n_872;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_890;
input n_162;
input n_960;
input n_64;
input n_759;
input n_1018;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_1011;
input n_904;
input n_985;
input n_869;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_827;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_925;
input n_424;
input n_1003;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_950;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_4411;

wire n_1263;
wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_2380;
wire n_1166;
wire n_1751;
wire n_2771;
wire n_1508;
wire n_3241;
wire n_4129;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_2899;
wire n_2955;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4127;
wire n_4138;
wire n_3086;
wire n_3297;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_4217;
wire n_4395;
wire n_2683;
wire n_2347;
wire n_1292;
wire n_2520;
wire n_2821;
wire n_1370;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_2487;
wire n_1466;
wire n_1695;
wire n_3766;
wire n_1353;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_3813;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4238;
wire n_1451;
wire n_4109;
wire n_2302;
wire n_4038;
wire n_1545;
wire n_2374;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1462;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_4013;
wire n_2011;
wire n_2096;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_2483;
wire n_1696;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_4155;
wire n_1359;
wire n_3695;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_3036;
wire n_3891;
wire n_2482;
wire n_1728;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4061;
wire n_4131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_4315;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1633;
wire n_1236;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_2466;
wire n_2091;
wire n_2652;
wire n_1289;
wire n_2635;
wire n_1517;
wire n_4311;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_1484;
wire n_2071;
wire n_2643;
wire n_2561;
wire n_1328;
wire n_1374;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_3049;
wire n_1598;
wire n_4394;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1547;
wire n_1070;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1071;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_3985;
wire n_1801;
wire n_1391;
wire n_1034;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_3744;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_3980;
wire n_2915;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_1587;
wire n_2682;
wire n_1473;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_4258;
wire n_1521;
wire n_1284;
wire n_1744;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2506;
wire n_2699;
wire n_4064;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3550;
wire n_2615;
wire n_3940;
wire n_1556;
wire n_1384;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_2118;
wire n_2985;
wire n_1151;
wire n_2944;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_2358;
wire n_3986;
wire n_4376;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_3837;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_3915;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_4385;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_1058;
wire n_1667;
wire n_3359;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_4405;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4375;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_1052;
wire n_3781;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_2987;
wire n_2042;
wire n_1527;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_3328;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_3433;
wire n_4024;
wire n_3392;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_2305;
wire n_3430;
wire n_3975;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_4151;
wire n_4148;
wire n_1906;
wire n_1883;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_1156;
wire n_4331;
wire n_4160;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_3989;
wire n_2837;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_2319;
wire n_1393;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_3655;
wire n_2808;
wire n_3009;
wire n_1276;
wire n_2548;
wire n_1412;
wire n_2679;
wire n_2676;
wire n_1709;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_2930;
wire n_1538;
wire n_1162;
wire n_4206;
wire n_1838;
wire n_1847;
wire n_1199;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_3923;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_2454;
wire n_4371;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_2801;
wire n_1293;
wire n_3120;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_2763;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_2009;
wire n_1888;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_3819;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_2064;
wire n_3978;
wire n_4325;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4372;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_1537;
wire n_3833;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_2671;
wire n_4262;
wire n_4184;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_2629;
wire n_1415;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_4379;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2838;
wire n_2181;
wire n_2479;
wire n_1647;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_4397;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_4391;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_3855;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_2054;
wire n_3765;
wire n_1503;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_3816;
wire n_2623;
wire n_1617;
wire n_1994;
wire n_3113;
wire n_1231;
wire n_1406;
wire n_1279;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_2960;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_3205;
wire n_4156;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_4404;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_3396;
wire n_3701;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_2666;
wire n_2982;
wire n_1692;
wire n_3385;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_2320;
wire n_2339;
wire n_2038;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_4396;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3820;
wire n_4367;
wire n_3741;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_4232;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2457;
wire n_2346;
wire n_4387;
wire n_2312;
wire n_3990;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_2536;
wire n_1592;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_2725;
wire n_1548;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_3787;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_4392;
wire n_3149;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_2897;
wire n_2077;
wire n_1416;
wire n_3614;
wire n_2909;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_1724;
wire n_4285;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_4329;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_3200;
wire n_1664;
wire n_4271;
wire n_1486;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2879;
wire n_2474;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_2033;
wire n_1591;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3077;
wire n_3929;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_3474;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_3984;
wire n_1140;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_3679;
wire n_3779;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_1456;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_4305;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4207;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_3154;
wire n_1551;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_4313;
wire n_4037;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_2240;
wire n_2696;
wire n_1351;
wire n_4063;
wire n_4198;
wire n_1044;
wire n_2436;
wire n_1205;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4339;
wire n_4041;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_2658;
wire n_1684;
wire n_3590;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_2555;
wire n_1381;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_2419;
wire n_1708;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_1082;
wire n_3961;
wire n_2122;
wire n_2512;
wire n_1630;
wire n_3589;
wire n_4102;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_3195;
wire n_3190;
wire n_1519;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3569;
wire n_3548;
wire n_4348;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_1442;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_3953;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_1050;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_4384;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_2701;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2415;
wire n_2309;
wire n_2948;
wire n_3299;
wire n_3041;
wire n_3274;
wire n_2646;
wire n_3715;
wire n_1560;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1363;
wire n_1301;
wire n_3737;
wire n_3913;
wire n_1668;
wire n_1185;
wire n_2903;
wire n_3482;
wire n_3417;
wire n_3866;
wire n_1967;
wire n_1143;
wire n_2233;
wire n_3717;
wire n_3921;
wire n_1579;
wire n_4106;
wire n_1329;
wire n_4034;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_2827;
wire n_3052;
wire n_1688;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_4400;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_3734;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_4402;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_3529;
wire n_3854;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_2468;
wire n_1977;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_4338;
wire n_3492;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_3253;
wire n_2056;
wire n_1636;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_2318;
wire n_2393;
wire n_1575;
wire n_1697;
wire n_3689;
wire n_1735;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2707;
wire n_2793;
wire n_2751;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_2285;
wire n_1446;
wire n_4406;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_2471;
wire n_2298;
wire n_1472;
wire n_1176;
wire n_1807;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_2795;
wire n_4091;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3460;
wire n_3409;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_4316;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_4247;
wire n_2638;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_4409;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_2034;
wire n_1637;
wire n_1687;
wire n_2711;
wire n_1419;
wire n_4336;
wire n_3933;
wire n_2270;
wire n_1653;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_1256;
wire n_2259;
wire n_2794;
wire n_1702;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_2995;
wire n_2494;
wire n_1375;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1929;
wire n_1597;
wire n_2807;
wire n_1164;
wire n_1834;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_1659;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_3450;
wire n_1714;
wire n_1116;
wire n_2000;
wire n_3402;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_3174;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1731;
wire n_2217;
wire n_1453;
wire n_3746;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_1253;
wire n_2201;
wire n_2745;
wire n_2722;
wire n_2117;
wire n_1737;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1777;
wire n_1335;
wire n_1514;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2437;
wire n_2219;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_1726;
wire n_3654;
wire n_1835;
wire n_3035;
wire n_3839;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_3972;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_2532;
wire n_2605;
wire n_1310;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1991;
wire n_2224;
wire n_1399;
wire n_1979;
wire n_1543;
wire n_1533;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_2484;
wire n_4111;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_3928;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_3534;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_3438;
wire n_4098;
wire n_2012;
wire n_3792;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1753;
wire n_1297;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_2806;
wire n_1485;
wire n_4269;
wire n_1184;
wire n_2184;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_2814;
wire n_1570;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_2213;
wire n_2023;
wire n_1170;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_3968;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_2697;
wire n_1461;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_2861;
wire n_1372;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_4380;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2284;
wire n_2187;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_3239;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_2850;
wire n_1747;
wire n_4220;
wire n_4251;
wire n_1817;
wire n_1944;
wire n_1683;
wire n_1530;
wire n_1497;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_3431;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_2996;
wire n_1268;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_4368;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_4393;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_2560;
wire n_2326;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_3584;
wire n_1425;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_3691;
wire n_2889;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_4382;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_4399;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_4401;
wire n_3904;
wire n_2250;
wire n_2678;
wire n_2778;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_2451;
wire n_1520;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_4363;
wire n_1262;
wire n_2691;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_1648;
wire n_4015;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_3627;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_3903;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3859;
wire n_3722;
wire n_3865;
wire n_4171;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_3117;
wire n_1555;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1396;
wire n_2744;
wire n_2030;
wire n_1348;
wire n_2453;
wire n_2397;
wire n_1752;
wire n_2883;
wire n_3115;
wire n_1525;
wire n_4287;
wire n_3509;
wire n_3352;
wire n_4390;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4270;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_3384;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1495;
wire n_1337;
wire n_4231;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1975;
wire n_1321;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_3114;
wire n_3125;
wire n_2594;
wire n_3234;
wire n_2394;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_4407;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_4389;
wire n_3930;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3997;
wire n_2513;
wire n_1275;
wire n_2525;
wire n_1604;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4343;
wire n_4319;
wire n_1493;
wire n_4212;
wire n_4320;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_3694;
wire n_2586;
wire n_1448;
wire n_4245;
wire n_4288;
wire n_4364;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1398;
wire n_1996;
wire n_1879;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_4216;
wire n_4222;
wire n_3939;
wire n_1634;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_1340;
wire n_1558;
wire n_4241;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_2689;
wire n_1990;
wire n_2920;
wire n_3259;
wire n_4265;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_3414;
wire n_2237;
wire n_1622;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_3693;
wire n_1542;
wire n_1251;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

INVx1_ASAP7_75t_L g1024 ( 
.A(n_62),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_884),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_726),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_514),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_813),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_950),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_956),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_165),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_268),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_611),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_419),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_489),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_438),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_473),
.Y(n_1037)
);

CKINVDCx16_ASAP7_75t_R g1038 ( 
.A(n_764),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_716),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_56),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_133),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_878),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_833),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1021),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_346),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_895),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_853),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_537),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_659),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_103),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_228),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_945),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_929),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_346),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_59),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_670),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_823),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_834),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_715),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_711),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_739),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_896),
.Y(n_1062)
);

BUFx10_ASAP7_75t_L g1063 ( 
.A(n_593),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_751),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_770),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_587),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_907),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_492),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_204),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_985),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_848),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_825),
.Y(n_1072)
);

BUFx8_ASAP7_75t_SL g1073 ( 
.A(n_772),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_545),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_257),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_694),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_741),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_868),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_731),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_808),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_844),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_842),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_903),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_496),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_13),
.Y(n_1085)
);

BUFx5_ASAP7_75t_L g1086 ( 
.A(n_696),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_832),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_163),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_914),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_753),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_607),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_607),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_395),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_342),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_934),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_210),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_250),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_548),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_169),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_409),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_992),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_829),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_464),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_423),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_719),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_430),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_251),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_720),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_725),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_239),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_947),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_78),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_988),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_217),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_976),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_951),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_26),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_160),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_297),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_369),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_535),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_35),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_197),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_740),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_595),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_388),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_139),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_854),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_498),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_971),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_804),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_864),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_883),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_578),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_722),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_567),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_560),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_1),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_972),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_647),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1007),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_916),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_979),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_712),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_544),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_623),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_666),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_987),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_850),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_391),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_109),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_341),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_577),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_835),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_736),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_702),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_107),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_974),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_899),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_784),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_695),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_667),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_782),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_481),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_682),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_373),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1015),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_799),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_264),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_15),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1011),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_685),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_409),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_193),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_539),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_503),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_696),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_710),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_452),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_860),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_721),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_890),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_967),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_516),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_955),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_874),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_157),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_977),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_852),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_91),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_13),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_633),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_961),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1002),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_839),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_14),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_640),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_434),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_350),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_52),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_982),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_171),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_547),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_263),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_411),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_905),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_801),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_674),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_713),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_737),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_229),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_818),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_685),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_879),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_525),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_783),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_61),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1004),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_952),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_932),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_918),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_435),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_67),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_503),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_904),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_290),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_996),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_997),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_230),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_908),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_146),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_824),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_857),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_983),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_962),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_661),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_893),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_676),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_270),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_157),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_9),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_958),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_922),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_815),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_316),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_401),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_898),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_939),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_64),
.Y(n_1249)
);

CKINVDCx14_ASAP7_75t_R g1250 ( 
.A(n_769),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_766),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_866),
.Y(n_1252)
);

BUFx5_ASAP7_75t_L g1253 ( 
.A(n_963),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_941),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_733),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_756),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_943),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_851),
.Y(n_1258)
);

CKINVDCx16_ASAP7_75t_R g1259 ( 
.A(n_305),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_240),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_98),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_807),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_674),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_625),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_790),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_109),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_456),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_560),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_697),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_830),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_701),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_183),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_888),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_856),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_708),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_510),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_249),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_287),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_504),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_302),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_998),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_810),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_121),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_923),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_450),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_46),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_50),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_443),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_779),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_841),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_577),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_965),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_466),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1012),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_159),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_949),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_776),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_728),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_569),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_376),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_353),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1001),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_570),
.Y(n_1303)
);

CKINVDCx16_ASAP7_75t_R g1304 ( 
.A(n_894),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_748),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_849),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_553),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_261),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1018),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_97),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_755),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_479),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_730),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_378),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_910),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_798),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_863),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_960),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1006),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_793),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_984),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_887),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_437),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_909),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_153),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_175),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_872),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_110),
.Y(n_1328)
);

CKINVDCx14_ASAP7_75t_R g1329 ( 
.A(n_912),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_248),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_444),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_617),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_131),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1014),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_902),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_215),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_690),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_994),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_991),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_729),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_351),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_921),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_39),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1013),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_590),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1010),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_640),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_480),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_261),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_445),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_423),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_780),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_917),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_199),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_785),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_762),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_714),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_102),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_889),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_180),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_680),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_131),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_937),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_742),
.Y(n_1364)
);

BUFx10_ASAP7_75t_L g1365 ( 
.A(n_19),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_936),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_204),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_765),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_880),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_620),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_749),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_876),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_175),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_535),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_791),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_122),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_453),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_96),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_336),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_820),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_207),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_214),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_734),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_968),
.Y(n_1384)
);

CKINVDCx16_ASAP7_75t_R g1385 ( 
.A(n_700),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_235),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_773),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_375),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_393),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_940),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_892),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_113),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_17),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_698),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_74),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_511),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_752),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_33),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_403),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_846),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_287),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_693),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_678),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_680),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_858),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_964),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_855),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_635),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_100),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_677),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_18),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_135),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_211),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_659),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_817),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_568),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_717),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_120),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_402),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_235),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_202),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_675),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_33),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_590),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_325),
.Y(n_1425)
);

BUFx5_ASAP7_75t_L g1426 ( 
.A(n_582),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_58),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_561),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_316),
.Y(n_1429)
);

BUFx10_ASAP7_75t_L g1430 ( 
.A(n_567),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_156),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_915),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_911),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_620),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_757),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_812),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_390),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_690),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_311),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_794),
.Y(n_1440)
);

CKINVDCx14_ASAP7_75t_R g1441 ( 
.A(n_691),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_995),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_699),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_163),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_34),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_257),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_382),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_981),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_446),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_990),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_74),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_269),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_169),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_930),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1005),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_925),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_744),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_643),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_900),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_875),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_671),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_217),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_870),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_226),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_203),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_119),
.Y(n_1466)
);

INVx4_ASAP7_75t_R g1467 ( 
.A(n_787),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_621),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_437),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_481),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_862),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_684),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_828),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_676),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_709),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_667),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_805),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_547),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_178),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_589),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_331),
.Y(n_1481)
);

CKINVDCx16_ASAP7_75t_R g1482 ( 
.A(n_935),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_938),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_778),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_218),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1017),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_906),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_843),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_601),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_679),
.Y(n_1490)
);

CKINVDCx16_ASAP7_75t_R g1491 ( 
.A(n_8),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_683),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_777),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_262),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_767),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_973),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_989),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1016),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_37),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_873),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_865),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_975),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_761),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_395),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_747),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1023),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_247),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_624),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_361),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_673),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_871),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_745),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_58),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_624),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_732),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_268),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_638),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_600),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_999),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_673),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_455),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_822),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_252),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_79),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_724),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_329),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_459),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_628),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_275),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_788),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_133),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_180),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_424),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_201),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_978),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_78),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_881),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_99),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_532),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_347),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_240),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_605),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_565),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_457),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_517),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_758),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_759),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_304),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_313),
.Y(n_1549)
);

CKINVDCx14_ASAP7_75t_R g1550 ( 
.A(n_702),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_8),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_283),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_546),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_686),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_59),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_993),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_959),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_845),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_321),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_831),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_796),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_276),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_840),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_155),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_957),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_781),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_827),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_255),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_811),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_96),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_290),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_247),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_683),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_418),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_446),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_775),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_919),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_366),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_703),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_986),
.Y(n_1580)
);

CKINVDCx16_ASAP7_75t_R g1581 ( 
.A(n_589),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_681),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_541),
.Y(n_1583)
);

INVxp33_ASAP7_75t_SL g1584 ( 
.A(n_332),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_410),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_370),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1003),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_953),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_299),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_933),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_969),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_196),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_735),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_207),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1000),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_913),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_367),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_819),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_746),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_214),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_565),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_95),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_859),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_25),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_558),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_511),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_789),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_14),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_585),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_738),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_52),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_597),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_587),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_891),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_621),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_897),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_688),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_768),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_141),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_97),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_359),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_954),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_420),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_296),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_102),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_809),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_397),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_400),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_463),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_433),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_882),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_357),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_672),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_802),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_351),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_718),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_419),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_861),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_926),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_190),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_692),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_774),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_475),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_380),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_663),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_410),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_948),
.Y(n_1647)
);

CKINVDCx20_ASAP7_75t_R g1648 ( 
.A(n_1020),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_65),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_216),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_3),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_300),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_224),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_838),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_816),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_573),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_444),
.Y(n_1657)
);

BUFx10_ASAP7_75t_L g1658 ( 
.A(n_806),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_847),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_234),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_727),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_803),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_301),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_173),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_42),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_161),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_318),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_797),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_605),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_885),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_558),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_980),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_927),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_754),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_177),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_284),
.Y(n_1676)
);

BUFx10_ASAP7_75t_L g1677 ( 
.A(n_317),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_208),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1022),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_886),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1019),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_548),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1008),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_416),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_942),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_944),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_750),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_286),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_469),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_2),
.Y(n_1690)
);

BUFx5_ASAP7_75t_L g1691 ( 
.A(n_433),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_415),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_924),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_141),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_453),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_439),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_483),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_631),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_142),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_544),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_510),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_107),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_837),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_836),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_946),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_609),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_786),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_966),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_743),
.Y(n_1709)
);

BUFx10_ASAP7_75t_L g1710 ( 
.A(n_622),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_669),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_826),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_970),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_920),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_568),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_294),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_342),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_396),
.Y(n_1718)
);

INVxp67_ASAP7_75t_SL g1719 ( 
.A(n_901),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_877),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_689),
.Y(n_1721)
);

BUFx10_ASAP7_75t_L g1722 ( 
.A(n_652),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_357),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_760),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_771),
.Y(n_1725)
);

BUFx5_ASAP7_75t_L g1726 ( 
.A(n_795),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_814),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_723),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_251),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_484),
.Y(n_1730)
);

BUFx10_ASAP7_75t_L g1731 ( 
.A(n_867),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_328),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_591),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_205),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1009),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_800),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_427),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_931),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_353),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_792),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_928),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_80),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_603),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_763),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_586),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_SL g1746 ( 
.A(n_668),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_101),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_301),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_176),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_576),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_687),
.Y(n_1751)
);

BUFx10_ASAP7_75t_L g1752 ( 
.A(n_69),
.Y(n_1752)
);

CKINVDCx20_ASAP7_75t_R g1753 ( 
.A(n_391),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_400),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_178),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_332),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_362),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_408),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_56),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_821),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_213),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_869),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_324),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1086),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1319),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1073),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1029),
.Y(n_1767)
);

CKINVDCx14_ASAP7_75t_R g1768 ( 
.A(n_1441),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1086),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1030),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1086),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1042),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1065),
.Y(n_1773)
);

INVxp33_ASAP7_75t_L g1774 ( 
.A(n_1093),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1086),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1047),
.Y(n_1776)
);

INVxp33_ASAP7_75t_SL g1777 ( 
.A(n_1414),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1086),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1426),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1426),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1426),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1426),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1426),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1691),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1691),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1691),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1691),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1691),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1468),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1136),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1468),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1053),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1106),
.Y(n_1793)
);

INVxp33_ASAP7_75t_L g1794 ( 
.A(n_1287),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1063),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1106),
.Y(n_1796)
);

INVxp33_ASAP7_75t_SL g1797 ( 
.A(n_1464),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1727),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1106),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1090),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1140),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1095),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1140),
.Y(n_1803)
);

CKINVDCx16_ASAP7_75t_R g1804 ( 
.A(n_1037),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1140),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1063),
.Y(n_1806)
);

INVxp33_ASAP7_75t_SL g1807 ( 
.A(n_1540),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1165),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1165),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1165),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1059),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1283),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1283),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1283),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1188),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1721),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1721),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1124),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1721),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1097),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1260),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1061),
.Y(n_1822)
);

CKINVDCx16_ASAP7_75t_R g1823 ( 
.A(n_1123),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1057),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1377),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1062),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1253),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1064),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1303),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1378),
.B(n_0),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1360),
.Y(n_1831)
);

CKINVDCx16_ASAP7_75t_R g1832 ( 
.A(n_1259),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1669),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1067),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1761),
.Y(n_1835)
);

INVxp33_ASAP7_75t_SL g1836 ( 
.A(n_1748),
.Y(n_1836)
);

INVxp33_ASAP7_75t_L g1837 ( 
.A(n_1379),
.Y(n_1837)
);

INVxp67_ASAP7_75t_SL g1838 ( 
.A(n_1221),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1024),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1033),
.Y(n_1840)
);

CKINVDCx16_ASAP7_75t_R g1841 ( 
.A(n_1385),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1034),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1755),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_1218),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1281),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1451),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1057),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1071),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1758),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1078),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1079),
.Y(n_1851)
);

INVxp33_ASAP7_75t_SL g1852 ( 
.A(n_1538),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1035),
.Y(n_1853)
);

INVxp33_ASAP7_75t_SL g1854 ( 
.A(n_1573),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1686),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1180),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1051),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1054),
.Y(n_1858)
);

INVxp33_ASAP7_75t_SL g1859 ( 
.A(n_1027),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1081),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1258),
.Y(n_1861)
);

INVxp67_ASAP7_75t_SL g1862 ( 
.A(n_1180),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1074),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1076),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1091),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1096),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1098),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1103),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1083),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1087),
.Y(n_1870)
);

INVxp33_ASAP7_75t_L g1871 ( 
.A(n_1107),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1101),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1491),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1114),
.Y(n_1874)
);

INVxp33_ASAP7_75t_SL g1875 ( 
.A(n_1031),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1258),
.Y(n_1876)
);

INVxp67_ASAP7_75t_SL g1877 ( 
.A(n_1026),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1102),
.Y(n_1878)
);

NAND2xp33_ASAP7_75t_L g1879 ( 
.A(n_1830),
.B(n_1032),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1803),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1768),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1767),
.B(n_1250),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1824),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1770),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1846),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1824),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1852),
.A2(n_1550),
.B1(n_1329),
.B2(n_1581),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1861),
.B(n_1296),
.Y(n_1888)
);

BUFx8_ASAP7_75t_L g1889 ( 
.A(n_1795),
.Y(n_1889)
);

OA21x2_ASAP7_75t_L g1890 ( 
.A1(n_1764),
.A2(n_1043),
.B(n_1039),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1876),
.B(n_1450),
.Y(n_1891)
);

AND2x2_ASAP7_75t_SL g1892 ( 
.A(n_1804),
.B(n_1582),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1800),
.B(n_1547),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1793),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1877),
.B(n_1025),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1796),
.Y(n_1896)
);

OAI21x1_ASAP7_75t_L g1897 ( 
.A1(n_1827),
.A2(n_1089),
.B(n_1080),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1799),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1824),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1847),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1806),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1815),
.B(n_1580),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1838),
.B(n_1028),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1772),
.B(n_1159),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1847),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1845),
.B(n_1131),
.Y(n_1906)
);

AND2x2_ASAP7_75t_SL g1907 ( 
.A(n_1823),
.B(n_1038),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1855),
.B(n_1142),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1847),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1801),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1873),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_L g1912 ( 
.A(n_1776),
.B(n_1036),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1792),
.B(n_1193),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1805),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1808),
.Y(n_1915)
);

INVx6_ASAP7_75t_L g1916 ( 
.A(n_1832),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1765),
.B(n_1304),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1798),
.B(n_1220),
.Y(n_1918)
);

BUFx12f_ASAP7_75t_L g1919 ( 
.A(n_1766),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1809),
.Y(n_1920)
);

AND2x6_ASAP7_75t_L g1921 ( 
.A(n_1820),
.B(n_1174),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1810),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1825),
.B(n_1275),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1811),
.B(n_1339),
.Y(n_1924)
);

INVxp33_ASAP7_75t_SL g1925 ( 
.A(n_1822),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1812),
.Y(n_1926)
);

INVx4_ASAP7_75t_L g1927 ( 
.A(n_1826),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1813),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1828),
.B(n_1455),
.Y(n_1929)
);

OAI22x1_ASAP7_75t_R g1930 ( 
.A1(n_1773),
.A2(n_1121),
.B1(n_1229),
.B2(n_1056),
.Y(n_1930)
);

OAI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1856),
.A2(n_1232),
.B(n_1230),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1814),
.Y(n_1932)
);

BUFx12f_ASAP7_75t_L g1933 ( 
.A(n_1834),
.Y(n_1933)
);

OA21x2_ASAP7_75t_L g1934 ( 
.A1(n_1769),
.A2(n_1046),
.B(n_1044),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1816),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1821),
.Y(n_1936)
);

OAI22x1_ASAP7_75t_SL g1937 ( 
.A1(n_1854),
.A2(n_1241),
.B1(n_1249),
.B2(n_1240),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1848),
.B(n_1471),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1829),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1862),
.B(n_1352),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1771),
.A2(n_1344),
.B(n_1317),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1817),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1819),
.Y(n_1943)
);

INVx6_ASAP7_75t_L g1944 ( 
.A(n_1841),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1775),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1778),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1839),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1850),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1878),
.B(n_1482),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1851),
.B(n_1265),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1840),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1842),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1860),
.B(n_1869),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1870),
.B(n_1265),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1779),
.A2(n_1363),
.B(n_1346),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1780),
.Y(n_1956)
);

AOI22x1_ASAP7_75t_SL g1957 ( 
.A1(n_1802),
.A2(n_1330),
.B1(n_1331),
.B2(n_1312),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1872),
.B(n_1704),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1777),
.A2(n_1584),
.B1(n_1257),
.B2(n_1294),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1781),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1831),
.B(n_1405),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1833),
.Y(n_1962)
);

CKINVDCx16_ASAP7_75t_R g1963 ( 
.A(n_1818),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1837),
.B(n_1658),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1782),
.Y(n_1965)
);

OA21x2_ASAP7_75t_L g1966 ( 
.A1(n_1783),
.A2(n_1058),
.B(n_1052),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1843),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1835),
.B(n_1484),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1790),
.B(n_1435),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1784),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1859),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1774),
.B(n_1658),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1785),
.Y(n_1973)
);

BUFx8_ASAP7_75t_L g1974 ( 
.A(n_1849),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1853),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1789),
.B(n_1791),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1786),
.A2(n_1588),
.B(n_1567),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1857),
.B(n_1577),
.Y(n_1978)
);

INVxp33_ASAP7_75t_SL g1979 ( 
.A(n_1858),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1787),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1788),
.B(n_1599),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1794),
.B(n_1731),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1863),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1875),
.B(n_1655),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1871),
.B(n_1272),
.Y(n_1985)
);

INVx6_ASAP7_75t_L g1986 ( 
.A(n_1797),
.Y(n_1986)
);

AND2x6_ASAP7_75t_L g1987 ( 
.A(n_1864),
.B(n_1286),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1865),
.B(n_1731),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1866),
.B(n_1060),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1867),
.B(n_1670),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1868),
.B(n_1072),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1807),
.A2(n_1383),
.B1(n_1417),
.B2(n_1227),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1874),
.B(n_1719),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1844),
.B(n_1077),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1836),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1852),
.A2(n_1332),
.B1(n_1394),
.B2(n_1389),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1768),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1803),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1803),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1852),
.A2(n_1475),
.B1(n_1495),
.B2(n_1457),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1803),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1803),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1803),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1827),
.A2(n_1105),
.B(n_1082),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1861),
.B(n_1108),
.Y(n_2005)
);

BUFx6f_ASAP7_75t_L g2006 ( 
.A(n_1803),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1803),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1852),
.A2(n_1401),
.B1(n_1516),
.B2(n_1404),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1767),
.B(n_1113),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1803),
.Y(n_2010)
);

INVx4_ASAP7_75t_L g2011 ( 
.A(n_1767),
.Y(n_2011)
);

AND2x6_ASAP7_75t_L g2012 ( 
.A(n_1861),
.B(n_1299),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1803),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1803),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1803),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1859),
.B(n_1115),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1803),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1803),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1861),
.Y(n_2019)
);

BUFx8_ASAP7_75t_SL g2020 ( 
.A(n_1766),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1768),
.B(n_1138),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1803),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1852),
.A2(n_1566),
.B1(n_1610),
.B2(n_1506),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1767),
.B(n_1116),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1803),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1803),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1861),
.B(n_1139),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1803),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1803),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1803),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1768),
.B(n_1333),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1803),
.Y(n_2032)
);

OA21x2_ASAP7_75t_L g2033 ( 
.A1(n_1764),
.A2(n_1143),
.B(n_1141),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1803),
.Y(n_2034)
);

OA21x2_ASAP7_75t_L g2035 ( 
.A1(n_1764),
.A2(n_1149),
.B(n_1148),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1803),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1803),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1861),
.B(n_1155),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1803),
.Y(n_2039)
);

BUFx8_ASAP7_75t_L g2040 ( 
.A(n_1795),
.Y(n_2040)
);

AOI22x1_ASAP7_75t_SL g2041 ( 
.A1(n_1773),
.A2(n_1627),
.B1(n_1633),
.B2(n_1601),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1767),
.B(n_1171),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1852),
.A2(n_1638),
.B1(n_1642),
.B2(n_1614),
.Y(n_2043)
);

INVx4_ASAP7_75t_L g2044 ( 
.A(n_1767),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1803),
.Y(n_2045)
);

OA21x2_ASAP7_75t_L g2046 ( 
.A1(n_1764),
.A2(n_1182),
.B(n_1181),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1861),
.B(n_1185),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1803),
.Y(n_2048)
);

INVx4_ASAP7_75t_L g2049 ( 
.A(n_1767),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1803),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1803),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1803),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1803),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1767),
.B(n_1189),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1768),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1803),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1767),
.B(n_1194),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1820),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1767),
.B(n_1207),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1803),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1803),
.Y(n_2061)
);

BUFx12f_ASAP7_75t_L g2062 ( 
.A(n_1766),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1852),
.A2(n_1418),
.B1(n_1041),
.B2(n_1045),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1767),
.B(n_1212),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1767),
.B(n_1225),
.Y(n_2065)
);

CKINVDCx6p67_ASAP7_75t_R g2066 ( 
.A(n_1804),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1803),
.Y(n_2067)
);

CKINVDCx8_ASAP7_75t_R g2068 ( 
.A(n_1804),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1768),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1803),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1803),
.Y(n_2071)
);

OA21x2_ASAP7_75t_L g2072 ( 
.A1(n_1764),
.A2(n_1243),
.B(n_1237),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1803),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1803),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1803),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1803),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1852),
.A2(n_1654),
.B1(n_1720),
.B2(n_1648),
.Y(n_2077)
);

INVx5_ASAP7_75t_L g2078 ( 
.A(n_1824),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1767),
.B(n_1255),
.Y(n_2079)
);

XNOR2xp5_ASAP7_75t_L g2080 ( 
.A(n_1773),
.B(n_1675),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1790),
.B(n_1408),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1803),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1852),
.A2(n_1048),
.B1(n_1049),
.B2(n_1040),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_1766),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1768),
.B(n_1373),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1803),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1768),
.B(n_1445),
.Y(n_2087)
);

BUFx12f_ASAP7_75t_L g2088 ( 
.A(n_1766),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1803),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1803),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1824),
.Y(n_2091)
);

OA21x2_ASAP7_75t_L g2092 ( 
.A1(n_1764),
.A2(n_1273),
.B(n_1256),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1803),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_L g2094 ( 
.A(n_1861),
.B(n_1306),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1861),
.B(n_1311),
.Y(n_2095)
);

OA21x2_ASAP7_75t_L g2096 ( 
.A1(n_1764),
.A2(n_1321),
.B(n_1318),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1803),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1767),
.B(n_1322),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1803),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1803),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1803),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1767),
.B(n_1324),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1803),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1803),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1767),
.B(n_1327),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1824),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1803),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1767),
.B(n_1335),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_1820),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1852),
.A2(n_1055),
.B1(n_1066),
.B2(n_1050),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1803),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1803),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1804),
.B(n_1094),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1767),
.B(n_1355),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1861),
.B(n_1356),
.Y(n_2115)
);

BUFx3_ASAP7_75t_L g2116 ( 
.A(n_1820),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1803),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1803),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1767),
.B(n_1359),
.Y(n_2119)
);

BUFx8_ASAP7_75t_L g2120 ( 
.A(n_1795),
.Y(n_2120)
);

OA21x2_ASAP7_75t_L g2121 ( 
.A1(n_1764),
.A2(n_1387),
.B(n_1366),
.Y(n_2121)
);

XNOR2x1_ASAP7_75t_L g2122 ( 
.A(n_1790),
.B(n_1068),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1824),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1803),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_1861),
.B(n_1391),
.Y(n_2125)
);

INVx4_ASAP7_75t_L g2126 ( 
.A(n_1767),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_1846),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1803),
.Y(n_2128)
);

BUFx12f_ASAP7_75t_L g2129 ( 
.A(n_1766),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1803),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1803),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1767),
.B(n_1397),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1803),
.Y(n_2133)
);

BUFx6f_ASAP7_75t_L g2134 ( 
.A(n_1803),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1852),
.A2(n_1069),
.B1(n_1084),
.B2(n_1075),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1803),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1803),
.Y(n_2137)
);

OA21x2_ASAP7_75t_L g2138 ( 
.A1(n_1764),
.A2(n_1432),
.B(n_1406),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_1861),
.B(n_1436),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1803),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1767),
.B(n_1440),
.Y(n_2141)
);

CKINVDCx20_ASAP7_75t_R g2142 ( 
.A(n_1773),
.Y(n_2142)
);

OA21x2_ASAP7_75t_L g2143 ( 
.A1(n_1764),
.A2(n_1463),
.B(n_1442),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1803),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1803),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1803),
.Y(n_2146)
);

OAI21x1_ASAP7_75t_L g2147 ( 
.A1(n_1827),
.A2(n_1483),
.B(n_1477),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_L g2148 ( 
.A(n_1803),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1803),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1803),
.Y(n_2150)
);

INVxp33_ASAP7_75t_L g2151 ( 
.A(n_2081),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_2091),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1947),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1886),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1936),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1951),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1884),
.Y(n_2157)
);

BUFx3_ASAP7_75t_L g2158 ( 
.A(n_1939),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_R g2159 ( 
.A(n_1948),
.B(n_1109),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1952),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_2020),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1900),
.Y(n_2162)
);

CKINVDCx20_ASAP7_75t_R g2163 ( 
.A(n_2142),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1967),
.Y(n_2164)
);

NAND2xp33_ASAP7_75t_R g2165 ( 
.A(n_1994),
.B(n_1085),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1969),
.B(n_1111),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1925),
.Y(n_2167)
);

CKINVDCx20_ASAP7_75t_R g2168 ( 
.A(n_1963),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1946),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1933),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1909),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1919),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1956),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_2062),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1960),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1965),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_2084),
.Y(n_2177)
);

CKINVDCx20_ASAP7_75t_R g2178 ( 
.A(n_2066),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2091),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_SL g2180 ( 
.A1(n_1996),
.A2(n_1753),
.B1(n_1428),
.B2(n_1545),
.Y(n_2180)
);

BUFx10_ASAP7_75t_L g2181 ( 
.A(n_1986),
.Y(n_2181)
);

CKINVDCx20_ASAP7_75t_R g2182 ( 
.A(n_2068),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_2088),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_R g2184 ( 
.A(n_2129),
.B(n_1128),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1927),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_2011),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_2044),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_2049),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_2106),
.Y(n_2189)
);

BUFx10_ASAP7_75t_L g2190 ( 
.A(n_1916),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1998),
.Y(n_2191)
);

INVx3_ASAP7_75t_L g2192 ( 
.A(n_2106),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_2126),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1881),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_1944),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1980),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1985),
.Y(n_2197)
);

CKINVDCx20_ASAP7_75t_R g2198 ( 
.A(n_2080),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1997),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2001),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1945),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1970),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2002),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1973),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_2055),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2006),
.Y(n_2206)
);

INVx2_ASAP7_75t_SL g2207 ( 
.A(n_2021),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_2069),
.Y(n_2208)
);

CKINVDCx5p33_ASAP7_75t_R g2209 ( 
.A(n_1953),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1889),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_2040),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_2120),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1971),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2018),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_2122),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_2058),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1895),
.B(n_1130),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1906),
.B(n_1132),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_2000),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_2023),
.Y(n_2220)
);

AND3x2_ASAP7_75t_L g2221 ( 
.A(n_2016),
.B(n_1190),
.C(n_1184),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2109),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2061),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1972),
.B(n_1094),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_2043),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_2077),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2116),
.Y(n_2227)
);

NOR2xp67_ASAP7_75t_L g2228 ( 
.A(n_1882),
.B(n_1133),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1983),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1899),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1976),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_1885),
.Y(n_2232)
);

OAI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_1959),
.A2(n_1559),
.B1(n_1409),
.B2(n_1092),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_R g2234 ( 
.A(n_1912),
.B(n_2019),
.Y(n_2234)
);

CKINVDCx20_ASAP7_75t_R g2235 ( 
.A(n_1992),
.Y(n_2235)
);

CKINVDCx20_ASAP7_75t_R g2236 ( 
.A(n_1911),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1975),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2123),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2067),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2076),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_1907),
.Y(n_2241)
);

BUFx10_ASAP7_75t_L g2242 ( 
.A(n_1923),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1894),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1896),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_R g2245 ( 
.A(n_1879),
.B(n_1949),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_2127),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1898),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1979),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_2123),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1950),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1954),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1915),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1904),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1913),
.Y(n_2254)
);

CKINVDCx20_ASAP7_75t_R g2255 ( 
.A(n_1995),
.Y(n_2255)
);

CKINVDCx20_ASAP7_75t_R g2256 ( 
.A(n_1930),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2089),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1924),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1982),
.B(n_1349),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_1883),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2009),
.B(n_1532),
.Y(n_2261)
);

CKINVDCx20_ASAP7_75t_R g2262 ( 
.A(n_2008),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1905),
.Y(n_2263)
);

BUFx2_ASAP7_75t_L g2264 ( 
.A(n_2012),
.Y(n_2264)
);

CKINVDCx20_ASAP7_75t_R g2265 ( 
.A(n_1903),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1929),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1942),
.Y(n_2267)
);

CKINVDCx20_ASAP7_75t_R g2268 ( 
.A(n_1957),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_1964),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2090),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1943),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1880),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1938),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_1958),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2103),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2031),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2003),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_2111),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_1892),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_2117),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_2041),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2133),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_2024),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1940),
.B(n_1135),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2010),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_1917),
.B(n_1349),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_2134),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2013),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2017),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2022),
.Y(n_2290)
);

CKINVDCx20_ASAP7_75t_R g2291 ( 
.A(n_2113),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_2042),
.Y(n_2292)
);

NAND2xp33_ASAP7_75t_R g2293 ( 
.A(n_1908),
.B(n_1088),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2030),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_2054),
.Y(n_2295)
);

CKINVDCx20_ASAP7_75t_R g2296 ( 
.A(n_2083),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_2057),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2148),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_2059),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2032),
.Y(n_2300)
);

NAND2xp33_ASAP7_75t_R g2301 ( 
.A(n_1918),
.B(n_1099),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2034),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_2064),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_2065),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_2079),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2098),
.Y(n_2306)
);

AOI21x1_ASAP7_75t_L g2307 ( 
.A1(n_1981),
.A2(n_1501),
.B(n_1486),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2036),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_R g2309 ( 
.A(n_1901),
.B(n_1154),
.Y(n_2309)
);

CKINVDCx20_ASAP7_75t_R g2310 ( 
.A(n_2135),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2102),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2105),
.B(n_1158),
.Y(n_2312)
);

HB1xp67_ASAP7_75t_L g2313 ( 
.A(n_2085),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_2108),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2050),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_2114),
.Y(n_2316)
);

AOI22x1_ASAP7_75t_SL g2317 ( 
.A1(n_1937),
.A2(n_1104),
.B1(n_1110),
.B2(n_1100),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_2119),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_R g2319 ( 
.A(n_1984),
.B(n_1160),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_2132),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_2141),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_2110),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2051),
.Y(n_2323)
);

AOI22x1_ASAP7_75t_L g2324 ( 
.A1(n_1893),
.A2(n_1530),
.B1(n_1537),
.B2(n_1512),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_1887),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_1888),
.Y(n_2326)
);

AOI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_1902),
.A2(n_1167),
.B1(n_1168),
.B2(n_1163),
.Y(n_2327)
);

INVxp67_ASAP7_75t_L g2328 ( 
.A(n_1988),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_R g2329 ( 
.A(n_2087),
.B(n_1178),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_1891),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_2063),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2056),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2073),
.Y(n_2333)
);

INVxp67_ASAP7_75t_L g2334 ( 
.A(n_1987),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2012),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2075),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_SL g2337 ( 
.A(n_1987),
.B(n_1746),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2082),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1993),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_1921),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2086),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_1921),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2093),
.Y(n_2343)
);

CKINVDCx20_ASAP7_75t_R g2344 ( 
.A(n_1974),
.Y(n_2344)
);

CKINVDCx20_ASAP7_75t_R g2345 ( 
.A(n_1990),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_2005),
.Y(n_2346)
);

CKINVDCx20_ASAP7_75t_R g2347 ( 
.A(n_1961),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_2027),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_2038),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2100),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_2047),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_R g2352 ( 
.A(n_1962),
.B(n_1183),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_2095),
.Y(n_2353)
);

CKINVDCx20_ASAP7_75t_R g2354 ( 
.A(n_1968),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2101),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_1910),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2115),
.Y(n_2357)
);

CKINVDCx20_ASAP7_75t_R g2358 ( 
.A(n_1989),
.Y(n_2358)
);

CKINVDCx20_ASAP7_75t_R g2359 ( 
.A(n_1991),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2107),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_2125),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2139),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1978),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_1935),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_2112),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_2124),
.Y(n_2366)
);

CKINVDCx16_ASAP7_75t_R g2367 ( 
.A(n_2094),
.Y(n_2367)
);

NOR2xp67_ASAP7_75t_L g2368 ( 
.A(n_2014),
.B(n_1186),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2131),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2137),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2144),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2145),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_1914),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_1920),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_1922),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2004),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_1926),
.Y(n_2377)
);

BUFx2_ASAP7_75t_L g2378 ( 
.A(n_2029),
.Y(n_2378)
);

NOR2xp67_ASAP7_75t_L g2379 ( 
.A(n_2060),
.B(n_1195),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1928),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2147),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_1897),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_1932),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_2104),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1999),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_2007),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2015),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2025),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_2026),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2028),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2037),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_L g2392 ( 
.A(n_2283),
.B(n_1201),
.Y(n_2392)
);

INVx3_ASAP7_75t_L g2393 ( 
.A(n_2263),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2292),
.B(n_1206),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2295),
.B(n_1112),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2297),
.B(n_2299),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2263),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2303),
.B(n_1209),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2300),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2304),
.B(n_1890),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2243),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2308),
.Y(n_2402)
);

INVx3_ASAP7_75t_L g2403 ( 
.A(n_2263),
.Y(n_2403)
);

AND2x4_ASAP7_75t_L g2404 ( 
.A(n_2280),
.B(n_2039),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2315),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2305),
.B(n_1117),
.Y(n_2406)
);

BUFx6f_ASAP7_75t_L g2407 ( 
.A(n_2152),
.Y(n_2407)
);

INVx5_ASAP7_75t_L g2408 ( 
.A(n_2190),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2244),
.Y(n_2409)
);

BUFx4f_ASAP7_75t_L g2410 ( 
.A(n_2195),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2155),
.B(n_2045),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2197),
.B(n_2048),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2323),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2306),
.B(n_1934),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2247),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2158),
.B(n_2216),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2333),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2252),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2151),
.B(n_2052),
.Y(n_2419)
);

AND2x6_ASAP7_75t_L g2420 ( 
.A(n_2286),
.B(n_1119),
.Y(n_2420)
);

HB1xp67_ASAP7_75t_L g2421 ( 
.A(n_2363),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2338),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2311),
.B(n_1210),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2345),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2242),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2372),
.Y(n_2426)
);

BUFx2_ASAP7_75t_L g2427 ( 
.A(n_2236),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2267),
.Y(n_2428)
);

BUFx10_ASAP7_75t_L g2429 ( 
.A(n_2161),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_2287),
.B(n_2053),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2152),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2271),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_2152),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2314),
.B(n_1966),
.Y(n_2434)
);

INVx4_ASAP7_75t_L g2435 ( 
.A(n_2278),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_2278),
.Y(n_2436)
);

BUFx10_ASAP7_75t_L g2437 ( 
.A(n_2167),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2316),
.B(n_2318),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2272),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2277),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2369),
.Y(n_2441)
);

INVxp67_ASAP7_75t_L g2442 ( 
.A(n_2301),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2278),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2320),
.A2(n_1216),
.B1(n_1219),
.B2(n_1214),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2369),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2380),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2390),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2321),
.B(n_2033),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2285),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2253),
.B(n_1118),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2288),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2287),
.B(n_2070),
.Y(n_2452)
);

BUFx8_ASAP7_75t_SL g2453 ( 
.A(n_2182),
.Y(n_2453)
);

INVxp67_ASAP7_75t_SL g2454 ( 
.A(n_2189),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_2254),
.B(n_1228),
.Y(n_2455)
);

AND2x6_ASAP7_75t_L g2456 ( 
.A(n_2224),
.B(n_1120),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2258),
.B(n_2035),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2289),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2215),
.B(n_1553),
.Y(n_2459)
);

AND2x4_ASAP7_75t_L g2460 ( 
.A(n_2356),
.B(n_2071),
.Y(n_2460)
);

NOR2x1p5_ASAP7_75t_L g2461 ( 
.A(n_2210),
.B(n_1122),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2364),
.B(n_2074),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2290),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2266),
.B(n_1233),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2294),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2302),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2273),
.B(n_2274),
.Y(n_2467)
);

AND2x6_ASAP7_75t_L g2468 ( 
.A(n_2259),
.B(n_1125),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2209),
.B(n_1127),
.Y(n_2469)
);

NAND3x1_ASAP7_75t_L g2470 ( 
.A(n_2327),
.B(n_2261),
.C(n_2217),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2378),
.B(n_2097),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2260),
.Y(n_2472)
);

BUFx2_ASAP7_75t_L g2473 ( 
.A(n_2265),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2179),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2269),
.B(n_1129),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2312),
.B(n_2046),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2332),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2336),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2328),
.B(n_1145),
.Y(n_2479)
);

INVx4_ASAP7_75t_SL g2480 ( 
.A(n_2180),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2169),
.A2(n_2072),
.B1(n_2096),
.B2(n_2092),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2190),
.Y(n_2482)
);

OR2x2_ASAP7_75t_L g2483 ( 
.A(n_2232),
.B(n_1621),
.Y(n_2483)
);

BUFx2_ASAP7_75t_L g2484 ( 
.A(n_2347),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_2242),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2201),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2179),
.Y(n_2487)
);

INVx3_ASAP7_75t_L g2488 ( 
.A(n_2260),
.Y(n_2488)
);

INVx4_ASAP7_75t_L g2489 ( 
.A(n_2384),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2157),
.Y(n_2490)
);

OR2x6_ASAP7_75t_L g2491 ( 
.A(n_2264),
.B(n_1246),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2202),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2341),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_2248),
.B(n_1151),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2343),
.Y(n_2495)
);

BUFx2_ASAP7_75t_L g2496 ( 
.A(n_2354),
.Y(n_2496)
);

INVx3_ASAP7_75t_L g2497 ( 
.A(n_2179),
.Y(n_2497)
);

BUFx10_ASAP7_75t_L g2498 ( 
.A(n_2170),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2191),
.B(n_2099),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2181),
.Y(n_2500)
);

BUFx8_ASAP7_75t_SL g2501 ( 
.A(n_2178),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2173),
.B(n_2121),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_2255),
.Y(n_2503)
);

INVx1_ASAP7_75t_SL g2504 ( 
.A(n_2358),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2350),
.Y(n_2505)
);

INVx3_ASAP7_75t_L g2506 ( 
.A(n_2189),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2200),
.B(n_2118),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2355),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2360),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2204),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2370),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2192),
.Y(n_2512)
);

BUFx10_ASAP7_75t_L g2513 ( 
.A(n_2172),
.Y(n_2513)
);

OR2x6_ASAP7_75t_L g2514 ( 
.A(n_2207),
.B(n_1278),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_L g2515 ( 
.A1(n_2175),
.A2(n_2196),
.B1(n_2176),
.B2(n_2138),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2371),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2229),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2276),
.B(n_2128),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2181),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2385),
.Y(n_2520)
);

AND2x6_ASAP7_75t_L g2521 ( 
.A(n_2231),
.B(n_1126),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2163),
.Y(n_2522)
);

AND2x6_ASAP7_75t_L g2523 ( 
.A(n_2222),
.B(n_1134),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2391),
.Y(n_2524)
);

AO22x2_ASAP7_75t_L g2525 ( 
.A1(n_2317),
.A2(n_1146),
.B1(n_1147),
.B2(n_1137),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2154),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2153),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_2156),
.Y(n_2528)
);

INVx4_ASAP7_75t_L g2529 ( 
.A(n_2373),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2228),
.B(n_2143),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2162),
.Y(n_2531)
);

AND2x6_ASAP7_75t_L g2532 ( 
.A(n_2227),
.B(n_1150),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2171),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2245),
.B(n_1234),
.Y(n_2534)
);

INVxp67_ASAP7_75t_L g2535 ( 
.A(n_2293),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2230),
.Y(n_2536)
);

BUFx10_ASAP7_75t_L g2537 ( 
.A(n_2174),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2237),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_SL g2539 ( 
.A(n_2177),
.B(n_1746),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2313),
.B(n_1152),
.Y(n_2540)
);

AND2x6_ASAP7_75t_L g2541 ( 
.A(n_2203),
.B(n_1162),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2284),
.B(n_1931),
.Y(n_2542)
);

AOI22xp5_ASAP7_75t_L g2543 ( 
.A1(n_2359),
.A2(n_1242),
.B1(n_1244),
.B2(n_1235),
.Y(n_2543)
);

AOI21x1_ASAP7_75t_L g2544 ( 
.A1(n_2376),
.A2(n_1955),
.B(n_1941),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2365),
.Y(n_2545)
);

OAI22xp33_ASAP7_75t_SL g2546 ( 
.A1(n_2219),
.A2(n_1557),
.B1(n_1565),
.B2(n_1556),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_L g2547 ( 
.A(n_2334),
.B(n_1153),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2192),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2366),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2238),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2250),
.B(n_2130),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2374),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2234),
.B(n_1247),
.Y(n_2553)
);

AND2x4_ASAP7_75t_L g2554 ( 
.A(n_2206),
.B(n_2136),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2319),
.B(n_1587),
.Y(n_2555)
);

OR2x2_ASAP7_75t_L g2556 ( 
.A(n_2246),
.B(n_2140),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2238),
.Y(n_2557)
);

BUFx4f_ASAP7_75t_L g2558 ( 
.A(n_2500),
.Y(n_2558)
);

INVxp67_ASAP7_75t_L g2559 ( 
.A(n_2540),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2401),
.Y(n_2560)
);

AO22x2_ASAP7_75t_L g2561 ( 
.A1(n_2480),
.A2(n_2233),
.B1(n_1173),
.B2(n_1177),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2438),
.B(n_2251),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2399),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2396),
.B(n_2220),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_2408),
.B(n_2214),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2409),
.Y(n_2566)
);

INVx4_ASAP7_75t_L g2567 ( 
.A(n_2482),
.Y(n_2567)
);

INVxp67_ASAP7_75t_L g2568 ( 
.A(n_2419),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2402),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2415),
.Y(n_2570)
);

A2O1A1Ixp33_ASAP7_75t_L g2571 ( 
.A1(n_2400),
.A2(n_2381),
.B(n_2226),
.C(n_2225),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2418),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2414),
.A2(n_2322),
.B1(n_2324),
.B2(n_2331),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2467),
.B(n_2367),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2428),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2432),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2395),
.B(n_2213),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2520),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2442),
.B(n_2535),
.Y(n_2579)
);

INVxp67_ASAP7_75t_L g2580 ( 
.A(n_2412),
.Y(n_2580)
);

INVxp67_ASAP7_75t_L g2581 ( 
.A(n_2556),
.Y(n_2581)
);

AOI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2470),
.A2(n_2325),
.B1(n_2310),
.B2(n_2296),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2524),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_2471),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2434),
.B(n_2185),
.Y(n_2585)
);

INVx2_ASAP7_75t_SL g2586 ( 
.A(n_2551),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2406),
.B(n_2186),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2439),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2448),
.A2(n_2235),
.B1(n_2262),
.B2(n_2382),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2405),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2413),
.Y(n_2591)
);

OAI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2457),
.A2(n_2339),
.B1(n_2187),
.B2(n_2193),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2440),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2504),
.B(n_2279),
.Y(n_2594)
);

NAND2x1p5_ASAP7_75t_L g2595 ( 
.A(n_2416),
.B(n_2435),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2449),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2451),
.Y(n_2597)
);

NAND2x1p5_ASAP7_75t_L g2598 ( 
.A(n_2489),
.B(n_2249),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2458),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2502),
.A2(n_2382),
.B1(n_2218),
.B2(n_1590),
.Y(n_2600)
);

A2O1A1Ixp33_ASAP7_75t_L g2601 ( 
.A1(n_2469),
.A2(n_2166),
.B(n_2241),
.C(n_2188),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2479),
.Y(n_2602)
);

INVxp67_ASAP7_75t_L g2603 ( 
.A(n_2475),
.Y(n_2603)
);

INVxp67_ASAP7_75t_L g2604 ( 
.A(n_2484),
.Y(n_2604)
);

NAND2x1p5_ASAP7_75t_L g2605 ( 
.A(n_2529),
.B(n_2249),
.Y(n_2605)
);

AO22x2_ASAP7_75t_L g2606 ( 
.A1(n_2459),
.A2(n_1187),
.B1(n_1191),
.B2(n_1164),
.Y(n_2606)
);

OAI22xp33_ASAP7_75t_L g2607 ( 
.A1(n_2545),
.A2(n_2337),
.B1(n_2335),
.B2(n_2165),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2463),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2465),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2417),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2422),
.Y(n_2611)
);

BUFx3_ASAP7_75t_L g2612 ( 
.A(n_2397),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2426),
.Y(n_2613)
);

BUFx2_ASAP7_75t_L g2614 ( 
.A(n_2424),
.Y(n_2614)
);

NAND2x1p5_ASAP7_75t_L g2615 ( 
.A(n_2552),
.B(n_2160),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2450),
.B(n_2375),
.Y(n_2616)
);

NOR2x1p5_ASAP7_75t_L g2617 ( 
.A(n_2490),
.B(n_2211),
.Y(n_2617)
);

NAND2x1p5_ASAP7_75t_L g2618 ( 
.A(n_2497),
.B(n_2164),
.Y(n_2618)
);

AO22x2_ASAP7_75t_L g2619 ( 
.A1(n_2549),
.A2(n_1197),
.B1(n_1198),
.B2(n_1196),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2446),
.Y(n_2620)
);

OR2x2_ASAP7_75t_SL g2621 ( 
.A(n_2421),
.B(n_2256),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2494),
.B(n_2340),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2491),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2519),
.B(n_2223),
.Y(n_2624)
);

OAI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2546),
.A2(n_2342),
.B1(n_2387),
.B2(n_2388),
.C(n_2386),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2407),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_L g2627 ( 
.A1(n_2515),
.A2(n_2382),
.B1(n_1593),
.B2(n_1607),
.Y(n_2627)
);

BUFx3_ASAP7_75t_L g2628 ( 
.A(n_2522),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2531),
.Y(n_2629)
);

INVx3_ASAP7_75t_L g2630 ( 
.A(n_2431),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2486),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2555),
.B(n_2444),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2427),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2466),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2477),
.Y(n_2635)
);

AO22x2_ASAP7_75t_L g2636 ( 
.A1(n_2483),
.A2(n_1203),
.B1(n_1217),
.B2(n_1200),
.Y(n_2636)
);

CKINVDCx20_ASAP7_75t_R g2637 ( 
.A(n_2453),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2478),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2420),
.A2(n_2291),
.B1(n_2383),
.B2(n_2377),
.Y(n_2639)
);

AOI22x1_ASAP7_75t_L g2640 ( 
.A1(n_2538),
.A2(n_2389),
.B1(n_2348),
.B2(n_2349),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2518),
.B(n_2346),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2394),
.B(n_2194),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2492),
.Y(n_2643)
);

BUFx6f_ASAP7_75t_L g2644 ( 
.A(n_2433),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_2501),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2493),
.B(n_2159),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2441),
.B(n_2329),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2495),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2547),
.B(n_2351),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2505),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2510),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2411),
.B(n_2239),
.Y(n_2652)
);

INVxp67_ASAP7_75t_L g2653 ( 
.A(n_2496),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_2398),
.B(n_2199),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2445),
.B(n_2353),
.Y(n_2655)
);

OR2x2_ASAP7_75t_L g2656 ( 
.A(n_2473),
.B(n_2205),
.Y(n_2656)
);

AOI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2627),
.A2(n_2476),
.B(n_2542),
.Y(n_2657)
);

OAI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2616),
.A2(n_2543),
.B1(n_2514),
.B2(n_2425),
.Y(n_2658)
);

AOI21xp5_ASAP7_75t_L g2659 ( 
.A1(n_2632),
.A2(n_2530),
.B(n_2534),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2560),
.Y(n_2660)
);

OAI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2571),
.A2(n_2481),
.B(n_2508),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2602),
.B(n_2603),
.Y(n_2662)
);

OAI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2585),
.A2(n_2511),
.B(n_2509),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2559),
.B(n_2456),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2566),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2587),
.B(n_2456),
.Y(n_2666)
);

INVx4_ASAP7_75t_L g2667 ( 
.A(n_2558),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2564),
.A2(n_2392),
.B1(n_2420),
.B2(n_2468),
.Y(n_2668)
);

OAI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2600),
.A2(n_2516),
.B(n_2423),
.Y(n_2669)
);

AOI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2647),
.A2(n_2553),
.B(n_2454),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2586),
.B(n_2437),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2644),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2589),
.B(n_2410),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2570),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2577),
.B(n_2641),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2568),
.B(n_2468),
.Y(n_2676)
);

OAI21xp33_ASAP7_75t_L g2677 ( 
.A1(n_2580),
.A2(n_2539),
.B(n_2464),
.Y(n_2677)
);

INVx5_ASAP7_75t_L g2678 ( 
.A(n_2644),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2572),
.B(n_2455),
.Y(n_2679)
);

O2A1O1Ixp33_ASAP7_75t_L g2680 ( 
.A1(n_2607),
.A2(n_2517),
.B(n_2447),
.C(n_2526),
.Y(n_2680)
);

AOI21xp5_ASAP7_75t_L g2681 ( 
.A1(n_2646),
.A2(n_2533),
.B(n_2536),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2574),
.B(n_2485),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2563),
.Y(n_2683)
);

INVx3_ASAP7_75t_L g2684 ( 
.A(n_2612),
.Y(n_2684)
);

A2O1A1Ixp33_ASAP7_75t_L g2685 ( 
.A1(n_2573),
.A2(n_2557),
.B(n_2550),
.C(n_2512),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2645),
.Y(n_2686)
);

NOR2x1p5_ASAP7_75t_SL g2687 ( 
.A(n_2569),
.B(n_2544),
.Y(n_2687)
);

AOI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2579),
.A2(n_2521),
.B1(n_2198),
.B2(n_2523),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2655),
.A2(n_2548),
.B(n_2506),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2575),
.B(n_2576),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2581),
.B(n_2622),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2578),
.B(n_2521),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2583),
.B(n_2523),
.Y(n_2693)
);

AOI21xp5_ASAP7_75t_L g2694 ( 
.A1(n_2590),
.A2(n_2361),
.B(n_2357),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2649),
.B(n_2503),
.Y(n_2695)
);

AND2x2_ASAP7_75t_SL g2696 ( 
.A(n_2582),
.B(n_2474),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2594),
.B(n_2208),
.Y(n_2697)
);

NAND2x1_ASAP7_75t_L g2698 ( 
.A(n_2591),
.B(n_2487),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2588),
.B(n_2532),
.Y(n_2699)
);

AOI21xp5_ASAP7_75t_L g2700 ( 
.A1(n_2610),
.A2(n_2362),
.B(n_2330),
.Y(n_2700)
);

AOI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2611),
.A2(n_2326),
.B(n_2436),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2642),
.A2(n_2654),
.B1(n_2592),
.B2(n_2562),
.Y(n_2702)
);

AOI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2625),
.A2(n_2532),
.B1(n_2168),
.B2(n_2379),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2604),
.B(n_2443),
.Y(n_2704)
);

INVx4_ASAP7_75t_L g2705 ( 
.A(n_2628),
.Y(n_2705)
);

A2O1A1Ixp33_ASAP7_75t_L g2706 ( 
.A1(n_2593),
.A2(n_2596),
.B(n_2599),
.C(n_2597),
.Y(n_2706)
);

AOI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2613),
.A2(n_2462),
.B(n_2460),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2608),
.B(n_2352),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2614),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2620),
.A2(n_2404),
.B(n_2527),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2609),
.B(n_2472),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2629),
.Y(n_2712)
);

AOI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_2631),
.A2(n_2528),
.B(n_2488),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2634),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2635),
.B(n_2368),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2643),
.A2(n_2403),
.B(n_2393),
.Y(n_2716)
);

AOI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2651),
.A2(n_2507),
.B(n_2499),
.Y(n_2717)
);

AOI21xp33_ASAP7_75t_L g2718 ( 
.A1(n_2656),
.A2(n_2554),
.B(n_2452),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2639),
.B(n_2498),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2638),
.B(n_2430),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2648),
.A2(n_1467),
.B(n_1977),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2650),
.A2(n_1070),
.B(n_1057),
.Y(n_2722)
);

O2A1O1Ixp33_ASAP7_75t_L g2723 ( 
.A1(n_2601),
.A2(n_1616),
.B(n_1626),
.C(n_1596),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2618),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2584),
.A2(n_1144),
.B(n_1070),
.Y(n_2725)
);

OAI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2595),
.A2(n_1673),
.B1(n_1679),
.B2(n_1639),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2640),
.B(n_2513),
.Y(n_2727)
);

AOI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2652),
.A2(n_1144),
.B(n_1070),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2619),
.B(n_2309),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2619),
.B(n_2221),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2626),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2606),
.B(n_2537),
.Y(n_2732)
);

INVx4_ASAP7_75t_L g2733 ( 
.A(n_2567),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2630),
.Y(n_2734)
);

BUFx4f_ASAP7_75t_L g2735 ( 
.A(n_2615),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2624),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2598),
.B(n_2605),
.Y(n_2737)
);

AOI21x1_ASAP7_75t_L g2738 ( 
.A1(n_2636),
.A2(n_2307),
.B(n_1685),
.Y(n_2738)
);

AOI21xp5_ASAP7_75t_L g2739 ( 
.A1(n_2653),
.A2(n_1254),
.B(n_1144),
.Y(n_2739)
);

OAI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2623),
.A2(n_1703),
.B(n_1681),
.Y(n_2740)
);

OAI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2661),
.A2(n_1725),
.B(n_1708),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2714),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2702),
.A2(n_2621),
.B1(n_2633),
.B2(n_2561),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2675),
.A2(n_2268),
.B1(n_2617),
.B2(n_2281),
.Y(n_2744)
);

A2O1A1Ixp33_ASAP7_75t_L g2745 ( 
.A1(n_2723),
.A2(n_1741),
.B(n_1760),
.C(n_1740),
.Y(n_2745)
);

OAI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2659),
.A2(n_2565),
.B(n_1251),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2662),
.B(n_2691),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2690),
.B(n_2561),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2660),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2682),
.B(n_2184),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2657),
.A2(n_1369),
.B(n_1254),
.Y(n_2751)
);

BUFx12f_ASAP7_75t_SL g2752 ( 
.A(n_2667),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2663),
.A2(n_1369),
.B(n_1254),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2695),
.B(n_2636),
.Y(n_2754)
);

INVx1_ASAP7_75t_SL g2755 ( 
.A(n_2709),
.Y(n_2755)
);

A2O1A1Ixp33_ASAP7_75t_L g2756 ( 
.A1(n_2669),
.A2(n_2257),
.B(n_2270),
.C(n_2240),
.Y(n_2756)
);

AO21x1_ASAP7_75t_L g2757 ( 
.A1(n_2670),
.A2(n_1226),
.B(n_1224),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2665),
.B(n_2606),
.Y(n_2758)
);

A2O1A1Ixp33_ASAP7_75t_L g2759 ( 
.A1(n_2668),
.A2(n_2282),
.B(n_2298),
.C(n_2275),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2674),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2679),
.B(n_2146),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_SL g2762 ( 
.A(n_2658),
.B(n_2183),
.Y(n_2762)
);

A2O1A1Ixp33_ASAP7_75t_SL g2763 ( 
.A1(n_2740),
.A2(n_2150),
.B(n_2149),
.C(n_1245),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2666),
.B(n_2429),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2706),
.B(n_2461),
.Y(n_2765)
);

AOI222xp33_ASAP7_75t_L g2766 ( 
.A1(n_2673),
.A2(n_1677),
.B1(n_1421),
.B2(n_1710),
.C1(n_1430),
.C2(n_1365),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2683),
.Y(n_2767)
);

OAI21x1_ASAP7_75t_L g2768 ( 
.A1(n_2721),
.A2(n_2716),
.B(n_2681),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2708),
.B(n_2541),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2715),
.A2(n_1683),
.B(n_1369),
.Y(n_2770)
);

CKINVDCx16_ASAP7_75t_R g2771 ( 
.A(n_2705),
.Y(n_2771)
);

O2A1O1Ixp33_ASAP7_75t_L g2772 ( 
.A1(n_2729),
.A2(n_1263),
.B(n_1267),
.C(n_1236),
.Y(n_2772)
);

OAI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2711),
.A2(n_2525),
.B1(n_1252),
.B2(n_1262),
.Y(n_2773)
);

A2O1A1Ixp33_ASAP7_75t_L g2774 ( 
.A1(n_2677),
.A2(n_1269),
.B(n_1288),
.C(n_1285),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2712),
.B(n_2541),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2720),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2680),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2710),
.A2(n_1736),
.B(n_1683),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2686),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2717),
.A2(n_1736),
.B(n_1683),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2688),
.A2(n_2637),
.B1(n_2212),
.B2(n_2344),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2696),
.B(n_1248),
.Y(n_2782)
);

OAI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2664),
.A2(n_1274),
.B1(n_1282),
.B2(n_1270),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2697),
.B(n_1365),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2692),
.A2(n_1289),
.B1(n_1290),
.B2(n_1284),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2707),
.B(n_1292),
.Y(n_2786)
);

A2O1A1Ixp33_ASAP7_75t_L g2787 ( 
.A1(n_2693),
.A2(n_1314),
.B(n_1325),
.C(n_1291),
.Y(n_2787)
);

AND2x2_ASAP7_75t_SL g2788 ( 
.A(n_2735),
.B(n_1736),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2687),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2724),
.B(n_1354),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2736),
.Y(n_2791)
);

AOI22xp33_ASAP7_75t_SL g2792 ( 
.A1(n_2732),
.A2(n_1430),
.B1(n_1710),
.B2(n_1677),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2719),
.B(n_1156),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2703),
.B(n_2730),
.C(n_2676),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2734),
.B(n_1421),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2699),
.B(n_1297),
.Y(n_2796)
);

CKINVDCx20_ASAP7_75t_R g2797 ( 
.A(n_2671),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2685),
.A2(n_1302),
.B1(n_1305),
.B2(n_1298),
.Y(n_2798)
);

AOI21x1_ASAP7_75t_L g2799 ( 
.A1(n_2738),
.A2(n_1395),
.B(n_1392),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2698),
.Y(n_2800)
);

A2O1A1Ixp33_ASAP7_75t_L g2801 ( 
.A1(n_2713),
.A2(n_1399),
.B(n_1402),
.C(n_1398),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2704),
.B(n_2689),
.Y(n_2802)
);

AOI22xp5_ASAP7_75t_L g2803 ( 
.A1(n_2718),
.A2(n_1762),
.B1(n_1313),
.B2(n_1315),
.Y(n_2803)
);

O2A1O1Ixp33_ASAP7_75t_L g2804 ( 
.A1(n_2727),
.A2(n_1413),
.B(n_1420),
.C(n_1411),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2731),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2779),
.Y(n_2806)
);

INVxp67_ASAP7_75t_SL g2807 ( 
.A(n_2776),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2755),
.Y(n_2808)
);

BUFx3_ASAP7_75t_L g2809 ( 
.A(n_2797),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2742),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2749),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2805),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2760),
.Y(n_2813)
);

INVxp67_ASAP7_75t_SL g2814 ( 
.A(n_2747),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2767),
.Y(n_2815)
);

INVx3_ASAP7_75t_SL g2816 ( 
.A(n_2771),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2789),
.Y(n_2817)
);

BUFx2_ASAP7_75t_L g2818 ( 
.A(n_2752),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_2790),
.Y(n_2819)
);

INVx8_ASAP7_75t_L g2820 ( 
.A(n_2790),
.Y(n_2820)
);

BUFx2_ASAP7_75t_SL g2821 ( 
.A(n_2791),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2758),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2748),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2801),
.Y(n_2824)
);

INVx8_ASAP7_75t_L g2825 ( 
.A(n_2795),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2775),
.Y(n_2826)
);

INVxp33_ASAP7_75t_L g2827 ( 
.A(n_2754),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2766),
.A2(n_2726),
.B1(n_2701),
.B2(n_2739),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2802),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2800),
.B(n_2684),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2793),
.B(n_2694),
.Y(n_2831)
);

HB1xp67_ASAP7_75t_L g2832 ( 
.A(n_2794),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_2744),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2777),
.Y(n_2834)
);

BUFx6f_ASAP7_75t_L g2835 ( 
.A(n_2788),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2761),
.Y(n_2836)
);

BUFx2_ASAP7_75t_SL g2837 ( 
.A(n_2750),
.Y(n_2837)
);

BUFx12f_ASAP7_75t_L g2838 ( 
.A(n_2781),
.Y(n_2838)
);

INVx4_ASAP7_75t_L g2839 ( 
.A(n_2759),
.Y(n_2839)
);

INVx5_ASAP7_75t_SL g2840 ( 
.A(n_2764),
.Y(n_2840)
);

CKINVDCx11_ASAP7_75t_R g2841 ( 
.A(n_2743),
.Y(n_2841)
);

NAND2x1p5_ASAP7_75t_L g2842 ( 
.A(n_2762),
.B(n_2678),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2765),
.Y(n_2843)
);

BUFx3_ASAP7_75t_L g2844 ( 
.A(n_2769),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2784),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2756),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2782),
.B(n_2700),
.Y(n_2847)
);

INVx4_ASAP7_75t_L g2848 ( 
.A(n_2787),
.Y(n_2848)
);

INVx2_ASAP7_75t_SL g2849 ( 
.A(n_2796),
.Y(n_2849)
);

AND2x4_ASAP7_75t_L g2850 ( 
.A(n_2774),
.B(n_2678),
.Y(n_2850)
);

INVx6_ASAP7_75t_L g2851 ( 
.A(n_2792),
.Y(n_2851)
);

CKINVDCx11_ASAP7_75t_R g2852 ( 
.A(n_2773),
.Y(n_2852)
);

BUFx2_ASAP7_75t_SL g2853 ( 
.A(n_2757),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2783),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2803),
.B(n_2672),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2799),
.Y(n_2856)
);

BUFx3_ASAP7_75t_L g2857 ( 
.A(n_2786),
.Y(n_2857)
);

HB1xp67_ASAP7_75t_L g2858 ( 
.A(n_2746),
.Y(n_2858)
);

BUFx4f_ASAP7_75t_SL g2859 ( 
.A(n_2804),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_2768),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2785),
.Y(n_2861)
);

CKINVDCx11_ASAP7_75t_R g2862 ( 
.A(n_2798),
.Y(n_2862)
);

BUFx6f_ASAP7_75t_SL g2863 ( 
.A(n_2772),
.Y(n_2863)
);

BUFx12f_ASAP7_75t_L g2864 ( 
.A(n_2763),
.Y(n_2864)
);

INVx3_ASAP7_75t_L g2865 ( 
.A(n_2770),
.Y(n_2865)
);

NAND2x1p5_ASAP7_75t_L g2866 ( 
.A(n_2778),
.B(n_2678),
.Y(n_2866)
);

OAI211xp5_ASAP7_75t_SL g2867 ( 
.A1(n_2841),
.A2(n_2741),
.B(n_1424),
.C(n_1427),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2814),
.B(n_2737),
.Y(n_2868)
);

OAI22xp33_ASAP7_75t_SL g2869 ( 
.A1(n_2851),
.A2(n_2753),
.B1(n_1429),
.B2(n_1434),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2836),
.B(n_2745),
.Y(n_2870)
);

INVx4_ASAP7_75t_L g2871 ( 
.A(n_2825),
.Y(n_2871)
);

OA21x2_ASAP7_75t_L g2872 ( 
.A1(n_2856),
.A2(n_2751),
.B(n_2780),
.Y(n_2872)
);

OR2x2_ASAP7_75t_L g2873 ( 
.A(n_2823),
.B(n_2672),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2831),
.B(n_2733),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2829),
.B(n_1763),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2827),
.B(n_1253),
.Y(n_2876)
);

OAI21x1_ASAP7_75t_L g2877 ( 
.A1(n_2865),
.A2(n_2722),
.B(n_2728),
.Y(n_2877)
);

OAI21x1_ASAP7_75t_L g2878 ( 
.A1(n_2846),
.A2(n_2725),
.B(n_1438),
.Y(n_2878)
);

AND2x4_ASAP7_75t_L g2879 ( 
.A(n_2808),
.B(n_704),
.Y(n_2879)
);

CKINVDCx20_ASAP7_75t_R g2880 ( 
.A(n_2816),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2810),
.Y(n_2881)
);

AOI221xp5_ASAP7_75t_L g2882 ( 
.A1(n_2863),
.A2(n_1166),
.B1(n_1169),
.B2(n_1161),
.C(n_1157),
.Y(n_2882)
);

INVx6_ASAP7_75t_L g2883 ( 
.A(n_2820),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2812),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2815),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2807),
.B(n_1745),
.Y(n_2886)
);

BUFx3_ASAP7_75t_L g2887 ( 
.A(n_2818),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2817),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2811),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2854),
.B(n_1309),
.Y(n_2890)
);

O2A1O1Ixp33_ASAP7_75t_SL g2891 ( 
.A1(n_2858),
.A2(n_1439),
.B(n_1446),
.C(n_1423),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_L g2892 ( 
.A1(n_2866),
.A2(n_1461),
.B(n_1452),
.Y(n_2892)
);

AOI21xp33_ASAP7_75t_SL g2893 ( 
.A1(n_2845),
.A2(n_1756),
.B(n_1172),
.Y(n_2893)
);

CKINVDCx16_ASAP7_75t_R g2894 ( 
.A(n_2809),
.Y(n_2894)
);

OAI21x1_ASAP7_75t_SL g2895 ( 
.A1(n_2834),
.A2(n_1361),
.B(n_1326),
.Y(n_2895)
);

OAI21x1_ASAP7_75t_L g2896 ( 
.A1(n_2813),
.A2(n_1472),
.B(n_1462),
.Y(n_2896)
);

AOI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_2859),
.A2(n_1722),
.B1(n_1752),
.B2(n_1726),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2806),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2843),
.A2(n_1175),
.B1(n_1176),
.B2(n_1170),
.Y(n_2899)
);

AOI21x1_ASAP7_75t_L g2900 ( 
.A1(n_2832),
.A2(n_1489),
.B(n_1474),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2822),
.Y(n_2901)
);

OAI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2828),
.A2(n_1536),
.B(n_1518),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2847),
.A2(n_1320),
.B(n_1316),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2862),
.A2(n_2852),
.B1(n_2848),
.B2(n_2861),
.Y(n_2904)
);

BUFx2_ASAP7_75t_L g2905 ( 
.A(n_2844),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2849),
.B(n_1754),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2857),
.B(n_1757),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2821),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2853),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2806),
.Y(n_2910)
);

OAI21x1_ASAP7_75t_L g2911 ( 
.A1(n_2824),
.A2(n_1494),
.B(n_1492),
.Y(n_2911)
);

A2O1A1Ixp33_ASAP7_75t_L g2912 ( 
.A1(n_2833),
.A2(n_1509),
.B(n_1517),
.C(n_1504),
.Y(n_2912)
);

OAI21x1_ASAP7_75t_L g2913 ( 
.A1(n_2842),
.A2(n_1542),
.B(n_1539),
.Y(n_2913)
);

OAI21x1_ASAP7_75t_L g2914 ( 
.A1(n_2860),
.A2(n_1575),
.B(n_1572),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2837),
.B(n_1742),
.Y(n_2915)
);

AOI221xp5_ASAP7_75t_L g2916 ( 
.A1(n_2835),
.A2(n_1199),
.B1(n_1202),
.B2(n_1192),
.C(n_1179),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2826),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2835),
.A2(n_1205),
.B1(n_1208),
.B2(n_1204),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2819),
.B(n_705),
.Y(n_2919)
);

OAI21x1_ASAP7_75t_L g2920 ( 
.A1(n_2855),
.A2(n_1592),
.B(n_1589),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2838),
.B(n_1334),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2888),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2885),
.Y(n_2923)
);

INVx4_ASAP7_75t_L g2924 ( 
.A(n_2898),
.Y(n_2924)
);

INVx4_ASAP7_75t_L g2925 ( 
.A(n_2883),
.Y(n_2925)
);

AO21x2_ASAP7_75t_L g2926 ( 
.A1(n_2909),
.A2(n_2850),
.B(n_1604),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2889),
.Y(n_2927)
);

AO21x1_ASAP7_75t_L g2928 ( 
.A1(n_2869),
.A2(n_2839),
.B(n_1615),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2901),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2883),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2881),
.Y(n_2931)
);

AO21x1_ASAP7_75t_L g2932 ( 
.A1(n_2902),
.A2(n_1609),
.B(n_1602),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2876),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2873),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2908),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2905),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2896),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2917),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2868),
.Y(n_2939)
);

INVx3_ASAP7_75t_L g2940 ( 
.A(n_2871),
.Y(n_2940)
);

BUFx2_ASAP7_75t_SL g2941 ( 
.A(n_2880),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2874),
.B(n_2840),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2884),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2895),
.Y(n_2944)
);

OAI21x1_ASAP7_75t_L g2945 ( 
.A1(n_2877),
.A2(n_1620),
.B(n_1619),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2920),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2911),
.Y(n_2947)
);

INVx1_ASAP7_75t_SL g2948 ( 
.A(n_2887),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_2886),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2900),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2870),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2912),
.Y(n_2952)
);

BUFx10_ASAP7_75t_L g2953 ( 
.A(n_2921),
.Y(n_2953)
);

AOI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2867),
.A2(n_2864),
.B1(n_2826),
.B2(n_1726),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2872),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2914),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2892),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2894),
.B(n_2830),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2875),
.Y(n_2959)
);

INVx2_ASAP7_75t_SL g2960 ( 
.A(n_2910),
.Y(n_2960)
);

OAI21x1_ASAP7_75t_L g2961 ( 
.A1(n_2878),
.A2(n_1632),
.B(n_1630),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2879),
.Y(n_2962)
);

HB1xp67_ASAP7_75t_L g2963 ( 
.A(n_2913),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2919),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2891),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2890),
.A2(n_2897),
.B1(n_2882),
.B2(n_2904),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2907),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2899),
.Y(n_2968)
);

AO21x2_ASAP7_75t_L g2969 ( 
.A1(n_2955),
.A2(n_2903),
.B(n_2915),
.Y(n_2969)
);

INVxp67_ASAP7_75t_L g2970 ( 
.A(n_2949),
.Y(n_2970)
);

AND2x4_ASAP7_75t_L g2971 ( 
.A(n_2943),
.B(n_2936),
.Y(n_2971)
);

OR2x2_ASAP7_75t_SL g2972 ( 
.A(n_2934),
.B(n_2942),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2922),
.Y(n_2973)
);

HB1xp67_ASAP7_75t_L g2974 ( 
.A(n_2933),
.Y(n_2974)
);

NAND2xp33_ASAP7_75t_R g2975 ( 
.A(n_2940),
.B(n_2906),
.Y(n_2975)
);

INVx4_ASAP7_75t_L g2976 ( 
.A(n_2924),
.Y(n_2976)
);

CKINVDCx5p33_ASAP7_75t_R g2977 ( 
.A(n_2941),
.Y(n_2977)
);

O2A1O1Ixp33_ASAP7_75t_SL g2978 ( 
.A1(n_2959),
.A2(n_1649),
.B(n_1656),
.C(n_1643),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2927),
.Y(n_2979)
);

HB1xp67_ASAP7_75t_L g2980 ( 
.A(n_2935),
.Y(n_2980)
);

INVx1_ASAP7_75t_SL g2981 ( 
.A(n_2948),
.Y(n_2981)
);

OAI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2966),
.A2(n_2893),
.B1(n_2916),
.B2(n_2918),
.Y(n_2982)
);

AO31x2_ASAP7_75t_L g2983 ( 
.A1(n_2956),
.A2(n_1667),
.A3(n_1676),
.B(n_1666),
.Y(n_2983)
);

OR2x2_ASAP7_75t_L g2984 ( 
.A(n_2939),
.B(n_1682),
.Y(n_2984)
);

CKINVDCx16_ASAP7_75t_R g2985 ( 
.A(n_2953),
.Y(n_2985)
);

OR2x6_ASAP7_75t_L g2986 ( 
.A(n_2925),
.B(n_1684),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2923),
.Y(n_2987)
);

INVxp67_ASAP7_75t_L g2988 ( 
.A(n_2967),
.Y(n_2988)
);

BUFx3_ASAP7_75t_L g2989 ( 
.A(n_2958),
.Y(n_2989)
);

CKINVDCx16_ASAP7_75t_R g2990 ( 
.A(n_2962),
.Y(n_2990)
);

NAND2xp33_ASAP7_75t_SL g2991 ( 
.A(n_2962),
.B(n_1211),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2938),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2929),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2960),
.B(n_1698),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2930),
.Y(n_2995)
);

CKINVDCx8_ASAP7_75t_R g2996 ( 
.A(n_2964),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2931),
.Y(n_2997)
);

AND2x2_ASAP7_75t_L g2998 ( 
.A(n_2951),
.B(n_1701),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2950),
.Y(n_2999)
);

OAI221xp5_ASAP7_75t_L g3000 ( 
.A1(n_2954),
.A2(n_1716),
.B1(n_1730),
.B2(n_1706),
.C(n_1702),
.Y(n_3000)
);

OAI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2945),
.A2(n_1732),
.B(n_1586),
.Y(n_3001)
);

INVx1_ASAP7_75t_SL g3002 ( 
.A(n_2926),
.Y(n_3002)
);

CKINVDCx20_ASAP7_75t_R g3003 ( 
.A(n_2968),
.Y(n_3003)
);

AND2x4_ASAP7_75t_L g3004 ( 
.A(n_2944),
.B(n_706),
.Y(n_3004)
);

INVx3_ASAP7_75t_L g3005 ( 
.A(n_2957),
.Y(n_3005)
);

NAND2xp33_ASAP7_75t_R g3006 ( 
.A(n_2952),
.B(n_2965),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2946),
.B(n_1253),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2963),
.B(n_1253),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2937),
.B(n_1253),
.Y(n_3009)
);

NOR2xp33_ASAP7_75t_R g3010 ( 
.A(n_2947),
.B(n_0),
.Y(n_3010)
);

OR2x6_ASAP7_75t_L g3011 ( 
.A(n_2928),
.B(n_1370),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2961),
.B(n_1726),
.Y(n_3012)
);

OR2x6_ASAP7_75t_L g3013 ( 
.A(n_2932),
.B(n_1443),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2932),
.B(n_1726),
.Y(n_3014)
);

AO31x2_ASAP7_75t_L g3015 ( 
.A1(n_2956),
.A2(n_1640),
.A3(n_1641),
.B(n_1564),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2943),
.B(n_707),
.Y(n_3016)
);

NAND2xp33_ASAP7_75t_SL g3017 ( 
.A(n_2924),
.B(n_1213),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2932),
.A2(n_1726),
.B1(n_1739),
.B2(n_1697),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2922),
.Y(n_3019)
);

NAND2xp33_ASAP7_75t_R g3020 ( 
.A(n_2940),
.B(n_1),
.Y(n_3020)
);

NOR3xp33_ASAP7_75t_SL g3021 ( 
.A(n_2968),
.B(n_1750),
.C(n_1749),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2943),
.B(n_1747),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2943),
.B(n_1722),
.Y(n_3023)
);

CKINVDCx16_ASAP7_75t_R g3024 ( 
.A(n_2941),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2935),
.Y(n_3025)
);

AO31x2_ASAP7_75t_L g3026 ( 
.A1(n_2956),
.A2(n_1752),
.A3(n_4),
.B(n_2),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2970),
.B(n_3),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2988),
.B(n_1215),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2973),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2992),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2979),
.Y(n_3031)
);

INVx2_ASAP7_75t_SL g3032 ( 
.A(n_2989),
.Y(n_3032)
);

BUFx6f_ASAP7_75t_L g3033 ( 
.A(n_2995),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2980),
.B(n_4),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2999),
.B(n_5),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_3019),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2987),
.B(n_1222),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_3025),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2971),
.B(n_5),
.Y(n_3039)
);

OR2x2_ASAP7_75t_L g3040 ( 
.A(n_2974),
.B(n_6),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2972),
.B(n_6),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_3024),
.B(n_7),
.Y(n_3042)
);

OAI22xp5_ASAP7_75t_SL g3043 ( 
.A1(n_2985),
.A2(n_1231),
.B1(n_1238),
.B2(n_1223),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2993),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2997),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_3008),
.B(n_1239),
.Y(n_3046)
);

INVx3_ASAP7_75t_L g3047 ( 
.A(n_2976),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_3007),
.B(n_1261),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_3009),
.B(n_1264),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_3005),
.Y(n_3050)
);

OR2x2_ASAP7_75t_L g3051 ( 
.A(n_2981),
.B(n_7),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2996),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2990),
.B(n_9),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_3022),
.B(n_1266),
.Y(n_3054)
);

OAI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_3006),
.A2(n_1271),
.B1(n_1276),
.B2(n_1268),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2984),
.Y(n_3056)
);

BUFx2_ASAP7_75t_L g3057 ( 
.A(n_2977),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_3026),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_3003),
.B(n_10),
.Y(n_3059)
);

BUFx2_ASAP7_75t_L g3060 ( 
.A(n_3010),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_3015),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_3023),
.B(n_10),
.Y(n_3062)
);

NAND2x1_ASAP7_75t_L g3063 ( 
.A(n_2998),
.B(n_11),
.Y(n_3063)
);

OAI31xp33_ASAP7_75t_L g3064 ( 
.A1(n_2982),
.A2(n_15),
.A3(n_11),
.B(n_12),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_3015),
.Y(n_3065)
);

OR2x2_ASAP7_75t_L g3066 ( 
.A(n_3002),
.B(n_12),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2983),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2994),
.B(n_16),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2983),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2969),
.B(n_3014),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_3026),
.Y(n_3071)
);

OR2x2_ASAP7_75t_L g3072 ( 
.A(n_3012),
.B(n_2986),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3016),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2978),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_2975),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3001),
.Y(n_3076)
);

NOR2x1_ASAP7_75t_SL g3077 ( 
.A(n_3013),
.B(n_2078),
.Y(n_3077)
);

OR2x2_ASAP7_75t_L g3078 ( 
.A(n_2986),
.B(n_16),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_3004),
.Y(n_3079)
);

AND2x4_ASAP7_75t_L g3080 ( 
.A(n_3011),
.B(n_17),
.Y(n_3080)
);

OR2x2_ASAP7_75t_L g3081 ( 
.A(n_3013),
.B(n_18),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_3011),
.B(n_19),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3018),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_3075),
.A2(n_3000),
.B1(n_2991),
.B2(n_3017),
.Y(n_3084)
);

A2O1A1Ixp33_ASAP7_75t_L g3085 ( 
.A1(n_3064),
.A2(n_3021),
.B(n_3020),
.C(n_1350),
.Y(n_3085)
);

AOI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_3070),
.A2(n_1351),
.B(n_1301),
.Y(n_3086)
);

OAI21x1_ASAP7_75t_L g3087 ( 
.A1(n_3071),
.A2(n_20),
.B(n_21),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_3045),
.B(n_20),
.Y(n_3088)
);

OAI22xp5_ASAP7_75t_SL g3089 ( 
.A1(n_3060),
.A2(n_1279),
.B1(n_1280),
.B2(n_1277),
.Y(n_3089)
);

BUFx3_ASAP7_75t_L g3090 ( 
.A(n_3057),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_3032),
.B(n_21),
.Y(n_3091)
);

BUFx2_ASAP7_75t_L g3092 ( 
.A(n_3052),
.Y(n_3092)
);

HB1xp67_ASAP7_75t_L g3093 ( 
.A(n_3058),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_3056),
.B(n_1293),
.Y(n_3094)
);

AOI221xp5_ASAP7_75t_L g3095 ( 
.A1(n_3055),
.A2(n_1307),
.B1(n_1308),
.B2(n_1300),
.C(n_1295),
.Y(n_3095)
);

BUFx3_ASAP7_75t_L g3096 ( 
.A(n_3033),
.Y(n_3096)
);

HB1xp67_ASAP7_75t_L g3097 ( 
.A(n_3030),
.Y(n_3097)
);

AOI221xp5_ASAP7_75t_L g3098 ( 
.A1(n_3043),
.A2(n_1328),
.B1(n_1336),
.B2(n_1323),
.C(n_1310),
.Y(n_3098)
);

AND2x4_ASAP7_75t_L g3099 ( 
.A(n_3079),
.B(n_22),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3029),
.Y(n_3100)
);

OAI31xp33_ASAP7_75t_SL g3101 ( 
.A1(n_3059),
.A2(n_3042),
.A3(n_3053),
.B(n_3039),
.Y(n_3101)
);

INVx3_ASAP7_75t_L g3102 ( 
.A(n_3033),
.Y(n_3102)
);

AOI22xp33_ASAP7_75t_L g3103 ( 
.A1(n_3083),
.A2(n_3072),
.B1(n_3074),
.B2(n_3076),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3031),
.Y(n_3104)
);

BUFx2_ASAP7_75t_L g3105 ( 
.A(n_3047),
.Y(n_3105)
);

OR2x2_ASAP7_75t_SL g3106 ( 
.A(n_3041),
.B(n_3066),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_3077),
.A2(n_1348),
.B(n_1337),
.Y(n_3107)
);

OA21x2_ASAP7_75t_L g3108 ( 
.A1(n_3036),
.A2(n_1343),
.B(n_1341),
.Y(n_3108)
);

NAND2x1_ASAP7_75t_L g3109 ( 
.A(n_3050),
.B(n_22),
.Y(n_3109)
);

A2O1A1Ixp33_ASAP7_75t_L g3110 ( 
.A1(n_3063),
.A2(n_1419),
.B(n_1465),
.C(n_1396),
.Y(n_3110)
);

BUFx3_ASAP7_75t_L g3111 ( 
.A(n_3062),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3044),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3038),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_3034),
.B(n_3046),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3035),
.Y(n_3115)
);

BUFx3_ASAP7_75t_L g3116 ( 
.A(n_3051),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_3073),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3040),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_3027),
.Y(n_3119)
);

OAI21x1_ASAP7_75t_L g3120 ( 
.A1(n_3067),
.A2(n_23),
.B(n_24),
.Y(n_3120)
);

HB1xp67_ASAP7_75t_L g3121 ( 
.A(n_3069),
.Y(n_3121)
);

AO21x2_ASAP7_75t_L g3122 ( 
.A1(n_3061),
.A2(n_23),
.B(n_24),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3065),
.Y(n_3123)
);

AOI221xp5_ASAP7_75t_L g3124 ( 
.A1(n_3082),
.A2(n_1358),
.B1(n_1362),
.B2(n_1347),
.C(n_1345),
.Y(n_3124)
);

AO21x2_ASAP7_75t_L g3125 ( 
.A1(n_3028),
.A2(n_3037),
.B(n_3048),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_3049),
.Y(n_3126)
);

OAI21x1_ASAP7_75t_L g3127 ( 
.A1(n_3081),
.A2(n_25),
.B(n_26),
.Y(n_3127)
);

OAI21x1_ASAP7_75t_L g3128 ( 
.A1(n_3054),
.A2(n_27),
.B(n_28),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_3068),
.Y(n_3129)
);

AND4x1_ASAP7_75t_L g3130 ( 
.A(n_3078),
.B(n_3080),
.C(n_29),
.D(n_27),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_3031),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_3075),
.A2(n_1374),
.B1(n_1376),
.B2(n_1367),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_3056),
.B(n_1381),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3029),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_3031),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3029),
.Y(n_3136)
);

OAI211xp5_ASAP7_75t_L g3137 ( 
.A1(n_3064),
.A2(n_1386),
.B(n_1388),
.C(n_1382),
.Y(n_3137)
);

AND2x4_ASAP7_75t_L g3138 ( 
.A(n_3056),
.B(n_28),
.Y(n_3138)
);

BUFx2_ASAP7_75t_L g3139 ( 
.A(n_3075),
.Y(n_3139)
);

OAI21x1_ASAP7_75t_L g3140 ( 
.A1(n_3071),
.A2(n_29),
.B(n_30),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_3056),
.B(n_1393),
.Y(n_3141)
);

A2O1A1Ixp33_ASAP7_75t_L g3142 ( 
.A1(n_3064),
.A2(n_1410),
.B(n_1458),
.C(n_1437),
.Y(n_3142)
);

BUFx2_ASAP7_75t_L g3143 ( 
.A(n_3075),
.Y(n_3143)
);

AND2x4_ASAP7_75t_L g3144 ( 
.A(n_3056),
.B(n_30),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_3032),
.B(n_31),
.Y(n_3145)
);

INVxp67_ASAP7_75t_L g3146 ( 
.A(n_3075),
.Y(n_3146)
);

AO31x2_ASAP7_75t_L g3147 ( 
.A1(n_3071),
.A2(n_34),
.A3(n_31),
.B(n_32),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_3056),
.B(n_32),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3031),
.Y(n_3149)
);

OAI21x1_ASAP7_75t_L g3150 ( 
.A1(n_3071),
.A2(n_35),
.B(n_36),
.Y(n_3150)
);

INVx2_ASAP7_75t_SL g3151 ( 
.A(n_3033),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3029),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_3031),
.Y(n_3153)
);

INVx2_ASAP7_75t_SL g3154 ( 
.A(n_3033),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3029),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_3058),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_3031),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_3029),
.Y(n_3158)
);

BUFx8_ASAP7_75t_L g3159 ( 
.A(n_3053),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3029),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_3070),
.A2(n_1478),
.B(n_1431),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_3032),
.B(n_36),
.Y(n_3162)
);

AO31x2_ASAP7_75t_L g3163 ( 
.A1(n_3071),
.A2(n_39),
.A3(n_37),
.B(n_38),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_3075),
.A2(n_1412),
.B1(n_1416),
.B2(n_1403),
.Y(n_3164)
);

INVx2_ASAP7_75t_SL g3165 ( 
.A(n_3033),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3029),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_3058),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_3075),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_3056),
.B(n_1422),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_3031),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_3031),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_3031),
.Y(n_3172)
);

OAI211xp5_ASAP7_75t_L g3173 ( 
.A1(n_3064),
.A2(n_1444),
.B(n_1447),
.C(n_1425),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_3031),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3029),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3031),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_3075),
.Y(n_3177)
);

INVx4_ASAP7_75t_L g3178 ( 
.A(n_3033),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_3075),
.A2(n_1453),
.B1(n_1466),
.B2(n_1449),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3032),
.B(n_38),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_3031),
.Y(n_3181)
);

BUFx2_ASAP7_75t_L g3182 ( 
.A(n_3075),
.Y(n_3182)
);

BUFx6f_ASAP7_75t_L g3183 ( 
.A(n_3033),
.Y(n_3183)
);

INVxp67_ASAP7_75t_L g3184 ( 
.A(n_3075),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3029),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3029),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_3032),
.B(n_40),
.Y(n_3187)
);

OAI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_3075),
.A2(n_1470),
.B(n_1469),
.Y(n_3188)
);

A2O1A1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_3064),
.A2(n_1508),
.B(n_1521),
.C(n_1480),
.Y(n_3189)
);

INVxp67_ASAP7_75t_SL g3190 ( 
.A(n_3075),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_3056),
.B(n_1476),
.Y(n_3191)
);

OA21x2_ASAP7_75t_L g3192 ( 
.A1(n_3075),
.A2(n_1481),
.B(n_1479),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3029),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_3070),
.A2(n_1543),
.B(n_1527),
.Y(n_3194)
);

OAI222xp33_ASAP7_75t_L g3195 ( 
.A1(n_3146),
.A2(n_3184),
.B1(n_3177),
.B2(n_3139),
.C1(n_3182),
.C2(n_3168),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3100),
.Y(n_3196)
);

HB1xp67_ASAP7_75t_L g3197 ( 
.A(n_3143),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3190),
.B(n_40),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_3092),
.B(n_41),
.Y(n_3199)
);

BUFx2_ASAP7_75t_L g3200 ( 
.A(n_3105),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3131),
.Y(n_3201)
);

INVx2_ASAP7_75t_SL g3202 ( 
.A(n_3090),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_3135),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_3149),
.Y(n_3204)
);

AOI222xp33_ASAP7_75t_L g3205 ( 
.A1(n_3085),
.A2(n_1507),
.B1(n_1490),
.B2(n_1510),
.C1(n_1499),
.C2(n_1485),
.Y(n_3205)
);

XNOR2xp5_ASAP7_75t_L g3206 ( 
.A(n_3130),
.B(n_41),
.Y(n_3206)
);

BUFx3_ASAP7_75t_L g3207 ( 
.A(n_3159),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3134),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3119),
.B(n_42),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3136),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3152),
.Y(n_3211)
);

AO21x2_ASAP7_75t_L g3212 ( 
.A1(n_3093),
.A2(n_43),
.B(n_44),
.Y(n_3212)
);

BUFx3_ASAP7_75t_L g3213 ( 
.A(n_3096),
.Y(n_3213)
);

OR2x2_ASAP7_75t_L g3214 ( 
.A(n_3106),
.B(n_43),
.Y(n_3214)
);

INVxp67_ASAP7_75t_SL g3215 ( 
.A(n_3109),
.Y(n_3215)
);

AOI211xp5_ASAP7_75t_L g3216 ( 
.A1(n_3194),
.A2(n_3161),
.B(n_3086),
.C(n_3137),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3117),
.B(n_44),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3155),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3125),
.B(n_1513),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3116),
.B(n_45),
.Y(n_3220)
);

INVxp67_ASAP7_75t_SL g3221 ( 
.A(n_3192),
.Y(n_3221)
);

BUFx2_ASAP7_75t_L g3222 ( 
.A(n_3178),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_L g3223 ( 
.A1(n_3126),
.A2(n_1520),
.B1(n_1523),
.B2(n_1514),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3158),
.Y(n_3224)
);

BUFx2_ASAP7_75t_L g3225 ( 
.A(n_3183),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3103),
.B(n_45),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3153),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3188),
.A2(n_1526),
.B1(n_1528),
.B2(n_1524),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3115),
.B(n_46),
.Y(n_3229)
);

AND2x2_ASAP7_75t_L g3230 ( 
.A(n_3118),
.B(n_47),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3157),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_3170),
.Y(n_3232)
);

NAND2xp33_ASAP7_75t_R g3233 ( 
.A(n_3108),
.B(n_47),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3160),
.Y(n_3234)
);

NAND3xp33_ASAP7_75t_L g3235 ( 
.A(n_3142),
.B(n_1531),
.C(n_1529),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_3114),
.B(n_1533),
.Y(n_3236)
);

OR2x6_ASAP7_75t_L g3237 ( 
.A(n_3183),
.B(n_48),
.Y(n_3237)
);

INVx1_ASAP7_75t_SL g3238 ( 
.A(n_3102),
.Y(n_3238)
);

HB1xp67_ASAP7_75t_L g3239 ( 
.A(n_3156),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_3097),
.B(n_48),
.Y(n_3240)
);

HB1xp67_ASAP7_75t_L g3241 ( 
.A(n_3167),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3171),
.Y(n_3242)
);

OR2x2_ASAP7_75t_L g3243 ( 
.A(n_3113),
.B(n_49),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3172),
.B(n_49),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_3174),
.Y(n_3245)
);

OAI31xp33_ASAP7_75t_SL g3246 ( 
.A1(n_3173),
.A2(n_53),
.A3(n_50),
.B(n_51),
.Y(n_3246)
);

NAND2x1_ASAP7_75t_L g3247 ( 
.A(n_3176),
.B(n_53),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3181),
.B(n_51),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_3084),
.A2(n_1541),
.B1(n_1544),
.B2(n_1534),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_3166),
.Y(n_3250)
);

HB1xp67_ASAP7_75t_L g3251 ( 
.A(n_3175),
.Y(n_3251)
);

BUFx2_ASAP7_75t_L g3252 ( 
.A(n_3111),
.Y(n_3252)
);

O2A1O1Ixp5_ASAP7_75t_L g3253 ( 
.A1(n_3104),
.A2(n_57),
.B(n_54),
.C(n_55),
.Y(n_3253)
);

INVx2_ASAP7_75t_SL g3254 ( 
.A(n_3151),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3185),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3112),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3186),
.Y(n_3257)
);

HB1xp67_ASAP7_75t_L g3258 ( 
.A(n_3193),
.Y(n_3258)
);

BUFx2_ASAP7_75t_L g3259 ( 
.A(n_3154),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3165),
.B(n_54),
.Y(n_3260)
);

OAI211xp5_ASAP7_75t_SL g3261 ( 
.A1(n_3132),
.A2(n_3164),
.B(n_3179),
.C(n_3101),
.Y(n_3261)
);

OR2x2_ASAP7_75t_L g3262 ( 
.A(n_3088),
.B(n_55),
.Y(n_3262)
);

INVx3_ASAP7_75t_L g3263 ( 
.A(n_3138),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3123),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3144),
.B(n_57),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3121),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3148),
.B(n_60),
.Y(n_3267)
);

NAND3xp33_ASAP7_75t_SL g3268 ( 
.A(n_3189),
.B(n_1549),
.C(n_1548),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3147),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3147),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3163),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_3094),
.B(n_1551),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3091),
.B(n_60),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3133),
.B(n_1552),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3099),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3163),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3145),
.B(n_61),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3162),
.B(n_62),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3141),
.Y(n_3279)
);

OAI211xp5_ASAP7_75t_L g3280 ( 
.A1(n_3098),
.A2(n_1555),
.B(n_1562),
.C(n_1554),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3169),
.B(n_1568),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_3127),
.B(n_63),
.Y(n_3282)
);

AO31x2_ASAP7_75t_L g3283 ( 
.A1(n_3191),
.A2(n_65),
.A3(n_63),
.B(n_64),
.Y(n_3283)
);

HB1xp67_ASAP7_75t_L g3284 ( 
.A(n_3122),
.Y(n_3284)
);

NOR2xp33_ASAP7_75t_L g3285 ( 
.A(n_3089),
.B(n_1570),
.Y(n_3285)
);

OAI211xp5_ASAP7_75t_L g3286 ( 
.A1(n_3124),
.A2(n_3095),
.B(n_3110),
.C(n_3107),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3180),
.B(n_1571),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3187),
.B(n_66),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3087),
.Y(n_3289)
);

HB1xp67_ASAP7_75t_L g3290 ( 
.A(n_3150),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3140),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3120),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3129),
.B(n_66),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3128),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3139),
.B(n_67),
.Y(n_3295)
);

BUFx2_ASAP7_75t_SL g3296 ( 
.A(n_3090),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3100),
.Y(n_3297)
);

BUFx2_ASAP7_75t_L g3298 ( 
.A(n_3139),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3139),
.B(n_68),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3139),
.B(n_68),
.Y(n_3300)
);

BUFx2_ASAP7_75t_L g3301 ( 
.A(n_3139),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3092),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3100),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3125),
.B(n_1574),
.Y(n_3304)
);

AND4x1_ASAP7_75t_L g3305 ( 
.A(n_3084),
.B(n_71),
.C(n_69),
.D(n_70),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3100),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3125),
.B(n_1578),
.Y(n_3307)
);

OR2x2_ASAP7_75t_L g3308 ( 
.A(n_3190),
.B(n_70),
.Y(n_3308)
);

INVx2_ASAP7_75t_SL g3309 ( 
.A(n_3090),
.Y(n_3309)
);

HB1xp67_ASAP7_75t_L g3310 ( 
.A(n_3139),
.Y(n_3310)
);

BUFx3_ASAP7_75t_L g3311 ( 
.A(n_3159),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3139),
.B(n_71),
.Y(n_3312)
);

INVxp67_ASAP7_75t_SL g3313 ( 
.A(n_3146),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3092),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3092),
.Y(n_3315)
);

AOI22xp33_ASAP7_75t_SL g3316 ( 
.A1(n_3190),
.A2(n_1723),
.B1(n_1729),
.B2(n_1718),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3100),
.Y(n_3317)
);

INVx4_ASAP7_75t_L g3318 ( 
.A(n_3183),
.Y(n_3318)
);

NAND2x1_ASAP7_75t_L g3319 ( 
.A(n_3139),
.B(n_73),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_3190),
.B(n_72),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3100),
.Y(n_3321)
);

OR2x2_ASAP7_75t_L g3322 ( 
.A(n_3190),
.B(n_72),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3190),
.B(n_73),
.Y(n_3323)
);

AND2x4_ASAP7_75t_L g3324 ( 
.A(n_3092),
.B(n_75),
.Y(n_3324)
);

AOI221xp5_ASAP7_75t_L g3325 ( 
.A1(n_3194),
.A2(n_1594),
.B1(n_1597),
.B2(n_1585),
.C(n_1583),
.Y(n_3325)
);

OAI21x1_ASAP7_75t_SL g3326 ( 
.A1(n_3188),
.A2(n_75),
.B(n_76),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3092),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3139),
.B(n_76),
.Y(n_3328)
);

INVx4_ASAP7_75t_L g3329 ( 
.A(n_3183),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3139),
.B(n_77),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3139),
.B(n_77),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3100),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3139),
.B(n_79),
.Y(n_3333)
);

OR2x2_ASAP7_75t_L g3334 ( 
.A(n_3190),
.B(n_80),
.Y(n_3334)
);

BUFx2_ASAP7_75t_L g3335 ( 
.A(n_3139),
.Y(n_3335)
);

INVxp67_ASAP7_75t_SL g3336 ( 
.A(n_3146),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3100),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3190),
.B(n_81),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_3183),
.Y(n_3339)
);

INVxp67_ASAP7_75t_L g3340 ( 
.A(n_3139),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3139),
.B(n_81),
.Y(n_3341)
);

AOI31xp33_ASAP7_75t_L g3342 ( 
.A1(n_3190),
.A2(n_1605),
.A3(n_1606),
.B(n_1600),
.Y(n_3342)
);

BUFx6f_ASAP7_75t_L g3343 ( 
.A(n_3183),
.Y(n_3343)
);

NAND3xp33_ASAP7_75t_L g3344 ( 
.A(n_3086),
.B(n_1611),
.C(n_1608),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3139),
.B(n_82),
.Y(n_3345)
);

INVxp67_ASAP7_75t_SL g3346 ( 
.A(n_3146),
.Y(n_3346)
);

AO21x2_ASAP7_75t_L g3347 ( 
.A1(n_3190),
.A2(n_82),
.B(n_83),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_3092),
.B(n_1612),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3100),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3296),
.B(n_83),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3313),
.B(n_1613),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3222),
.B(n_84),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_3336),
.B(n_84),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3250),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3251),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3200),
.B(n_85),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3346),
.B(n_1617),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3298),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3294),
.B(n_1623),
.Y(n_3359)
);

HB1xp67_ASAP7_75t_L g3360 ( 
.A(n_3197),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3302),
.B(n_85),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3258),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3314),
.B(n_3315),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_3301),
.B(n_1624),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3340),
.B(n_1625),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3327),
.B(n_86),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3252),
.B(n_86),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3196),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_3335),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3259),
.B(n_87),
.Y(n_3370)
);

AND2x4_ASAP7_75t_SL g3371 ( 
.A(n_3318),
.B(n_87),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_3207),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3225),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3310),
.B(n_3202),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3208),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3309),
.B(n_88),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3238),
.B(n_88),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3215),
.B(n_89),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3254),
.B(n_89),
.Y(n_3379)
);

AND3x1_ASAP7_75t_L g3380 ( 
.A(n_3246),
.B(n_90),
.C(n_91),
.Y(n_3380)
);

NAND2x1p5_ASAP7_75t_L g3381 ( 
.A(n_3319),
.B(n_3247),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3289),
.B(n_1628),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3279),
.B(n_90),
.Y(n_3383)
);

CKINVDCx16_ASAP7_75t_R g3384 ( 
.A(n_3311),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3291),
.B(n_1629),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3210),
.Y(n_3386)
);

NAND2x1p5_ASAP7_75t_L g3387 ( 
.A(n_3217),
.B(n_3329),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3263),
.B(n_92),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3213),
.B(n_3292),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_3275),
.B(n_92),
.Y(n_3390)
);

HB1xp67_ASAP7_75t_L g3391 ( 
.A(n_3239),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3290),
.B(n_1635),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_R g3393 ( 
.A(n_3233),
.B(n_93),
.Y(n_3393)
);

NOR4xp25_ASAP7_75t_SL g3394 ( 
.A(n_3195),
.B(n_1644),
.C(n_1645),
.D(n_1637),
.Y(n_3394)
);

OAI221xp5_ASAP7_75t_L g3395 ( 
.A1(n_3216),
.A2(n_1651),
.B1(n_1652),
.B2(n_1650),
.C(n_1646),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3229),
.B(n_93),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3339),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3221),
.B(n_1653),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3226),
.B(n_1657),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3211),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3230),
.B(n_94),
.Y(n_3401)
);

OR2x2_ASAP7_75t_L g3402 ( 
.A(n_3201),
.B(n_94),
.Y(n_3402)
);

OR2x2_ASAP7_75t_L g3403 ( 
.A(n_3203),
.B(n_95),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3214),
.B(n_1660),
.Y(n_3404)
);

NOR4xp25_ASAP7_75t_L g3405 ( 
.A(n_3261),
.B(n_100),
.C(n_98),
.D(n_99),
.Y(n_3405)
);

NOR2x1_ASAP7_75t_L g3406 ( 
.A(n_3347),
.B(n_101),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_3204),
.B(n_103),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3218),
.Y(n_3408)
);

AND2x4_ASAP7_75t_L g3409 ( 
.A(n_3339),
.B(n_104),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3198),
.B(n_1663),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3227),
.B(n_104),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3343),
.Y(n_3412)
);

AND2x4_ASAP7_75t_L g3413 ( 
.A(n_3343),
.B(n_105),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3224),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3231),
.B(n_105),
.Y(n_3415)
);

AND2x2_ASAP7_75t_L g3416 ( 
.A(n_3232),
.B(n_106),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3242),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3295),
.B(n_1664),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3234),
.Y(n_3419)
);

AND2x4_ASAP7_75t_L g3420 ( 
.A(n_3324),
.B(n_3260),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3299),
.B(n_1665),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3245),
.B(n_106),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3255),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3300),
.B(n_108),
.Y(n_3424)
);

HB1xp67_ASAP7_75t_L g3425 ( 
.A(n_3241),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3257),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3312),
.B(n_1671),
.Y(n_3427)
);

AND2x4_ASAP7_75t_L g3428 ( 
.A(n_3199),
.B(n_108),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3256),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3297),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3328),
.B(n_3330),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3303),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3331),
.B(n_110),
.Y(n_3433)
);

AND2x2_ASAP7_75t_L g3434 ( 
.A(n_3333),
.B(n_3341),
.Y(n_3434)
);

AND2x4_ASAP7_75t_SL g3435 ( 
.A(n_3237),
.B(n_111),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3306),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3317),
.Y(n_3437)
);

INVx2_ASAP7_75t_SL g3438 ( 
.A(n_3345),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_3266),
.B(n_111),
.Y(n_3439)
);

AND2x4_ASAP7_75t_L g3440 ( 
.A(n_3240),
.B(n_112),
.Y(n_3440)
);

OR2x2_ASAP7_75t_L g3441 ( 
.A(n_3321),
.B(n_112),
.Y(n_3441)
);

OR2x2_ASAP7_75t_L g3442 ( 
.A(n_3332),
.B(n_113),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_3342),
.B(n_1734),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3209),
.B(n_114),
.Y(n_3444)
);

INVx1_ASAP7_75t_SL g3445 ( 
.A(n_3308),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3219),
.B(n_1678),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3284),
.B(n_114),
.Y(n_3447)
);

BUFx2_ASAP7_75t_L g3448 ( 
.A(n_3237),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3304),
.B(n_1688),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_3269),
.B(n_3270),
.Y(n_3450)
);

AND2x4_ASAP7_75t_L g3451 ( 
.A(n_3220),
.B(n_115),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3337),
.Y(n_3452)
);

OR2x2_ASAP7_75t_L g3453 ( 
.A(n_3349),
.B(n_115),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3271),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3276),
.B(n_116),
.Y(n_3455)
);

INVxp67_ASAP7_75t_SL g3456 ( 
.A(n_3320),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3264),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3243),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3244),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3248),
.B(n_116),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3212),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3282),
.Y(n_3462)
);

HB1xp67_ASAP7_75t_L g3463 ( 
.A(n_3322),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3323),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3334),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3338),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3262),
.Y(n_3467)
);

HB1xp67_ASAP7_75t_L g3468 ( 
.A(n_3307),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3273),
.B(n_117),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3277),
.B(n_1689),
.Y(n_3470)
);

NAND2x1_ASAP7_75t_L g3471 ( 
.A(n_3293),
.B(n_117),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3283),
.Y(n_3472)
);

OR2x2_ASAP7_75t_L g3473 ( 
.A(n_3283),
.B(n_118),
.Y(n_3473)
);

HB1xp67_ASAP7_75t_L g3474 ( 
.A(n_3278),
.Y(n_3474)
);

INVxp67_ASAP7_75t_L g3475 ( 
.A(n_3348),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_3287),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3253),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3288),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3265),
.B(n_118),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3267),
.B(n_119),
.Y(n_3480)
);

INVx2_ASAP7_75t_SL g3481 ( 
.A(n_3206),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3326),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3249),
.B(n_3236),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3223),
.B(n_1690),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_3305),
.B(n_1692),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3272),
.Y(n_3486)
);

BUFx6f_ASAP7_75t_L g3487 ( 
.A(n_3274),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3281),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3316),
.B(n_120),
.Y(n_3489)
);

BUFx2_ASAP7_75t_L g3490 ( 
.A(n_3344),
.Y(n_3490)
);

NAND3xp33_ASAP7_75t_L g3491 ( 
.A(n_3325),
.B(n_1717),
.C(n_1695),
.Y(n_3491)
);

INVx4_ASAP7_75t_L g3492 ( 
.A(n_3285),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3286),
.Y(n_3493)
);

AOI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3268),
.A2(n_1696),
.B1(n_1699),
.B2(n_1694),
.Y(n_3494)
);

AND2x4_ASAP7_75t_L g3495 ( 
.A(n_3235),
.B(n_121),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3205),
.B(n_122),
.Y(n_3496)
);

HB1xp67_ASAP7_75t_L g3497 ( 
.A(n_3280),
.Y(n_3497)
);

AND2x2_ASAP7_75t_SL g3498 ( 
.A(n_3228),
.B(n_123),
.Y(n_3498)
);

AND2x4_ASAP7_75t_SL g3499 ( 
.A(n_3318),
.B(n_123),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3296),
.B(n_124),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3250),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3296),
.B(n_124),
.Y(n_3502)
);

BUFx2_ASAP7_75t_L g3503 ( 
.A(n_3298),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3222),
.B(n_125),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3250),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3222),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3313),
.B(n_1700),
.Y(n_3507)
);

INVx1_ASAP7_75t_SL g3508 ( 
.A(n_3296),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3296),
.B(n_125),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3313),
.B(n_1711),
.Y(n_3510)
);

HB1xp67_ASAP7_75t_L g3511 ( 
.A(n_3197),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3313),
.B(n_126),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3296),
.B(n_126),
.Y(n_3513)
);

AND2x4_ASAP7_75t_L g3514 ( 
.A(n_3222),
.B(n_127),
.Y(n_3514)
);

HB1xp67_ASAP7_75t_L g3515 ( 
.A(n_3197),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3313),
.B(n_1715),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3222),
.Y(n_3517)
);

INVx4_ASAP7_75t_L g3518 ( 
.A(n_3207),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3313),
.B(n_1733),
.Y(n_3519)
);

OR2x2_ASAP7_75t_L g3520 ( 
.A(n_3313),
.B(n_127),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3313),
.B(n_1737),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3313),
.B(n_1743),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3250),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_3197),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_3296),
.B(n_128),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3250),
.Y(n_3526)
);

INVxp67_ASAP7_75t_SL g3527 ( 
.A(n_3215),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3296),
.B(n_128),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3222),
.Y(n_3529)
);

INVx1_ASAP7_75t_SL g3530 ( 
.A(n_3296),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3296),
.B(n_129),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_SL g3532 ( 
.A(n_3195),
.B(n_1751),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_3296),
.B(n_129),
.Y(n_3533)
);

NOR2xp67_ASAP7_75t_L g3534 ( 
.A(n_3197),
.B(n_130),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3296),
.B(n_130),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3296),
.B(n_132),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3313),
.B(n_1759),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3296),
.B(n_132),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3222),
.Y(n_3539)
);

OR2x2_ASAP7_75t_L g3540 ( 
.A(n_3456),
.B(n_3445),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3477),
.B(n_134),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3508),
.B(n_3530),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3391),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3448),
.B(n_134),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3425),
.Y(n_3545)
);

OR2x2_ASAP7_75t_L g3546 ( 
.A(n_3463),
.B(n_135),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3527),
.B(n_136),
.Y(n_3547)
);

OAI22xp5_ASAP7_75t_L g3548 ( 
.A1(n_3380),
.A2(n_1340),
.B1(n_1342),
.B2(n_1338),
.Y(n_3548)
);

HB1xp67_ASAP7_75t_L g3549 ( 
.A(n_3503),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3454),
.Y(n_3550)
);

INVxp67_ASAP7_75t_L g3551 ( 
.A(n_3532),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3372),
.Y(n_3552)
);

OAI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_3394),
.A2(n_1357),
.B1(n_1364),
.B2(n_1353),
.Y(n_3553)
);

BUFx2_ASAP7_75t_L g3554 ( 
.A(n_3387),
.Y(n_3554)
);

NOR2xp67_ASAP7_75t_L g3555 ( 
.A(n_3518),
.B(n_136),
.Y(n_3555)
);

AND2x2_ASAP7_75t_SL g3556 ( 
.A(n_3405),
.B(n_137),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3384),
.Y(n_3557)
);

INVxp67_ASAP7_75t_L g3558 ( 
.A(n_3406),
.Y(n_3558)
);

INVxp67_ASAP7_75t_L g3559 ( 
.A(n_3360),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3381),
.Y(n_3560)
);

INVxp67_ASAP7_75t_L g3561 ( 
.A(n_3511),
.Y(n_3561)
);

AND2x2_ASAP7_75t_L g3562 ( 
.A(n_3374),
.B(n_137),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3515),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3524),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3438),
.B(n_138),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3450),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3539),
.B(n_138),
.Y(n_3567)
);

INVx1_ASAP7_75t_SL g3568 ( 
.A(n_3393),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3467),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3506),
.B(n_139),
.Y(n_3570)
);

OR2x2_ASAP7_75t_L g3571 ( 
.A(n_3474),
.B(n_3465),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3517),
.Y(n_3572)
);

AND2x2_ASAP7_75t_L g3573 ( 
.A(n_3529),
.B(n_140),
.Y(n_3573)
);

HB1xp67_ASAP7_75t_L g3574 ( 
.A(n_3534),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3373),
.B(n_140),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3358),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3458),
.Y(n_3577)
);

OAI21xp33_ASAP7_75t_SL g3578 ( 
.A1(n_3461),
.A2(n_3472),
.B(n_3493),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3369),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3478),
.B(n_142),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3389),
.B(n_143),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_SL g3582 ( 
.A1(n_3482),
.A2(n_1433),
.B1(n_1488),
.B2(n_1372),
.Y(n_3582)
);

CKINVDCx16_ASAP7_75t_R g3583 ( 
.A(n_3492),
.Y(n_3583)
);

OR2x2_ASAP7_75t_L g3584 ( 
.A(n_3462),
.B(n_143),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3397),
.B(n_3412),
.Y(n_3585)
);

INVxp67_ASAP7_75t_L g3586 ( 
.A(n_3431),
.Y(n_3586)
);

A2O1A1Ixp33_ASAP7_75t_L g3587 ( 
.A1(n_3473),
.A2(n_1371),
.B(n_1375),
.C(n_1368),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3363),
.B(n_144),
.Y(n_3588)
);

HB1xp67_ASAP7_75t_L g3589 ( 
.A(n_3464),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3459),
.B(n_144),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3434),
.B(n_3466),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3447),
.B(n_145),
.Y(n_3592)
);

INVx1_ASAP7_75t_SL g3593 ( 
.A(n_3371),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3420),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3457),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3402),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3488),
.B(n_145),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3368),
.Y(n_3598)
);

INVxp67_ASAP7_75t_SL g3599 ( 
.A(n_3471),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3375),
.Y(n_3600)
);

OR2x2_ASAP7_75t_L g3601 ( 
.A(n_3468),
.B(n_146),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3486),
.B(n_147),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3476),
.B(n_147),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3386),
.Y(n_3604)
);

OR2x2_ASAP7_75t_L g3605 ( 
.A(n_3354),
.B(n_148),
.Y(n_3605)
);

BUFx2_ASAP7_75t_L g3606 ( 
.A(n_3350),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3400),
.Y(n_3607)
);

OR2x2_ASAP7_75t_L g3608 ( 
.A(n_3355),
.B(n_148),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3500),
.B(n_149),
.Y(n_3609)
);

OR2x2_ASAP7_75t_L g3610 ( 
.A(n_3362),
.B(n_149),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3408),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3414),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3419),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3378),
.B(n_150),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3423),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3455),
.B(n_150),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3403),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3426),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3430),
.Y(n_3619)
);

HB1xp67_ASAP7_75t_L g3620 ( 
.A(n_3501),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3490),
.B(n_151),
.Y(n_3621)
);

OR2x2_ASAP7_75t_L g3622 ( 
.A(n_3505),
.B(n_151),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3432),
.Y(n_3623)
);

OAI22xp33_ASAP7_75t_SL g3624 ( 
.A1(n_3364),
.A2(n_1384),
.B1(n_1390),
.B2(n_1380),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3504),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3356),
.B(n_152),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3352),
.B(n_152),
.Y(n_3627)
);

AND2x2_ASAP7_75t_L g3628 ( 
.A(n_3502),
.B(n_153),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3436),
.Y(n_3629)
);

INVx2_ASAP7_75t_SL g3630 ( 
.A(n_3499),
.Y(n_3630)
);

OAI21xp33_ASAP7_75t_L g3631 ( 
.A1(n_3523),
.A2(n_1407),
.B(n_1400),
.Y(n_3631)
);

OR2x2_ASAP7_75t_L g3632 ( 
.A(n_3526),
.B(n_154),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3437),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3452),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3509),
.B(n_3513),
.Y(n_3635)
);

INVx4_ASAP7_75t_L g3636 ( 
.A(n_3514),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3370),
.B(n_154),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3429),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3441),
.Y(n_3639)
);

INVx4_ASAP7_75t_L g3640 ( 
.A(n_3435),
.Y(n_3640)
);

OR2x2_ASAP7_75t_L g3641 ( 
.A(n_3417),
.B(n_155),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3525),
.B(n_156),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3528),
.B(n_3531),
.Y(n_3643)
);

NAND3xp33_ASAP7_75t_SL g3644 ( 
.A(n_3485),
.B(n_1493),
.C(n_1415),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3383),
.B(n_3367),
.Y(n_3645)
);

OAI21xp33_ASAP7_75t_L g3646 ( 
.A1(n_3497),
.A2(n_1454),
.B(n_1448),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3361),
.B(n_158),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3442),
.Y(n_3648)
);

OR2x2_ASAP7_75t_L g3649 ( 
.A(n_3353),
.B(n_158),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3533),
.B(n_159),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3453),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3407),
.Y(n_3652)
);

AND3x1_ASAP7_75t_L g3653 ( 
.A(n_3535),
.B(n_160),
.C(n_161),
.Y(n_3653)
);

OR2x2_ASAP7_75t_L g3654 ( 
.A(n_3512),
.B(n_162),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3411),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3366),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3415),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_SL g3658 ( 
.A(n_3520),
.B(n_3487),
.Y(n_3658)
);

INVx2_ASAP7_75t_SL g3659 ( 
.A(n_3536),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3538),
.B(n_3439),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3416),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3422),
.Y(n_3662)
);

OR2x2_ASAP7_75t_L g3663 ( 
.A(n_3392),
.B(n_162),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3390),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3388),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3377),
.B(n_164),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3379),
.Y(n_3667)
);

INVxp67_ASAP7_75t_L g3668 ( 
.A(n_3351),
.Y(n_3668)
);

OR2x2_ASAP7_75t_L g3669 ( 
.A(n_3382),
.B(n_164),
.Y(n_3669)
);

OAI31xp33_ASAP7_75t_L g3670 ( 
.A1(n_3496),
.A2(n_167),
.A3(n_165),
.B(n_166),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3365),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3404),
.B(n_166),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3487),
.B(n_167),
.Y(n_3673)
);

INVx2_ASAP7_75t_SL g3674 ( 
.A(n_3542),
.Y(n_3674)
);

INVx2_ASAP7_75t_SL g3675 ( 
.A(n_3557),
.Y(n_3675)
);

OR2x2_ASAP7_75t_L g3676 ( 
.A(n_3540),
.B(n_3359),
.Y(n_3676)
);

INVxp67_ASAP7_75t_L g3677 ( 
.A(n_3574),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3549),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3635),
.B(n_3475),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3589),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3643),
.B(n_3376),
.Y(n_3681)
);

NAND2x1p5_ASAP7_75t_L g3682 ( 
.A(n_3653),
.B(n_3428),
.Y(n_3682)
);

AND2x2_ASAP7_75t_L g3683 ( 
.A(n_3583),
.B(n_3460),
.Y(n_3683)
);

OR2x2_ASAP7_75t_L g3684 ( 
.A(n_3606),
.B(n_3357),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3640),
.B(n_3444),
.Y(n_3685)
);

INVx1_ASAP7_75t_SL g3686 ( 
.A(n_3568),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3630),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_L g3688 ( 
.A(n_3636),
.B(n_3481),
.Y(n_3688)
);

OR2x2_ASAP7_75t_L g3689 ( 
.A(n_3571),
.B(n_3507),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3620),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3552),
.B(n_3396),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_L g3692 ( 
.A(n_3593),
.B(n_3446),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3543),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3554),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3545),
.Y(n_3695)
);

INVx1_ASAP7_75t_SL g3696 ( 
.A(n_3544),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3563),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3564),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_3551),
.B(n_3449),
.Y(n_3699)
);

OR2x6_ASAP7_75t_L g3700 ( 
.A(n_3555),
.B(n_3495),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3641),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3659),
.B(n_3401),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3599),
.B(n_3424),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3558),
.B(n_3398),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3625),
.B(n_3433),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3594),
.B(n_3585),
.Y(n_3706)
);

NAND2xp33_ASAP7_75t_L g3707 ( 
.A(n_3560),
.B(n_3510),
.Y(n_3707)
);

INVx2_ASAP7_75t_SL g3708 ( 
.A(n_3562),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3656),
.B(n_3469),
.Y(n_3709)
);

INVxp67_ASAP7_75t_L g3710 ( 
.A(n_3660),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3559),
.Y(n_3711)
);

NAND2x1p5_ASAP7_75t_L g3712 ( 
.A(n_3556),
.B(n_3409),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3586),
.B(n_3440),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3575),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3661),
.B(n_3479),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3561),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3664),
.B(n_3516),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3667),
.B(n_3519),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3591),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3550),
.Y(n_3720)
);

CKINVDCx16_ASAP7_75t_R g3721 ( 
.A(n_3644),
.Y(n_3721)
);

NAND3xp33_ASAP7_75t_L g3722 ( 
.A(n_3578),
.B(n_3491),
.C(n_3395),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3584),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3605),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3608),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3610),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3665),
.B(n_3480),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3652),
.B(n_3451),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3655),
.B(n_3521),
.Y(n_3729)
);

AND2x4_ASAP7_75t_L g3730 ( 
.A(n_3572),
.B(n_3413),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3576),
.B(n_3522),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3657),
.B(n_3537),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3579),
.B(n_3489),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3645),
.B(n_3399),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3622),
.Y(n_3735)
);

OR2x2_ASAP7_75t_L g3736 ( 
.A(n_3658),
.B(n_3385),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3662),
.B(n_3483),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3632),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3596),
.B(n_3470),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3639),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3648),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3651),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3617),
.B(n_3418),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3581),
.B(n_3410),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3546),
.Y(n_3745)
);

OAI211xp5_ASAP7_75t_L g3746 ( 
.A1(n_3670),
.A2(n_3494),
.B(n_3443),
.C(n_3484),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3668),
.B(n_3421),
.Y(n_3747)
);

OR2x2_ASAP7_75t_L g3748 ( 
.A(n_3541),
.B(n_3427),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3590),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3671),
.B(n_3498),
.Y(n_3750)
);

OAI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3547),
.A2(n_1459),
.B1(n_1460),
.B2(n_1456),
.Y(n_3751)
);

CKINVDCx16_ASAP7_75t_R g3752 ( 
.A(n_3609),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3588),
.B(n_168),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3567),
.B(n_168),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3566),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3570),
.B(n_170),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3598),
.Y(n_3757)
);

BUFx3_ASAP7_75t_L g3758 ( 
.A(n_3573),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3577),
.B(n_170),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3638),
.B(n_171),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3600),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3604),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_L g3763 ( 
.A(n_3686),
.B(n_3580),
.Y(n_3763)
);

INVx2_ASAP7_75t_SL g3764 ( 
.A(n_3685),
.Y(n_3764)
);

INVx1_ASAP7_75t_SL g3765 ( 
.A(n_3683),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3703),
.B(n_3628),
.Y(n_3766)
);

BUFx2_ASAP7_75t_L g3767 ( 
.A(n_3700),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3752),
.B(n_3621),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3678),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3674),
.B(n_3642),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3687),
.B(n_3650),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3675),
.B(n_3569),
.Y(n_3772)
);

NAND2x1p5_ASAP7_75t_L g3773 ( 
.A(n_3679),
.B(n_3601),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_SL g3774 ( 
.A(n_3682),
.B(n_3548),
.Y(n_3774)
);

INVxp33_ASAP7_75t_L g3775 ( 
.A(n_3712),
.Y(n_3775)
);

OR2x2_ASAP7_75t_L g3776 ( 
.A(n_3696),
.B(n_3595),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3677),
.Y(n_3777)
);

CKINVDCx16_ASAP7_75t_R g3778 ( 
.A(n_3721),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3680),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3681),
.B(n_3602),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3706),
.B(n_3603),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3688),
.B(n_3597),
.Y(n_3782)
);

OR2x2_ASAP7_75t_L g3783 ( 
.A(n_3684),
.B(n_3565),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3758),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3705),
.B(n_3582),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3708),
.B(n_3702),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3690),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3724),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3725),
.Y(n_3789)
);

INVxp67_ASAP7_75t_L g3790 ( 
.A(n_3700),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_L g3791 ( 
.A(n_3730),
.B(n_3669),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3726),
.Y(n_3792)
);

INVxp67_ASAP7_75t_L g3793 ( 
.A(n_3691),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3714),
.B(n_3663),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3733),
.B(n_3713),
.Y(n_3795)
);

INVxp67_ASAP7_75t_SL g3796 ( 
.A(n_3694),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3728),
.B(n_3646),
.Y(n_3797)
);

INVx1_ASAP7_75t_SL g3798 ( 
.A(n_3754),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3735),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3715),
.B(n_3607),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3745),
.B(n_3592),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3727),
.Y(n_3802)
);

INVx2_ASAP7_75t_SL g3803 ( 
.A(n_3709),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3750),
.B(n_3611),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3738),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3723),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3759),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3749),
.B(n_3701),
.Y(n_3808)
);

INVxp67_ASAP7_75t_L g3809 ( 
.A(n_3692),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3711),
.Y(n_3810)
);

INVx1_ASAP7_75t_SL g3811 ( 
.A(n_3756),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3739),
.B(n_3666),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3716),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3753),
.Y(n_3814)
);

INVx1_ASAP7_75t_SL g3815 ( 
.A(n_3689),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3747),
.B(n_3614),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3796),
.Y(n_3817)
);

OAI31xp33_ASAP7_75t_L g3818 ( 
.A1(n_3775),
.A2(n_3722),
.A3(n_3746),
.B(n_3774),
.Y(n_3818)
);

INVxp67_ASAP7_75t_L g3819 ( 
.A(n_3767),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3778),
.B(n_3734),
.Y(n_3820)
);

AOI321xp33_ASAP7_75t_L g3821 ( 
.A1(n_3777),
.A2(n_3719),
.A3(n_3742),
.B1(n_3741),
.B2(n_3740),
.C(n_3693),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3802),
.Y(n_3822)
);

INVx2_ASAP7_75t_SL g3823 ( 
.A(n_3770),
.Y(n_3823)
);

O2A1O1Ixp33_ASAP7_75t_L g3824 ( 
.A1(n_3768),
.A2(n_3704),
.B(n_3736),
.C(n_3697),
.Y(n_3824)
);

O2A1O1Ixp33_ASAP7_75t_L g3825 ( 
.A1(n_3790),
.A2(n_3698),
.B(n_3695),
.C(n_3707),
.Y(n_3825)
);

OR2x2_ASAP7_75t_L g3826 ( 
.A(n_3765),
.B(n_3737),
.Y(n_3826)
);

OAI21xp33_ASAP7_75t_L g3827 ( 
.A1(n_3763),
.A2(n_3710),
.B(n_3676),
.Y(n_3827)
);

OAI21xp5_ASAP7_75t_SL g3828 ( 
.A1(n_3809),
.A2(n_3718),
.B(n_3717),
.Y(n_3828)
);

OAI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3773),
.A2(n_3744),
.B1(n_3731),
.B2(n_3748),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3764),
.B(n_3699),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3766),
.B(n_3755),
.Y(n_3831)
);

OR2x2_ASAP7_75t_L g3832 ( 
.A(n_3798),
.B(n_3811),
.Y(n_3832)
);

OAI31xp33_ASAP7_75t_L g3833 ( 
.A1(n_3815),
.A2(n_3624),
.A3(n_3587),
.B(n_3743),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3782),
.B(n_3729),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3771),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3776),
.Y(n_3836)
);

NOR2xp67_ASAP7_75t_SL g3837 ( 
.A(n_3784),
.B(n_3649),
.Y(n_3837)
);

O2A1O1Ixp33_ASAP7_75t_L g3838 ( 
.A1(n_3769),
.A2(n_3760),
.B(n_3757),
.C(n_3720),
.Y(n_3838)
);

OAI21xp33_ASAP7_75t_L g3839 ( 
.A1(n_3786),
.A2(n_3732),
.B(n_3761),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3803),
.B(n_3751),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3781),
.B(n_3762),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3812),
.B(n_3612),
.Y(n_3842)
);

OAI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3795),
.A2(n_3626),
.B1(n_3654),
.B2(n_3672),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3816),
.B(n_3613),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3814),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3772),
.Y(n_3846)
);

XNOR2xp5_ASAP7_75t_L g3847 ( 
.A(n_3780),
.B(n_3627),
.Y(n_3847)
);

AOI22xp5_ASAP7_75t_L g3848 ( 
.A1(n_3793),
.A2(n_3615),
.B1(n_3619),
.B2(n_3618),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3794),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3791),
.B(n_3623),
.Y(n_3850)
);

A2O1A1Ixp33_ASAP7_75t_SL g3851 ( 
.A1(n_3810),
.A2(n_3813),
.B(n_3787),
.C(n_3779),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3808),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3807),
.B(n_3629),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_R g3854 ( 
.A1(n_3804),
.A2(n_3553),
.B(n_3633),
.Y(n_3854)
);

AOI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3785),
.A2(n_3634),
.B1(n_3631),
.B2(n_3616),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3800),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3823),
.B(n_3788),
.Y(n_3857)
);

NAND3xp33_ASAP7_75t_L g3858 ( 
.A(n_3818),
.B(n_3792),
.C(n_3789),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3832),
.B(n_3783),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3831),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3819),
.B(n_3799),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3817),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3835),
.B(n_3806),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3837),
.B(n_3805),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3820),
.B(n_3801),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3850),
.B(n_3797),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3849),
.B(n_3637),
.Y(n_3867)
);

INVxp33_ASAP7_75t_L g3868 ( 
.A(n_3847),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3836),
.B(n_3845),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3826),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3841),
.B(n_3647),
.Y(n_3871)
);

INVx1_ASAP7_75t_SL g3872 ( 
.A(n_3830),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3853),
.Y(n_3873)
);

HB1xp67_ASAP7_75t_L g3874 ( 
.A(n_3829),
.Y(n_3874)
);

INVxp67_ASAP7_75t_L g3875 ( 
.A(n_3834),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3822),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3843),
.B(n_3673),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3844),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3827),
.B(n_172),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3828),
.B(n_172),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3842),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3856),
.B(n_173),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3846),
.B(n_174),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3852),
.Y(n_3884)
);

NAND2x1_ASAP7_75t_L g3885 ( 
.A(n_3848),
.B(n_174),
.Y(n_3885)
);

OR2x2_ASAP7_75t_L g3886 ( 
.A(n_3851),
.B(n_176),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3825),
.Y(n_3887)
);

INVxp33_ASAP7_75t_L g3888 ( 
.A(n_3840),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3854),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3821),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3838),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3855),
.B(n_177),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_R g3893 ( 
.A(n_3824),
.B(n_181),
.Y(n_3893)
);

NOR2xp33_ASAP7_75t_L g3894 ( 
.A(n_3839),
.B(n_179),
.Y(n_3894)
);

NAND2x1_ASAP7_75t_L g3895 ( 
.A(n_3833),
.B(n_179),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3823),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3823),
.B(n_181),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3866),
.B(n_182),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3874),
.B(n_182),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3896),
.B(n_183),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3875),
.B(n_184),
.Y(n_3901)
);

HB1xp67_ASAP7_75t_L g3902 ( 
.A(n_3885),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3890),
.B(n_184),
.Y(n_3903)
);

OAI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3858),
.A2(n_1487),
.B(n_1473),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3870),
.B(n_185),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3859),
.Y(n_3906)
);

NOR2xp67_ASAP7_75t_L g3907 ( 
.A(n_3864),
.B(n_185),
.Y(n_3907)
);

NAND2xp33_ASAP7_75t_SL g3908 ( 
.A(n_3893),
.B(n_1496),
.Y(n_3908)
);

NOR2xp33_ASAP7_75t_L g3909 ( 
.A(n_3868),
.B(n_186),
.Y(n_3909)
);

AOI211xp5_ASAP7_75t_L g3910 ( 
.A1(n_3886),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3863),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3887),
.A2(n_1498),
.B1(n_1500),
.B2(n_1497),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3857),
.Y(n_3913)
);

NOR2x1_ASAP7_75t_L g3914 ( 
.A(n_3891),
.B(n_187),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3897),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3892),
.B(n_188),
.Y(n_3916)
);

AOI22xp33_ASAP7_75t_L g3917 ( 
.A1(n_3889),
.A2(n_1728),
.B1(n_1735),
.B2(n_1724),
.Y(n_3917)
);

NOR2xp67_ASAP7_75t_L g3918 ( 
.A(n_3873),
.B(n_189),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3882),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3872),
.B(n_189),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3888),
.B(n_190),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3883),
.Y(n_3922)
);

HB1xp67_ASAP7_75t_L g3923 ( 
.A(n_3895),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3862),
.B(n_191),
.Y(n_3924)
);

INVxp67_ASAP7_75t_L g3925 ( 
.A(n_3894),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3860),
.B(n_191),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3861),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3876),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_3865),
.B(n_3869),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3878),
.B(n_192),
.Y(n_3930)
);

INVx3_ASAP7_75t_L g3931 ( 
.A(n_3884),
.Y(n_3931)
);

XNOR2x1_ASAP7_75t_L g3932 ( 
.A(n_3871),
.B(n_193),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3880),
.B(n_192),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3881),
.B(n_194),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3867),
.B(n_194),
.Y(n_3935)
);

INVxp67_ASAP7_75t_SL g3936 ( 
.A(n_3877),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3879),
.Y(n_3937)
);

AOI211xp5_ASAP7_75t_L g3938 ( 
.A1(n_3890),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3864),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3874),
.B(n_195),
.Y(n_3940)
);

NOR2xp67_ASAP7_75t_SL g3941 ( 
.A(n_3874),
.B(n_1502),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3864),
.Y(n_3942)
);

NOR2x1_ASAP7_75t_L g3943 ( 
.A(n_3886),
.B(n_198),
.Y(n_3943)
);

INVxp67_ASAP7_75t_L g3944 ( 
.A(n_3874),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3866),
.B(n_198),
.Y(n_3945)
);

NOR2xp33_ASAP7_75t_L g3946 ( 
.A(n_3868),
.B(n_199),
.Y(n_3946)
);

NAND3xp33_ASAP7_75t_L g3947 ( 
.A(n_3886),
.B(n_1505),
.C(n_1503),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3944),
.B(n_200),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3923),
.B(n_200),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3906),
.B(n_201),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3907),
.B(n_1511),
.Y(n_3951)
);

NOR3xp33_ASAP7_75t_L g3952 ( 
.A(n_3929),
.B(n_3942),
.C(n_3939),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3918),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_L g3954 ( 
.A(n_3902),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3898),
.B(n_202),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3945),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_3911),
.B(n_203),
.Y(n_3957)
);

OAI21xp33_ASAP7_75t_L g3958 ( 
.A1(n_3903),
.A2(n_1519),
.B(n_1515),
.Y(n_3958)
);

NOR2xp33_ASAP7_75t_L g3959 ( 
.A(n_3919),
.B(n_3922),
.Y(n_3959)
);

NAND2x1_ASAP7_75t_L g3960 ( 
.A(n_3931),
.B(n_205),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3943),
.B(n_206),
.Y(n_3961)
);

AOI211xp5_ASAP7_75t_L g3962 ( 
.A1(n_3899),
.A2(n_209),
.B(n_206),
.C(n_208),
.Y(n_3962)
);

HB1xp67_ASAP7_75t_L g3963 ( 
.A(n_3914),
.Y(n_3963)
);

INVxp67_ASAP7_75t_L g3964 ( 
.A(n_3909),
.Y(n_3964)
);

NOR3xp33_ASAP7_75t_L g3965 ( 
.A(n_3946),
.B(n_1525),
.C(n_1522),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3905),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_SL g3967 ( 
.A(n_3931),
.B(n_1535),
.Y(n_3967)
);

HB1xp67_ASAP7_75t_L g3968 ( 
.A(n_3932),
.Y(n_3968)
);

NOR2xp33_ASAP7_75t_L g3969 ( 
.A(n_3916),
.B(n_209),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3920),
.B(n_210),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3921),
.Y(n_3971)
);

NAND3xp33_ASAP7_75t_L g3972 ( 
.A(n_3938),
.B(n_1558),
.C(n_1546),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3910),
.B(n_211),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3940),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3900),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3908),
.B(n_1560),
.Y(n_3976)
);

OR2x2_ASAP7_75t_L g3977 ( 
.A(n_3901),
.B(n_212),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3933),
.B(n_212),
.Y(n_3978)
);

NOR3xp33_ASAP7_75t_L g3979 ( 
.A(n_3936),
.B(n_1563),
.C(n_1561),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_L g3980 ( 
.A(n_3925),
.B(n_213),
.Y(n_3980)
);

INVxp67_ASAP7_75t_L g3981 ( 
.A(n_3926),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3904),
.A2(n_3935),
.B(n_3924),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3937),
.B(n_215),
.Y(n_3983)
);

NOR3x1_ASAP7_75t_L g3984 ( 
.A(n_3947),
.B(n_216),
.C(n_218),
.Y(n_3984)
);

NOR3xp33_ASAP7_75t_L g3985 ( 
.A(n_3913),
.B(n_1576),
.C(n_1569),
.Y(n_3985)
);

NOR3xp33_ASAP7_75t_L g3986 ( 
.A(n_3927),
.B(n_1591),
.C(n_1579),
.Y(n_3986)
);

NOR3xp33_ASAP7_75t_L g3987 ( 
.A(n_3915),
.B(n_1598),
.C(n_1595),
.Y(n_3987)
);

AOI21xp33_ASAP7_75t_L g3988 ( 
.A1(n_3941),
.A2(n_221),
.B(n_220),
.Y(n_3988)
);

NOR2xp67_ASAP7_75t_L g3989 ( 
.A(n_3928),
.B(n_219),
.Y(n_3989)
);

NOR3xp33_ASAP7_75t_L g3990 ( 
.A(n_3930),
.B(n_1618),
.C(n_1603),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3934),
.B(n_219),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3912),
.Y(n_3992)
);

NOR2xp33_ASAP7_75t_L g3993 ( 
.A(n_3917),
.B(n_220),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3918),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3923),
.B(n_221),
.Y(n_3995)
);

HB1xp67_ASAP7_75t_L g3996 ( 
.A(n_3918),
.Y(n_3996)
);

O2A1O1Ixp33_ASAP7_75t_L g3997 ( 
.A1(n_3944),
.A2(n_230),
.B(n_239),
.C(n_222),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3908),
.A2(n_1631),
.B(n_1622),
.Y(n_3998)
);

AOI321xp33_ASAP7_75t_L g3999 ( 
.A1(n_3936),
.A2(n_224),
.A3(n_226),
.B1(n_222),
.B2(n_223),
.C(n_225),
.Y(n_3999)
);

O2A1O1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_3944),
.A2(n_234),
.B(n_245),
.C(n_223),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3906),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3906),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_L g4003 ( 
.A(n_3923),
.B(n_225),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3923),
.B(n_227),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3906),
.B(n_1634),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3918),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3918),
.Y(n_4007)
);

OAI22x1_ASAP7_75t_L g4008 ( 
.A1(n_3944),
.A2(n_1647),
.B1(n_1659),
.B2(n_1636),
.Y(n_4008)
);

OAI21xp33_ASAP7_75t_SL g4009 ( 
.A1(n_3943),
.A2(n_227),
.B(n_228),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3918),
.Y(n_4010)
);

OAI21xp33_ASAP7_75t_L g4011 ( 
.A1(n_3944),
.A2(n_1662),
.B(n_1661),
.Y(n_4011)
);

AND3x4_ASAP7_75t_L g4012 ( 
.A(n_3943),
.B(n_229),
.C(n_231),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3923),
.B(n_231),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_L g4014 ( 
.A(n_3923),
.B(n_232),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3906),
.Y(n_4015)
);

AOI221xp5_ASAP7_75t_L g4016 ( 
.A1(n_3944),
.A2(n_1674),
.B1(n_1680),
.B2(n_1672),
.C(n_1668),
.Y(n_4016)
);

OR2x2_ASAP7_75t_L g4017 ( 
.A(n_3944),
.B(n_232),
.Y(n_4017)
);

NOR3xp33_ASAP7_75t_L g4018 ( 
.A(n_3906),
.B(n_1693),
.C(n_1687),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3918),
.Y(n_4019)
);

NAND3xp33_ASAP7_75t_L g4020 ( 
.A(n_3923),
.B(n_1707),
.C(n_1705),
.Y(n_4020)
);

XNOR2x2_ASAP7_75t_L g4021 ( 
.A(n_3914),
.B(n_233),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3906),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3908),
.A2(n_1712),
.B(n_1709),
.Y(n_4023)
);

NAND3xp33_ASAP7_75t_SL g4024 ( 
.A(n_3910),
.B(n_1714),
.C(n_1713),
.Y(n_4024)
);

NOR3xp33_ASAP7_75t_L g4025 ( 
.A(n_3906),
.B(n_1744),
.C(n_1738),
.Y(n_4025)
);

NAND4xp75_ASAP7_75t_L g4026 ( 
.A(n_3943),
.B(n_237),
.C(n_233),
.D(n_236),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3906),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3923),
.B(n_236),
.Y(n_4028)
);

AOI21x1_ASAP7_75t_L g4029 ( 
.A1(n_3918),
.A2(n_241),
.B(n_238),
.Y(n_4029)
);

XNOR2xp5_ASAP7_75t_L g4030 ( 
.A(n_3932),
.B(n_238),
.Y(n_4030)
);

AOI222xp33_ASAP7_75t_L g4031 ( 
.A1(n_3954),
.A2(n_242),
.B1(n_244),
.B2(n_237),
.C1(n_241),
.C2(n_243),
.Y(n_4031)
);

NOR3xp33_ASAP7_75t_L g4032 ( 
.A(n_4009),
.B(n_242),
.C(n_243),
.Y(n_4032)
);

OAI221xp5_ASAP7_75t_SL g4033 ( 
.A1(n_4001),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.C(n_248),
.Y(n_4033)
);

NAND2xp33_ASAP7_75t_R g4034 ( 
.A(n_3961),
.B(n_246),
.Y(n_4034)
);

NAND4xp25_ASAP7_75t_SL g4035 ( 
.A(n_3952),
.B(n_252),
.C(n_249),
.D(n_250),
.Y(n_4035)
);

AOI222xp33_ASAP7_75t_L g4036 ( 
.A1(n_3963),
.A2(n_255),
.B1(n_258),
.B2(n_253),
.C1(n_254),
.C2(n_256),
.Y(n_4036)
);

AOI211xp5_ASAP7_75t_L g4037 ( 
.A1(n_4003),
.A2(n_256),
.B(n_253),
.C(n_254),
.Y(n_4037)
);

AOI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_4002),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3951),
.A2(n_259),
.B(n_260),
.Y(n_4039)
);

OAI221xp5_ASAP7_75t_L g4040 ( 
.A1(n_4014),
.A2(n_4022),
.B1(n_4027),
.B2(n_4015),
.C(n_3996),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_4029),
.Y(n_4041)
);

A2O1A1Ixp33_ASAP7_75t_L g4042 ( 
.A1(n_3997),
.A2(n_4000),
.B(n_3989),
.C(n_3999),
.Y(n_4042)
);

INVx1_ASAP7_75t_SL g4043 ( 
.A(n_4021),
.Y(n_4043)
);

A2O1A1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_3959),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_4044)
);

NAND4xp25_ASAP7_75t_L g4045 ( 
.A(n_3956),
.B(n_3966),
.C(n_3982),
.D(n_3964),
.Y(n_4045)
);

AOI221xp5_ASAP7_75t_L g4046 ( 
.A1(n_3953),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_269),
.Y(n_4046)
);

AOI222xp33_ASAP7_75t_L g4047 ( 
.A1(n_3994),
.A2(n_267),
.B1(n_271),
.B2(n_265),
.C1(n_266),
.C2(n_270),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3960),
.Y(n_4048)
);

AOI322xp5_ASAP7_75t_L g4049 ( 
.A1(n_3968),
.A2(n_276),
.A3(n_275),
.B1(n_273),
.B2(n_271),
.C1(n_272),
.C2(n_274),
.Y(n_4049)
);

AND4x2_ASAP7_75t_L g4050 ( 
.A(n_4016),
.B(n_274),
.C(n_272),
.D(n_273),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_4006),
.A2(n_4010),
.B(n_4007),
.Y(n_4051)
);

AOI211xp5_ASAP7_75t_L g4052 ( 
.A1(n_4019),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_4052)
);

NAND4xp75_ASAP7_75t_L g4053 ( 
.A(n_4004),
.B(n_279),
.C(n_277),
.D(n_278),
.Y(n_4053)
);

AOI211xp5_ASAP7_75t_L g4054 ( 
.A1(n_3949),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_4054)
);

AOI22xp5_ASAP7_75t_L g4055 ( 
.A1(n_4012),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3995),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_4013),
.Y(n_4057)
);

AOI21xp33_ASAP7_75t_L g4058 ( 
.A1(n_4028),
.A2(n_283),
.B(n_284),
.Y(n_4058)
);

OAI211xp5_ASAP7_75t_SL g4059 ( 
.A1(n_3981),
.A2(n_288),
.B(n_285),
.C(n_286),
.Y(n_4059)
);

AOI221xp5_ASAP7_75t_L g4060 ( 
.A1(n_4024),
.A2(n_289),
.B1(n_285),
.B2(n_288),
.C(n_291),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3950),
.Y(n_4061)
);

NOR2xp33_ASAP7_75t_L g4062 ( 
.A(n_4026),
.B(n_289),
.Y(n_4062)
);

AOI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3976),
.A2(n_291),
.B(n_292),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_4030),
.B(n_292),
.Y(n_4064)
);

NOR3xp33_ASAP7_75t_L g4065 ( 
.A(n_3974),
.B(n_293),
.C(n_294),
.Y(n_4065)
);

AOI221xp5_ASAP7_75t_L g4066 ( 
.A1(n_4011),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.C(n_297),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3957),
.B(n_295),
.Y(n_4067)
);

AOI211xp5_ASAP7_75t_SL g4068 ( 
.A1(n_3948),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_4068)
);

AOI221xp5_ASAP7_75t_SL g4069 ( 
.A1(n_3971),
.A2(n_303),
.B1(n_298),
.B2(n_302),
.C(n_304),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3969),
.B(n_303),
.Y(n_4070)
);

NOR3xp33_ASAP7_75t_L g4071 ( 
.A(n_3972),
.B(n_305),
.C(n_306),
.Y(n_4071)
);

AOI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_3980),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_4072)
);

AOI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_3967),
.A2(n_307),
.B(n_308),
.Y(n_4073)
);

A2O1A1Ixp33_ASAP7_75t_L g4074 ( 
.A1(n_3993),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_4074)
);

AOI221x1_ASAP7_75t_L g4075 ( 
.A1(n_3979),
.A2(n_312),
.B1(n_309),
.B2(n_310),
.C(n_313),
.Y(n_4075)
);

AOI221xp5_ASAP7_75t_L g4076 ( 
.A1(n_3992),
.A2(n_315),
.B1(n_312),
.B2(n_314),
.C(n_317),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3984),
.B(n_314),
.Y(n_4077)
);

OAI211xp5_ASAP7_75t_SL g4078 ( 
.A1(n_3975),
.A2(n_319),
.B(n_315),
.C(n_318),
.Y(n_4078)
);

INVxp67_ASAP7_75t_SL g4079 ( 
.A(n_3955),
.Y(n_4079)
);

OAI221xp5_ASAP7_75t_SL g4080 ( 
.A1(n_4017),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.C(n_322),
.Y(n_4080)
);

CKINVDCx5p33_ASAP7_75t_R g4081 ( 
.A(n_3970),
.Y(n_4081)
);

OAI211xp5_ASAP7_75t_L g4082 ( 
.A1(n_3958),
.A2(n_329),
.B(n_338),
.C(n_320),
.Y(n_4082)
);

NAND4xp25_ASAP7_75t_L g4083 ( 
.A(n_4020),
.B(n_324),
.C(n_322),
.D(n_323),
.Y(n_4083)
);

NAND4xp25_ASAP7_75t_L g4084 ( 
.A(n_3962),
.B(n_326),
.C(n_323),
.D(n_325),
.Y(n_4084)
);

A2O1A1Ixp33_ASAP7_75t_L g4085 ( 
.A1(n_3988),
.A2(n_328),
.B(n_326),
.C(n_327),
.Y(n_4085)
);

O2A1O1Ixp5_ASAP7_75t_L g4086 ( 
.A1(n_4005),
.A2(n_331),
.B(n_327),
.C(n_330),
.Y(n_4086)
);

NAND4xp25_ASAP7_75t_L g4087 ( 
.A(n_3990),
.B(n_3973),
.C(n_3985),
.D(n_3986),
.Y(n_4087)
);

OAI221xp5_ASAP7_75t_SL g4088 ( 
.A1(n_3983),
.A2(n_334),
.B1(n_330),
.B2(n_333),
.C(n_335),
.Y(n_4088)
);

AOI221xp5_ASAP7_75t_L g4089 ( 
.A1(n_3987),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_4089)
);

AOI221xp5_ASAP7_75t_L g4090 ( 
.A1(n_3965),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.C(n_340),
.Y(n_4090)
);

AOI221xp5_ASAP7_75t_L g4091 ( 
.A1(n_4018),
.A2(n_340),
.B1(n_337),
.B2(n_339),
.C(n_341),
.Y(n_4091)
);

NAND3xp33_ASAP7_75t_L g4092 ( 
.A(n_4025),
.B(n_343),
.C(n_344),
.Y(n_4092)
);

AOI221x1_ASAP7_75t_L g4093 ( 
.A1(n_4008),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.C(n_347),
.Y(n_4093)
);

OAI211xp5_ASAP7_75t_L g4094 ( 
.A1(n_3991),
.A2(n_358),
.B(n_366),
.C(n_345),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3977),
.Y(n_4095)
);

AOI221xp5_ASAP7_75t_L g4096 ( 
.A1(n_3978),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.C(n_352),
.Y(n_4096)
);

O2A1O1Ixp33_ASAP7_75t_SL g4097 ( 
.A1(n_3998),
.A2(n_352),
.B(n_348),
.C(n_349),
.Y(n_4097)
);

AOI222xp33_ASAP7_75t_L g4098 ( 
.A1(n_4023),
.A2(n_356),
.B1(n_359),
.B2(n_354),
.C1(n_355),
.C2(n_358),
.Y(n_4098)
);

OAI22xp5_ASAP7_75t_L g4099 ( 
.A1(n_4001),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_4099)
);

AOI221xp5_ASAP7_75t_SL g4100 ( 
.A1(n_3953),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.C(n_363),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_4029),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4029),
.Y(n_4102)
);

O2A1O1Ixp5_ASAP7_75t_L g4103 ( 
.A1(n_3953),
.A2(n_364),
.B(n_360),
.C(n_363),
.Y(n_4103)
);

INVx4_ASAP7_75t_L g4104 ( 
.A(n_4001),
.Y(n_4104)
);

AOI221xp5_ASAP7_75t_L g4105 ( 
.A1(n_3952),
.A2(n_367),
.B1(n_364),
.B2(n_365),
.C(n_368),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_3954),
.B(n_365),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3954),
.B(n_368),
.Y(n_4107)
);

O2A1O1Ixp5_ASAP7_75t_SL g4108 ( 
.A1(n_3954),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_4108)
);

AOI221xp5_ASAP7_75t_SL g4109 ( 
.A1(n_3953),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_4109)
);

OAI21xp33_ASAP7_75t_L g4110 ( 
.A1(n_3959),
.A2(n_372),
.B(n_374),
.Y(n_4110)
);

AOI22xp33_ASAP7_75t_L g4111 ( 
.A1(n_4001),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4111)
);

OAI221xp5_ASAP7_75t_L g4112 ( 
.A1(n_4009),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.C(n_380),
.Y(n_4112)
);

NOR3xp33_ASAP7_75t_L g4113 ( 
.A(n_4009),
.B(n_379),
.C(n_381),
.Y(n_4113)
);

XNOR2xp5_ASAP7_75t_L g4114 ( 
.A(n_4055),
.B(n_381),
.Y(n_4114)
);

OAI21xp5_ASAP7_75t_L g4115 ( 
.A1(n_4051),
.A2(n_384),
.B(n_383),
.Y(n_4115)
);

AOI222xp33_ASAP7_75t_L g4116 ( 
.A1(n_4043),
.A2(n_384),
.B1(n_386),
.B2(n_382),
.C1(n_383),
.C2(n_385),
.Y(n_4116)
);

AOI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_4032),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_4117)
);

OAI211xp5_ASAP7_75t_SL g4118 ( 
.A1(n_4040),
.A2(n_4042),
.B(n_4061),
.C(n_4057),
.Y(n_4118)
);

NAND4xp25_ASAP7_75t_L g4119 ( 
.A(n_4045),
.B(n_389),
.C(n_387),
.D(n_388),
.Y(n_4119)
);

NAND4xp25_ASAP7_75t_L g4120 ( 
.A(n_4113),
.B(n_392),
.C(n_389),
.D(n_390),
.Y(n_4120)
);

INVx1_ASAP7_75t_SL g4121 ( 
.A(n_4048),
.Y(n_4121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g4122 ( 
.A1(n_4041),
.A2(n_394),
.B(n_392),
.C(n_393),
.D(n_396),
.Y(n_4122)
);

AOI221xp5_ASAP7_75t_L g4123 ( 
.A1(n_4101),
.A2(n_398),
.B1(n_394),
.B2(n_397),
.C(n_399),
.Y(n_4123)
);

AOI221xp5_ASAP7_75t_L g4124 ( 
.A1(n_4102),
.A2(n_401),
.B1(n_398),
.B2(n_399),
.C(n_402),
.Y(n_4124)
);

AOI221xp5_ASAP7_75t_L g4125 ( 
.A1(n_4104),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.C(n_406),
.Y(n_4125)
);

OAI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_4103),
.A2(n_4086),
.B(n_4106),
.Y(n_4126)
);

NAND4xp25_ASAP7_75t_L g4127 ( 
.A(n_4104),
.B(n_4095),
.C(n_4087),
.D(n_4034),
.Y(n_4127)
);

AOI221xp5_ASAP7_75t_L g4128 ( 
.A1(n_4112),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.C(n_407),
.Y(n_4128)
);

AOI211xp5_ASAP7_75t_L g4129 ( 
.A1(n_4035),
.A2(n_411),
.B(n_407),
.C(n_408),
.Y(n_4129)
);

AOI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_4062),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4130)
);

AOI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_4056),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4131)
);

OAI21x1_ASAP7_75t_SL g4132 ( 
.A1(n_4039),
.A2(n_415),
.B(n_416),
.Y(n_4132)
);

A2O1A1Ixp33_ASAP7_75t_SL g4133 ( 
.A1(n_4079),
.A2(n_4107),
.B(n_4068),
.C(n_4065),
.Y(n_4133)
);

OA22x2_ASAP7_75t_SL g4134 ( 
.A1(n_4050),
.A2(n_420),
.B1(n_421),
.B2(n_418),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_4077),
.Y(n_4135)
);

OAI321xp33_ASAP7_75t_L g4136 ( 
.A1(n_4084),
.A2(n_422),
.A3(n_425),
.B1(n_417),
.B2(n_421),
.C(n_424),
.Y(n_4136)
);

OAI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_4108),
.A2(n_425),
.B(n_422),
.Y(n_4137)
);

AND4x1_ASAP7_75t_L g4138 ( 
.A(n_4052),
.B(n_4054),
.C(n_4037),
.D(n_4031),
.Y(n_4138)
);

INVx1_ASAP7_75t_SL g4139 ( 
.A(n_4053),
.Y(n_4139)
);

OAI211xp5_ASAP7_75t_L g4140 ( 
.A1(n_4093),
.A2(n_427),
.B(n_417),
.C(n_426),
.Y(n_4140)
);

AOI22xp5_ASAP7_75t_L g4141 ( 
.A1(n_4081),
.A2(n_429),
.B1(n_426),
.B2(n_428),
.Y(n_4141)
);

NOR3xp33_ASAP7_75t_L g4142 ( 
.A(n_4092),
.B(n_430),
.C(n_429),
.Y(n_4142)
);

NAND3xp33_ASAP7_75t_SL g4143 ( 
.A(n_4071),
.B(n_428),
.C(n_431),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4064),
.Y(n_4144)
);

OAI211xp5_ASAP7_75t_L g4145 ( 
.A1(n_4036),
.A2(n_434),
.B(n_431),
.C(n_432),
.Y(n_4145)
);

OAI221xp5_ASAP7_75t_L g4146 ( 
.A1(n_4100),
.A2(n_4109),
.B1(n_4069),
.B2(n_4110),
.C(n_4085),
.Y(n_4146)
);

NOR3xp33_ASAP7_75t_L g4147 ( 
.A(n_4070),
.B(n_436),
.C(n_435),
.Y(n_4147)
);

AND4x1_ASAP7_75t_L g4148 ( 
.A(n_4075),
.B(n_438),
.C(n_432),
.D(n_436),
.Y(n_4148)
);

AOI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_4059),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_4097),
.A2(n_440),
.B(n_441),
.Y(n_4150)
);

AOI311xp33_ASAP7_75t_L g4151 ( 
.A1(n_4058),
.A2(n_4063),
.A3(n_4073),
.B(n_4094),
.C(n_4082),
.Y(n_4151)
);

OAI211xp5_ASAP7_75t_SL g4152 ( 
.A1(n_4060),
.A2(n_445),
.B(n_442),
.C(n_443),
.Y(n_4152)
);

NAND4xp75_ASAP7_75t_L g4153 ( 
.A(n_4105),
.B(n_448),
.C(n_442),
.D(n_447),
.Y(n_4153)
);

HB1xp67_ASAP7_75t_L g4154 ( 
.A(n_4099),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4047),
.B(n_447),
.Y(n_4155)
);

BUFx2_ASAP7_75t_L g4156 ( 
.A(n_4044),
.Y(n_4156)
);

O2A1O1Ixp33_ASAP7_75t_L g4157 ( 
.A1(n_4078),
.A2(n_450),
.B(n_448),
.C(n_449),
.Y(n_4157)
);

AOI211xp5_ASAP7_75t_L g4158 ( 
.A1(n_4080),
.A2(n_452),
.B(n_449),
.C(n_451),
.Y(n_4158)
);

AOI22xp33_ASAP7_75t_L g4159 ( 
.A1(n_4083),
.A2(n_455),
.B1(n_451),
.B2(n_454),
.Y(n_4159)
);

AOI211x1_ASAP7_75t_SL g4160 ( 
.A1(n_4074),
.A2(n_457),
.B(n_454),
.C(n_456),
.Y(n_4160)
);

INVxp67_ASAP7_75t_L g4161 ( 
.A(n_4067),
.Y(n_4161)
);

NOR4xp75_ASAP7_75t_SL g4162 ( 
.A(n_4088),
.B(n_466),
.C(n_474),
.D(n_458),
.Y(n_4162)
);

AOI221xp5_ASAP7_75t_L g4163 ( 
.A1(n_4033),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.C(n_461),
.Y(n_4163)
);

OAI221xp5_ASAP7_75t_L g4164 ( 
.A1(n_4046),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.C(n_463),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4072),
.Y(n_4165)
);

AOI21xp5_ASAP7_75t_L g4166 ( 
.A1(n_4096),
.A2(n_4066),
.B(n_4089),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_SL g4167 ( 
.A(n_4098),
.B(n_4076),
.Y(n_4167)
);

OAI211xp5_ASAP7_75t_L g4168 ( 
.A1(n_4111),
.A2(n_465),
.B(n_462),
.C(n_464),
.Y(n_4168)
);

OAI211xp5_ASAP7_75t_L g4169 ( 
.A1(n_4091),
.A2(n_468),
.B(n_465),
.C(n_467),
.Y(n_4169)
);

OAI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_4038),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_4170)
);

XOR2xp5_ASAP7_75t_L g4171 ( 
.A(n_4049),
.B(n_470),
.Y(n_4171)
);

AOI221xp5_ASAP7_75t_L g4172 ( 
.A1(n_4090),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.C(n_473),
.Y(n_4172)
);

OAI211xp5_ASAP7_75t_SL g4173 ( 
.A1(n_4040),
.A2(n_474),
.B(n_471),
.C(n_472),
.Y(n_4173)
);

OAI21xp5_ASAP7_75t_SL g4174 ( 
.A1(n_4043),
.A2(n_475),
.B(n_476),
.Y(n_4174)
);

OAI221xp5_ASAP7_75t_SL g4175 ( 
.A1(n_4043),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.C(n_479),
.Y(n_4175)
);

AOI21xp33_ASAP7_75t_L g4176 ( 
.A1(n_4034),
.A2(n_477),
.B(n_478),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4041),
.Y(n_4177)
);

NOR2xp33_ASAP7_75t_L g4178 ( 
.A(n_4043),
.B(n_480),
.Y(n_4178)
);

INVxp67_ASAP7_75t_SL g4179 ( 
.A(n_4048),
.Y(n_4179)
);

AOI22xp33_ASAP7_75t_L g4180 ( 
.A1(n_4043),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_4180)
);

AOI211xp5_ASAP7_75t_L g4181 ( 
.A1(n_4040),
.A2(n_486),
.B(n_482),
.C(n_485),
.Y(n_4181)
);

NAND4xp25_ASAP7_75t_L g4182 ( 
.A(n_4042),
.B(n_487),
.C(n_485),
.D(n_486),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4043),
.B(n_487),
.Y(n_4183)
);

OAI211xp5_ASAP7_75t_L g4184 ( 
.A1(n_4051),
.A2(n_490),
.B(n_488),
.C(n_489),
.Y(n_4184)
);

AOI211xp5_ASAP7_75t_L g4185 ( 
.A1(n_4040),
.A2(n_491),
.B(n_488),
.C(n_490),
.Y(n_4185)
);

BUFx6f_ASAP7_75t_L g4186 ( 
.A(n_4104),
.Y(n_4186)
);

AOI22xp5_ASAP7_75t_L g4187 ( 
.A1(n_4043),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_4187)
);

OAI21xp5_ASAP7_75t_L g4188 ( 
.A1(n_4051),
.A2(n_495),
.B(n_494),
.Y(n_4188)
);

BUFx2_ASAP7_75t_L g4189 ( 
.A(n_4048),
.Y(n_4189)
);

O2A1O1Ixp33_ASAP7_75t_L g4190 ( 
.A1(n_4043),
.A2(n_495),
.B(n_493),
.C(n_494),
.Y(n_4190)
);

HB1xp67_ASAP7_75t_L g4191 ( 
.A(n_4048),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4043),
.B(n_496),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4041),
.Y(n_4193)
);

NAND4xp25_ASAP7_75t_SL g4194 ( 
.A(n_4043),
.B(n_499),
.C(n_497),
.D(n_498),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4043),
.B(n_497),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4041),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4041),
.Y(n_4197)
);

AOI211xp5_ASAP7_75t_L g4198 ( 
.A1(n_4040),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_4198)
);

AOI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_4121),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_4199)
);

NOR4xp75_ASAP7_75t_L g4200 ( 
.A(n_4126),
.B(n_505),
.C(n_502),
.D(n_504),
.Y(n_4200)
);

OAI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_4180),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_SL g4202 ( 
.A(n_4162),
.B(n_2078),
.Y(n_4202)
);

AOI22xp33_ASAP7_75t_L g4203 ( 
.A1(n_4189),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_4203)
);

AOI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_4133),
.A2(n_508),
.B(n_509),
.Y(n_4204)
);

OAI211xp5_ASAP7_75t_L g4205 ( 
.A1(n_4174),
.A2(n_513),
.B(n_509),
.C(n_512),
.Y(n_4205)
);

NAND3x1_ASAP7_75t_L g4206 ( 
.A(n_4122),
.B(n_512),
.C(n_513),
.Y(n_4206)
);

OAI211xp5_ASAP7_75t_SL g4207 ( 
.A1(n_4167),
.A2(n_516),
.B(n_514),
.C(n_515),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4186),
.Y(n_4208)
);

NOR3xp33_ASAP7_75t_L g4209 ( 
.A(n_4118),
.B(n_515),
.C(n_517),
.Y(n_4209)
);

INVx1_ASAP7_75t_SL g4210 ( 
.A(n_4183),
.Y(n_4210)
);

AOI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_4139),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_4211)
);

AOI221xp5_ASAP7_75t_L g4212 ( 
.A1(n_4190),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.C(n_521),
.Y(n_4212)
);

AND3x1_ASAP7_75t_L g4213 ( 
.A(n_4129),
.B(n_521),
.C(n_522),
.Y(n_4213)
);

O2A1O1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_4173),
.A2(n_524),
.B(n_522),
.C(n_523),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4135),
.B(n_523),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4179),
.B(n_524),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4191),
.B(n_525),
.Y(n_4217)
);

XNOR2x1_ASAP7_75t_L g4218 ( 
.A(n_4114),
.B(n_526),
.Y(n_4218)
);

OAI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_4187),
.A2(n_528),
.B1(n_526),
.B2(n_527),
.Y(n_4219)
);

A2O1A1Ixp33_ASAP7_75t_L g4220 ( 
.A1(n_4178),
.A2(n_529),
.B(n_527),
.C(n_528),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_L g4221 ( 
.A(n_4182),
.B(n_4175),
.Y(n_4221)
);

OAI221xp5_ASAP7_75t_L g4222 ( 
.A1(n_4181),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.C(n_532),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4116),
.B(n_530),
.Y(n_4223)
);

NOR2xp67_ASAP7_75t_L g4224 ( 
.A(n_4194),
.B(n_531),
.Y(n_4224)
);

AOI322xp5_ASAP7_75t_L g4225 ( 
.A1(n_4192),
.A2(n_539),
.A3(n_538),
.B1(n_536),
.B2(n_533),
.C1(n_534),
.C2(n_537),
.Y(n_4225)
);

OAI211xp5_ASAP7_75t_L g4226 ( 
.A1(n_4140),
.A2(n_536),
.B(n_533),
.C(n_534),
.Y(n_4226)
);

NOR2x1_ASAP7_75t_L g4227 ( 
.A(n_4119),
.B(n_538),
.Y(n_4227)
);

INVx2_ASAP7_75t_SL g4228 ( 
.A(n_4186),
.Y(n_4228)
);

NOR2x1_ASAP7_75t_L g4229 ( 
.A(n_4127),
.B(n_540),
.Y(n_4229)
);

OAI22xp5_ASAP7_75t_L g4230 ( 
.A1(n_4149),
.A2(n_4159),
.B1(n_4130),
.B2(n_4117),
.Y(n_4230)
);

AOI22xp33_ASAP7_75t_L g4231 ( 
.A1(n_4156),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_4231)
);

AOI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_4171),
.A2(n_545),
.B1(n_542),
.B2(n_543),
.Y(n_4232)
);

AOI321xp33_ASAP7_75t_L g4233 ( 
.A1(n_4151),
.A2(n_549),
.A3(n_551),
.B1(n_543),
.B2(n_546),
.C(n_550),
.Y(n_4233)
);

NOR3xp33_ASAP7_75t_L g4234 ( 
.A(n_4120),
.B(n_549),
.C(n_550),
.Y(n_4234)
);

NOR3xp33_ASAP7_75t_SL g4235 ( 
.A(n_4143),
.B(n_551),
.C(n_552),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_4154),
.B(n_552),
.Y(n_4236)
);

INVx1_ASAP7_75t_SL g4237 ( 
.A(n_4195),
.Y(n_4237)
);

OR2x2_ASAP7_75t_L g4238 ( 
.A(n_4155),
.B(n_553),
.Y(n_4238)
);

NAND3x1_ASAP7_75t_L g4239 ( 
.A(n_4148),
.B(n_554),
.C(n_555),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4177),
.B(n_554),
.Y(n_4240)
);

A2O1A1Ixp33_ASAP7_75t_L g4241 ( 
.A1(n_4157),
.A2(n_557),
.B(n_555),
.C(n_556),
.Y(n_4241)
);

OAI221xp5_ASAP7_75t_L g4242 ( 
.A1(n_4185),
.A2(n_4198),
.B1(n_4134),
.B2(n_4158),
.C(n_4188),
.Y(n_4242)
);

O2A1O1Ixp33_ASAP7_75t_L g4243 ( 
.A1(n_4176),
.A2(n_559),
.B(n_556),
.C(n_557),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_4165),
.A2(n_562),
.B1(n_559),
.B2(n_561),
.Y(n_4244)
);

NOR2x1_ASAP7_75t_L g4245 ( 
.A(n_4184),
.B(n_4137),
.Y(n_4245)
);

O2A1O1Ixp33_ASAP7_75t_L g4246 ( 
.A1(n_4193),
.A2(n_4197),
.B(n_4196),
.C(n_4132),
.Y(n_4246)
);

NOR2x1_ASAP7_75t_L g4247 ( 
.A(n_4186),
.B(n_562),
.Y(n_4247)
);

NAND2x1p5_ASAP7_75t_L g4248 ( 
.A(n_4138),
.B(n_564),
.Y(n_4248)
);

AOI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_4150),
.A2(n_563),
.B(n_564),
.Y(n_4249)
);

AOI221xp5_ASAP7_75t_L g4250 ( 
.A1(n_4146),
.A2(n_569),
.B1(n_563),
.B2(n_566),
.C(n_570),
.Y(n_4250)
);

XNOR2xp5_ASAP7_75t_L g4251 ( 
.A(n_4153),
.B(n_566),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_4136),
.B(n_571),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4160),
.B(n_4163),
.Y(n_4253)
);

AOI221x1_ASAP7_75t_L g4254 ( 
.A1(n_4147),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.C(n_574),
.Y(n_4254)
);

OAI211xp5_ASAP7_75t_SL g4255 ( 
.A1(n_4166),
.A2(n_575),
.B(n_572),
.C(n_574),
.Y(n_4255)
);

NOR2xp33_ASAP7_75t_L g4256 ( 
.A(n_4145),
.B(n_575),
.Y(n_4256)
);

HB1xp67_ASAP7_75t_L g4257 ( 
.A(n_4115),
.Y(n_4257)
);

XOR2xp5_ASAP7_75t_L g4258 ( 
.A(n_4141),
.B(n_576),
.Y(n_4258)
);

AOI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_4142),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_4144),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.Y(n_4260)
);

AOI211xp5_ASAP7_75t_L g4261 ( 
.A1(n_4169),
.A2(n_583),
.B(n_581),
.C(n_582),
.Y(n_4261)
);

NAND4xp75_ASAP7_75t_L g4262 ( 
.A(n_4123),
.B(n_585),
.C(n_583),
.D(n_584),
.Y(n_4262)
);

AOI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_4164),
.A2(n_584),
.B(n_586),
.Y(n_4263)
);

NAND3xp33_ASAP7_75t_SL g4264 ( 
.A(n_4168),
.B(n_588),
.C(n_591),
.Y(n_4264)
);

NOR3xp33_ASAP7_75t_L g4265 ( 
.A(n_4128),
.B(n_588),
.C(n_592),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4124),
.B(n_592),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4161),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4131),
.B(n_4125),
.Y(n_4268)
);

OAI22xp33_ASAP7_75t_L g4269 ( 
.A1(n_4170),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.Y(n_4269)
);

AND2x4_ASAP7_75t_L g4270 ( 
.A(n_4152),
.B(n_594),
.Y(n_4270)
);

OAI211xp5_ASAP7_75t_L g4271 ( 
.A1(n_4172),
.A2(n_598),
.B(n_596),
.C(n_597),
.Y(n_4271)
);

AOI221xp5_ASAP7_75t_SL g4272 ( 
.A1(n_4121),
.A2(n_599),
.B1(n_596),
.B2(n_598),
.C(n_600),
.Y(n_4272)
);

INVx2_ASAP7_75t_SL g4273 ( 
.A(n_4186),
.Y(n_4273)
);

OAI221xp5_ASAP7_75t_L g4274 ( 
.A1(n_4174),
.A2(n_602),
.B1(n_599),
.B2(n_601),
.C(n_603),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4247),
.Y(n_4275)
);

NOR2xp67_ASAP7_75t_L g4276 ( 
.A(n_4226),
.B(n_604),
.Y(n_4276)
);

OAI22xp5_ASAP7_75t_L g4277 ( 
.A1(n_4232),
.A2(n_606),
.B1(n_602),
.B2(n_604),
.Y(n_4277)
);

NAND4xp75_ASAP7_75t_L g4278 ( 
.A(n_4229),
.B(n_4204),
.C(n_4217),
.D(n_4236),
.Y(n_4278)
);

NOR3xp33_ASAP7_75t_L g4279 ( 
.A(n_4228),
.B(n_615),
.C(n_606),
.Y(n_4279)
);

NAND3xp33_ASAP7_75t_SL g4280 ( 
.A(n_4209),
.B(n_608),
.C(n_609),
.Y(n_4280)
);

OAI31xp33_ASAP7_75t_L g4281 ( 
.A1(n_4205),
.A2(n_611),
.A3(n_608),
.B(n_610),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4248),
.B(n_610),
.Y(n_4282)
);

INVxp33_ASAP7_75t_SL g4283 ( 
.A(n_4251),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4215),
.Y(n_4284)
);

NAND5xp2_ASAP7_75t_L g4285 ( 
.A(n_4221),
.B(n_614),
.C(n_612),
.D(n_613),
.E(n_615),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4239),
.Y(n_4286)
);

NAND3xp33_ASAP7_75t_SL g4287 ( 
.A(n_4233),
.B(n_612),
.C(n_613),
.Y(n_4287)
);

AOI31xp33_ASAP7_75t_L g4288 ( 
.A1(n_4272),
.A2(n_4261),
.A3(n_4252),
.B(n_4245),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_SL g4289 ( 
.A(n_4224),
.B(n_614),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_4213),
.Y(n_4290)
);

NOR4xp75_ASAP7_75t_SL g4291 ( 
.A(n_4206),
.B(n_618),
.C(n_616),
.D(n_617),
.Y(n_4291)
);

NOR2x1_ASAP7_75t_L g4292 ( 
.A(n_4202),
.B(n_616),
.Y(n_4292)
);

NAND3xp33_ASAP7_75t_L g4293 ( 
.A(n_4254),
.B(n_618),
.C(n_619),
.Y(n_4293)
);

INVxp67_ASAP7_75t_SL g4294 ( 
.A(n_4214),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4216),
.Y(n_4295)
);

AO211x2_ASAP7_75t_L g4296 ( 
.A1(n_4265),
.A2(n_4249),
.B(n_4234),
.C(n_4208),
.Y(n_4296)
);

OR2x2_ASAP7_75t_L g4297 ( 
.A(n_4223),
.B(n_619),
.Y(n_4297)
);

AOI311xp33_ASAP7_75t_L g4298 ( 
.A1(n_4242),
.A2(n_625),
.A3(n_622),
.B(n_623),
.C(n_626),
.Y(n_4298)
);

NOR2x1_ASAP7_75t_L g4299 ( 
.A(n_4220),
.B(n_626),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4211),
.A2(n_4259),
.B1(n_4222),
.B2(n_4274),
.Y(n_4300)
);

NAND4xp25_ASAP7_75t_L g4301 ( 
.A(n_4253),
.B(n_629),
.C(n_627),
.D(n_628),
.Y(n_4301)
);

INVx1_ASAP7_75t_SL g4302 ( 
.A(n_4200),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4273),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4238),
.Y(n_4304)
);

NAND4xp75_ASAP7_75t_L g4305 ( 
.A(n_4227),
.B(n_630),
.C(n_627),
.D(n_629),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4240),
.Y(n_4306)
);

NAND3xp33_ASAP7_75t_SL g4307 ( 
.A(n_4212),
.B(n_630),
.C(n_631),
.Y(n_4307)
);

AOI21x1_ASAP7_75t_L g4308 ( 
.A1(n_4218),
.A2(n_632),
.B(n_633),
.Y(n_4308)
);

NAND4xp75_ASAP7_75t_L g4309 ( 
.A(n_4256),
.B(n_635),
.C(n_632),
.D(n_634),
.Y(n_4309)
);

AOI21xp33_ASAP7_75t_SL g4310 ( 
.A1(n_4219),
.A2(n_634),
.B(n_636),
.Y(n_4310)
);

NOR3xp33_ASAP7_75t_SL g4311 ( 
.A(n_4264),
.B(n_636),
.C(n_637),
.Y(n_4311)
);

NOR2x1p5_ASAP7_75t_L g4312 ( 
.A(n_4262),
.B(n_637),
.Y(n_4312)
);

AOI32xp33_ASAP7_75t_L g4313 ( 
.A1(n_4270),
.A2(n_641),
.A3(n_638),
.B1(n_639),
.B2(n_642),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4270),
.Y(n_4314)
);

AND3x4_ASAP7_75t_L g4315 ( 
.A(n_4235),
.B(n_639),
.C(n_641),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_4257),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4231),
.B(n_642),
.Y(n_4317)
);

OAI211xp5_ASAP7_75t_L g4318 ( 
.A1(n_4271),
.A2(n_645),
.B(n_643),
.C(n_644),
.Y(n_4318)
);

NAND3x1_ASAP7_75t_L g4319 ( 
.A(n_4266),
.B(n_644),
.C(n_645),
.Y(n_4319)
);

NAND5xp2_ASAP7_75t_L g4320 ( 
.A(n_4246),
.B(n_648),
.C(n_646),
.D(n_647),
.E(n_649),
.Y(n_4320)
);

HB1xp67_ASAP7_75t_L g4321 ( 
.A(n_4201),
.Y(n_4321)
);

OR2x2_ASAP7_75t_L g4322 ( 
.A(n_4210),
.B(n_646),
.Y(n_4322)
);

OR2x2_ASAP7_75t_L g4323 ( 
.A(n_4237),
.B(n_648),
.Y(n_4323)
);

AND2x4_ASAP7_75t_L g4324 ( 
.A(n_4267),
.B(n_649),
.Y(n_4324)
);

NOR3xp33_ASAP7_75t_L g4325 ( 
.A(n_4243),
.B(n_650),
.C(n_651),
.Y(n_4325)
);

NOR2xp67_ASAP7_75t_L g4326 ( 
.A(n_4199),
.B(n_650),
.Y(n_4326)
);

AND2x4_ASAP7_75t_L g4327 ( 
.A(n_4241),
.B(n_651),
.Y(n_4327)
);

OR2x2_ASAP7_75t_L g4328 ( 
.A(n_4268),
.B(n_652),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4258),
.Y(n_4329)
);

CKINVDCx5p33_ASAP7_75t_R g4330 ( 
.A(n_4283),
.Y(n_4330)
);

CKINVDCx5p33_ASAP7_75t_R g4331 ( 
.A(n_4316),
.Y(n_4331)
);

CKINVDCx5p33_ASAP7_75t_R g4332 ( 
.A(n_4303),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4324),
.Y(n_4333)
);

HB1xp67_ASAP7_75t_L g4334 ( 
.A(n_4275),
.Y(n_4334)
);

INVx1_ASAP7_75t_SL g4335 ( 
.A(n_4282),
.Y(n_4335)
);

CKINVDCx16_ASAP7_75t_R g4336 ( 
.A(n_4287),
.Y(n_4336)
);

CKINVDCx16_ASAP7_75t_R g4337 ( 
.A(n_4290),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4324),
.Y(n_4338)
);

AOI31xp33_ASAP7_75t_L g4339 ( 
.A1(n_4289),
.A2(n_4250),
.A3(n_4263),
.B(n_4230),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4308),
.Y(n_4340)
);

INVx1_ASAP7_75t_SL g4341 ( 
.A(n_4302),
.Y(n_4341)
);

HB1xp67_ASAP7_75t_L g4342 ( 
.A(n_4305),
.Y(n_4342)
);

AND4x1_ASAP7_75t_L g4343 ( 
.A(n_4298),
.B(n_4203),
.C(n_4244),
.D(n_4260),
.Y(n_4343)
);

INVx3_ASAP7_75t_SL g4344 ( 
.A(n_4322),
.Y(n_4344)
);

AOI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_4315),
.A2(n_4207),
.B1(n_4255),
.B2(n_4269),
.Y(n_4345)
);

HB1xp67_ASAP7_75t_L g4346 ( 
.A(n_4276),
.Y(n_4346)
);

CKINVDCx5p33_ASAP7_75t_R g4347 ( 
.A(n_4284),
.Y(n_4347)
);

HB1xp67_ASAP7_75t_L g4348 ( 
.A(n_4312),
.Y(n_4348)
);

CKINVDCx5p33_ASAP7_75t_R g4349 ( 
.A(n_4286),
.Y(n_4349)
);

INVx2_ASAP7_75t_SL g4350 ( 
.A(n_4323),
.Y(n_4350)
);

BUFx2_ASAP7_75t_L g4351 ( 
.A(n_4314),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4313),
.B(n_4225),
.Y(n_4352)
);

AND2x4_ASAP7_75t_L g4353 ( 
.A(n_4292),
.B(n_653),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4293),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_R g4355 ( 
.A(n_4280),
.B(n_654),
.Y(n_4355)
);

HB1xp67_ASAP7_75t_L g4356 ( 
.A(n_4278),
.Y(n_4356)
);

NAND4xp25_ASAP7_75t_L g4357 ( 
.A(n_4281),
.B(n_657),
.C(n_655),
.D(n_656),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4311),
.B(n_656),
.Y(n_4358)
);

CKINVDCx5p33_ASAP7_75t_R g4359 ( 
.A(n_4328),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4309),
.Y(n_4360)
);

BUFx2_ASAP7_75t_L g4361 ( 
.A(n_4299),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4317),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_4297),
.Y(n_4363)
);

XNOR2x1_ASAP7_75t_SL g4364 ( 
.A(n_4350),
.B(n_4329),
.Y(n_4364)
);

OAI22xp5_ASAP7_75t_SL g4365 ( 
.A1(n_4337),
.A2(n_4294),
.B1(n_4321),
.B2(n_4327),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4351),
.Y(n_4366)
);

AOI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_4341),
.A2(n_4288),
.B(n_4320),
.Y(n_4367)
);

NAND3xp33_ASAP7_75t_L g4368 ( 
.A(n_4331),
.B(n_4325),
.C(n_4279),
.Y(n_4368)
);

AND3x1_ASAP7_75t_L g4369 ( 
.A(n_4358),
.B(n_4285),
.C(n_4304),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4334),
.Y(n_4370)
);

OAI211xp5_ASAP7_75t_SL g4371 ( 
.A1(n_4352),
.A2(n_4295),
.B(n_4306),
.C(n_4300),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4332),
.A2(n_4349),
.B1(n_4330),
.B2(n_4336),
.Y(n_4372)
);

AOI22x1_ASAP7_75t_L g4373 ( 
.A1(n_4361),
.A2(n_4327),
.B1(n_4291),
.B2(n_4296),
.Y(n_4373)
);

NOR3xp33_ASAP7_75t_L g4374 ( 
.A(n_4356),
.B(n_4307),
.C(n_4318),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4333),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4353),
.B(n_4326),
.Y(n_4376)
);

CKINVDCx20_ASAP7_75t_R g4377 ( 
.A(n_4347),
.Y(n_4377)
);

XNOR2xp5_ASAP7_75t_L g4378 ( 
.A(n_4343),
.B(n_4319),
.Y(n_4378)
);

AOI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_4360),
.A2(n_4277),
.B1(n_4301),
.B2(n_4310),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4345),
.A2(n_660),
.B1(n_657),
.B2(n_658),
.Y(n_4380)
);

NOR3xp33_ASAP7_75t_L g4381 ( 
.A(n_4371),
.B(n_4338),
.C(n_4346),
.Y(n_4381)
);

HB1xp67_ASAP7_75t_L g4382 ( 
.A(n_4366),
.Y(n_4382)
);

XNOR2xp5_ASAP7_75t_L g4383 ( 
.A(n_4369),
.B(n_4342),
.Y(n_4383)
);

OAI21x1_ASAP7_75t_SL g4384 ( 
.A1(n_4373),
.A2(n_4354),
.B(n_4340),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4378),
.Y(n_4385)
);

INVx2_ASAP7_75t_SL g4386 ( 
.A(n_4375),
.Y(n_4386)
);

OAI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4372),
.A2(n_4339),
.B1(n_4357),
.B2(n_4344),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4370),
.B(n_4353),
.Y(n_4388)
);

OAI22x1_ASAP7_75t_L g4389 ( 
.A1(n_4379),
.A2(n_4335),
.B1(n_4348),
.B2(n_4359),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4365),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4376),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4382),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4386),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4388),
.Y(n_4394)
);

INVxp67_ASAP7_75t_SL g4395 ( 
.A(n_4383),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4384),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4385),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4390),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4392),
.Y(n_4399)
);

OAI22xp5_ASAP7_75t_SL g4400 ( 
.A1(n_4396),
.A2(n_4377),
.B1(n_4395),
.B2(n_4368),
.Y(n_4400)
);

OAI22xp5_ASAP7_75t_L g4401 ( 
.A1(n_4397),
.A2(n_4391),
.B1(n_4367),
.B2(n_4363),
.Y(n_4401)
);

OAI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4398),
.A2(n_4393),
.B1(n_4394),
.B2(n_4362),
.Y(n_4402)
);

INVx1_ASAP7_75t_SL g4403 ( 
.A(n_4392),
.Y(n_4403)
);

A2O1A1Ixp33_ASAP7_75t_L g4404 ( 
.A1(n_4399),
.A2(n_4381),
.B(n_4374),
.C(n_4380),
.Y(n_4404)
);

OA21x2_ASAP7_75t_L g4405 ( 
.A1(n_4403),
.A2(n_4364),
.B(n_4389),
.Y(n_4405)
);

OAI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4404),
.A2(n_4400),
.B1(n_4401),
.B2(n_4402),
.Y(n_4406)
);

AOI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_4406),
.A2(n_4405),
.B1(n_4387),
.B2(n_4355),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4407),
.B(n_658),
.Y(n_4408)
);

AOI21xp33_ASAP7_75t_L g4409 ( 
.A1(n_4408),
.A2(n_660),
.B(n_661),
.Y(n_4409)
);

OAI22xp5_ASAP7_75t_SL g4410 ( 
.A1(n_4409),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.Y(n_4410)
);

AOI211xp5_ASAP7_75t_L g4411 ( 
.A1(n_4410),
.A2(n_665),
.B(n_662),
.C(n_664),
.Y(n_4411)
);


endmodule