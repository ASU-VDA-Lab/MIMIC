module fake_jpeg_21437_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_21),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_38),
.B1(n_41),
.B2(n_36),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_11),
.B1(n_29),
.B2(n_27),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_4),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_64),
.B1(n_4),
.B2(n_6),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_85),
.A2(n_78),
.B(n_74),
.C(n_81),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_80),
.A3(n_86),
.B1(n_84),
.B2(n_82),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_31),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_12),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_14),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_18),
.CI(n_19),
.CON(n_96),
.SN(n_96)
);


endmodule