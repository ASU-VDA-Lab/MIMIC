module fake_netlist_6_674_n_184 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_184);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_184;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_1),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_32),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_7),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_9),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_10),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_33),
.B(n_51),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_75),
.B(n_73),
.C(n_71),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_66),
.B(n_56),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_45),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_43),
.B1(n_53),
.B2(n_50),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_40),
.B(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_50),
.C(n_34),
.Y(n_86)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_52),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_11),
.Y(n_87)
);

O2A1O1Ixp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_41),
.B(n_37),
.C(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_15),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_90)
);

NAND2x1p5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_29),
.Y(n_91)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_75),
.A3(n_73),
.B1(n_63),
.B2(n_68),
.C(n_71),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_72),
.B(n_59),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_59),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_69),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_83),
.Y(n_98)
);

NOR2xp67_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_69),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_64),
.B1(n_61),
.B2(n_74),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_61),
.B(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_94),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_91),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_111),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_104),
.Y(n_125)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_99),
.B(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_104),
.B1(n_115),
.B2(n_64),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_105),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_122),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_105),
.Y(n_142)
);

AOI222xp33_ASAP7_75t_SL g143 ( 
.A1(n_135),
.A2(n_90),
.B1(n_87),
.B2(n_64),
.C1(n_93),
.C2(n_92),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_87),
.C(n_88),
.Y(n_144)
);

NOR3x1_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_131),
.C(n_132),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_131),
.Y(n_148)
);

OAI211xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_77),
.B(n_136),
.C(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_129),
.Y(n_150)
);

AOI211xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_127),
.B(n_99),
.C(n_97),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_126),
.Y(n_152)
);

NOR4xp75_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_97),
.C(n_100),
.D(n_126),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_126),
.B1(n_100),
.B2(n_109),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_80),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_112),
.B1(n_113),
.B2(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_80),
.Y(n_166)
);

AO21x2_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_112),
.B(n_113),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_112),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_113),
.C(n_102),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NAND4xp25_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_81),
.C(n_111),
.D(n_107),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_163),
.B1(n_81),
.B2(n_111),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_81),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_81),
.Y(n_176)
);

NAND5xp2_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_81),
.C(n_107),
.D(n_169),
.E(n_172),
.Y(n_177)
);

OAI22x1_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_107),
.B1(n_171),
.B2(n_172),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_107),
.C(n_166),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_167),
.B(n_107),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_107),
.B(n_174),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_177),
.B(n_176),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_R g184 ( 
.A1(n_183),
.A2(n_175),
.B1(n_180),
.B2(n_181),
.C(n_60),
.Y(n_184)
);


endmodule