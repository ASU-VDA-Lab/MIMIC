module fake_jpeg_15211_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_33),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_2),
.C(n_3),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_31),
.C(n_17),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_19),
.C(n_17),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_32),
.B1(n_26),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_27),
.B1(n_34),
.B2(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_54),
.Y(n_80)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_38),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_20),
.B1(n_32),
.B2(n_26),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_46),
.B1(n_22),
.B2(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_28),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_36),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_16),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_42),
.B1(n_26),
.B2(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_63),
.B1(n_58),
.B2(n_16),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_58),
.B1(n_25),
.B2(n_19),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_62),
.B(n_56),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_24),
.B(n_22),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_55),
.B(n_48),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_71),
.C(n_74),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_94),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_56),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_103),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_93),
.B1(n_71),
.B2(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_46),
.B1(n_61),
.B2(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_83),
.B(n_79),
.C(n_66),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_81),
.B(n_65),
.C(n_80),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_57),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_67),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_126),
.B1(n_19),
.B2(n_31),
.Y(n_145)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_120),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_121),
.B(n_102),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_123),
.B(n_88),
.C(n_105),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_74),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_122),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_71),
.B1(n_16),
.B2(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_25),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_97),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_134),
.C(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_131),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_98),
.B1(n_86),
.B2(n_100),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_96),
.B1(n_93),
.B2(n_103),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_140),
.B1(n_121),
.B2(n_106),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_146),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_92),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_87),
.B(n_91),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_87),
.C(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_25),
.B1(n_19),
.B2(n_17),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_123),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_119),
.B1(n_115),
.B2(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_158),
.B1(n_161),
.B2(n_140),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_155),
.C(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_134),
.B(n_131),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_162),
.B(n_157),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_119),
.B(n_115),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_141),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_173),
.C(n_153),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_154),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_170),
.B(n_172),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_136),
.B(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_130),
.B1(n_146),
.B2(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_3),
.B(n_4),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_31),
.CI(n_4),
.CON(n_178),
.SN(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_152),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_178),
.B1(n_170),
.B2(n_176),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_185),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_175),
.B(n_166),
.Y(n_192)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_148),
.C(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_190),
.C(n_170),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_167),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_3),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_6),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_15),
.C(n_14),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_196),
.C(n_198),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_199),
.B(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_189),
.B1(n_180),
.B2(n_164),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_188),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_15),
.B(n_14),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_183),
.B(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_185),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_13),
.B(n_8),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_184),
.A3(n_186),
.B1(n_182),
.B2(n_187),
.C1(n_12),
.C2(n_13),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_197),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_207),
.B(n_10),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.C(n_9),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_200),
.B1(n_206),
.B2(n_195),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_6),
.B(n_9),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_215),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_211),
.B(n_6),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_9),
.B(n_11),
.C(n_217),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_11),
.Y(n_219)
);


endmodule