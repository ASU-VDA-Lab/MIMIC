module fake_jpeg_11634_n_460 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_460);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_460;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_9),
.B(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_58),
.Y(n_176)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_60),
.Y(n_123)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g161 ( 
.A(n_62),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_64),
.Y(n_178)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_70),
.B(n_78),
.Y(n_140)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_94),
.Y(n_118)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_15),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_18),
.B(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_97),
.Y(n_121)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_89),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_92),
.Y(n_166)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_26),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_102),
.Y(n_153)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_107),
.Y(n_119)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_103),
.B(n_104),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_26),
.B(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_43),
.A2(n_13),
.B1(n_12),
.B2(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_31),
.B1(n_34),
.B2(n_56),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_13),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_111),
.B(n_23),
.Y(n_141)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_115),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_50),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_120),
.B(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_180),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_28),
.B1(n_25),
.B2(n_37),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_126),
.A2(n_167),
.B1(n_161),
.B2(n_125),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_28),
.B1(n_25),
.B2(n_38),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_123),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_31),
.B1(n_34),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_145),
.B1(n_165),
.B2(n_168),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_50),
.B1(n_38),
.B2(n_54),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_78),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_138),
.B(n_139),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_62),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_141),
.B(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_27),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_144),
.B(n_148),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_50),
.B1(n_38),
.B2(n_54),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_84),
.A2(n_27),
.B(n_49),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_167),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_104),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_53),
.B1(n_48),
.B2(n_44),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_57),
.A2(n_22),
.B1(n_6),
.B2(n_7),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_66),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_173),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_115),
.A2(n_22),
.B1(n_6),
.B2(n_7),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_107),
.B1(n_109),
.B2(n_8),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_81),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_95),
.B(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_184),
.Y(n_273)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_185),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_124),
.A2(n_4),
.B(n_8),
.C(n_10),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_190),
.A2(n_199),
.B(n_204),
.C(n_222),
.Y(n_267)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_192),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_161),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_195),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_196),
.A2(n_209),
.B1(n_213),
.B2(n_219),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_128),
.A2(n_8),
.B1(n_11),
.B2(n_155),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_198),
.Y(n_290)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_140),
.A2(n_8),
.A3(n_118),
.B1(n_121),
.B2(n_119),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_240),
.Y(n_246)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

BUFx24_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_135),
.A3(n_143),
.B1(n_146),
.B2(n_123),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_126),
.A2(n_145),
.B1(n_172),
.B2(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_211),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_174),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_212),
.B(n_241),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_132),
.B1(n_157),
.B2(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_223),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_161),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_217),
.A2(n_230),
.B1(n_215),
.B2(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_152),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_164),
.C(n_150),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_225),
.C(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_181),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_150),
.B(n_116),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g226 ( 
.A1(n_159),
.A2(n_133),
.B1(n_170),
.B2(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_234),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_133),
.A2(n_162),
.B1(n_125),
.B2(n_137),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_217),
.B1(n_223),
.B2(n_200),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_116),
.A2(n_183),
.B1(n_171),
.B2(n_176),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_229),
.B1(n_236),
.B2(n_186),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_137),
.A2(n_162),
.B1(n_142),
.B2(n_171),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_142),
.A2(n_183),
.B1(n_166),
.B2(n_176),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_152),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_159),
.B(n_131),
.C(n_182),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_182),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_242),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_182),
.A2(n_131),
.B1(n_149),
.B2(n_46),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_149),
.Y(n_237)
);

AO22x2_ASAP7_75t_L g238 ( 
.A1(n_149),
.A2(n_132),
.B1(n_163),
.B2(n_141),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_240),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_118),
.B(n_134),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_202),
.Y(n_266)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_244),
.B(n_205),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_280),
.C(n_289),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_272),
.B1(n_274),
.B2(n_226),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_214),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_266),
.Y(n_295)
);

AOI32xp33_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_197),
.A3(n_215),
.B1(n_238),
.B2(n_201),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_265),
.B(n_249),
.Y(n_327)
);

NAND2x1p5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_238),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_277),
.B(n_291),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_187),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_270),
.B(n_278),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_233),
.B1(n_197),
.B2(n_219),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_189),
.B(n_221),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_194),
.B(n_241),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_242),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_208),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_282),
.B(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_191),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_190),
.B(n_237),
.C(n_229),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_193),
.A2(n_243),
.B(n_226),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_203),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_224),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_297),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_296),
.A2(n_321),
.B1(n_297),
.B2(n_295),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_244),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_298),
.B(n_309),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_245),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_300),
.B(n_303),
.Y(n_343)
);

OR2x2_ASAP7_75t_SL g301 ( 
.A(n_268),
.B(n_261),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_261),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_273),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_264),
.A2(n_259),
.B1(n_290),
.B2(n_277),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_304),
.A2(n_306),
.B1(n_322),
.B2(n_329),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_264),
.A2(n_268),
.B1(n_257),
.B2(n_267),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_273),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_308),
.B(n_310),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_246),
.B(n_248),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_250),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_275),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_312),
.B(n_314),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_291),
.B(n_290),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_328),
.B(n_298),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_262),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_262),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_249),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_324),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_252),
.B(n_251),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_320),
.Y(n_347)
);

A2O1A1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_267),
.A2(n_289),
.B(n_258),
.C(n_280),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_258),
.B1(n_286),
.B2(n_288),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_271),
.A2(n_251),
.B1(n_288),
.B2(n_287),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_283),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_325),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_258),
.B(n_256),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_283),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_249),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_327),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_306),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_254),
.A2(n_269),
.B1(n_279),
.B2(n_260),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_254),
.A2(n_269),
.B1(n_279),
.B2(n_260),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_330),
.A2(n_344),
.B(n_311),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_322),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_342),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_309),
.C(n_311),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_324),
.C(n_321),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_312),
.Y(n_337)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_339),
.B(n_300),
.Y(n_369)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_302),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_305),
.A2(n_329),
.B1(n_317),
.B2(n_313),
.Y(n_346)
);

OAI22x1_ASAP7_75t_L g358 ( 
.A1(n_346),
.A2(n_296),
.B1(n_305),
.B2(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_353),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_349),
.A2(n_304),
.B1(n_333),
.B2(n_342),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_326),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_301),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_299),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_375),
.B(n_377),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_299),
.C(n_301),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_373),
.C(n_364),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_368),
.B1(n_374),
.B2(n_376),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_351),
.A2(n_296),
.B1(n_299),
.B2(n_305),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_363),
.A2(n_379),
.B1(n_353),
.B2(n_341),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_367),
.B(n_369),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_305),
.B1(n_294),
.B2(n_320),
.Y(n_368)
);

OAI22x1_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_321),
.B1(n_320),
.B2(n_295),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_347),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_310),
.Y(n_372)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_317),
.B1(n_307),
.B2(n_319),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_330),
.A2(n_328),
.B(n_308),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_307),
.B1(n_303),
.B2(n_315),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_347),
.A2(n_328),
.B(n_352),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_351),
.A2(n_331),
.B1(n_352),
.B2(n_341),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_381),
.A2(n_375),
.B(n_368),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_383),
.A2(n_392),
.B1(n_362),
.B2(n_376),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_366),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_389),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_370),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_395),
.C(n_397),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_363),
.A2(n_331),
.B1(n_337),
.B2(n_350),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_343),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_343),
.Y(n_409)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_396),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_344),
.C(n_354),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_366),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_344),
.C(n_345),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_377),
.A2(n_350),
.B(n_338),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_398),
.A2(n_374),
.B(n_359),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_402),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_385),
.A2(n_379),
.B1(n_359),
.B2(n_358),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_371),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_412),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_385),
.B1(n_386),
.B2(n_389),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_357),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_408),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_371),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_409),
.B(n_415),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_361),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_390),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_355),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_410),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_416),
.A2(n_394),
.B(n_407),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g417 ( 
.A(n_411),
.B(n_367),
.CI(n_390),
.CON(n_417),
.SN(n_417)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_417),
.A2(n_423),
.B1(n_424),
.B2(n_392),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_355),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_419),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_SL g422 ( 
.A(n_403),
.B(n_408),
.Y(n_422)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_426),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_406),
.B(n_383),
.Y(n_427)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_425),
.A2(n_380),
.B(n_412),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_429),
.A2(n_400),
.B(n_407),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_416),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_436),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_398),
.B1(n_382),
.B2(n_358),
.Y(n_442)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_420),
.A2(n_387),
.B1(n_396),
.B2(n_382),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_411),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_438),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_SL g438 ( 
.A1(n_434),
.A2(n_380),
.B(n_405),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_427),
.C(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_440),
.B(n_444),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_442),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_429),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_418),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_439),
.A2(n_423),
.B1(n_436),
.B2(n_402),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_447),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_441),
.B(n_372),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_421),
.C(n_435),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_SL g452 ( 
.A1(n_446),
.A2(n_443),
.B(n_417),
.C(n_438),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_452),
.A2(n_453),
.B(n_454),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_450),
.A2(n_413),
.B(n_384),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_451),
.B(n_449),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_456),
.A2(n_452),
.B(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_457),
.B(n_455),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_458),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_401),
.B1(n_384),
.B2(n_365),
.Y(n_460)
);


endmodule