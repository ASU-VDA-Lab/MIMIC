module fake_netlist_1_12133_n_654 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_654);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_654;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_577;
wire n_216;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx10_ASAP7_75t_L g77 ( .A(n_0), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_45), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_46), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_38), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_7), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_35), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_62), .B(n_26), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_42), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_41), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_33), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_34), .Y(n_87) );
INVx1_ASAP7_75t_SL g88 ( .A(n_23), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_59), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_20), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_58), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_30), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_64), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_19), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_31), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_51), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_29), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_39), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_43), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_47), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
INVxp33_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_1), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_7), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_52), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_5), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_24), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_18), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_66), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_22), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_65), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_91), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_91), .B(n_1), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_95), .B(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_114), .Y(n_125) );
NAND2xp33_ASAP7_75t_L g126 ( .A(n_98), .B(n_76), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_114), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_81), .B(n_3), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_89), .A2(n_4), .B1(n_5), .B2(n_8), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_92), .B(n_8), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_102), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_94), .B(n_9), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_105), .B(n_9), .Y(n_142) );
NOR2x1_ASAP7_75t_L g143 ( .A(n_111), .B(n_10), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_94), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_112), .B(n_10), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_104), .A2(n_48), .B(n_74), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_103), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_101), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_78), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_118), .B(n_12), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_77), .B(n_13), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_96), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
NOR2x1p5_ASAP7_75t_L g160 ( .A(n_130), .B(n_108), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_134), .B(n_100), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_134), .B(n_120), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_152), .B(n_93), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_122), .A2(n_119), .B1(n_107), .B2(n_109), .Y(n_168) );
INVx6_ASAP7_75t_L g169 ( .A(n_122), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_132), .B(n_116), .Y(n_173) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_152), .B(n_93), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_130), .B(n_117), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_123), .B(n_77), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_123), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_142), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_124), .B(n_97), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_121), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_121), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_138), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_124), .B(n_97), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_133), .B(n_100), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_142), .B(n_77), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_190), .B(n_125), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_191), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_191), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_166), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_174), .B(n_178), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_163), .B(n_157), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_191), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_191), .Y(n_210) );
AOI21x1_ASAP7_75t_L g211 ( .A1(n_188), .A2(n_147), .B(n_137), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_183), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_183), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_176), .B(n_157), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_183), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_174), .B(n_135), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_181), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_174), .B(n_135), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_173), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_181), .B(n_154), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g224 ( .A1(n_201), .A2(n_150), .B1(n_154), .B2(n_106), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_169), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_174), .A2(n_87), .B1(n_79), .B2(n_99), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_201), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_184), .A2(n_126), .B1(n_129), .B2(n_153), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_169), .Y(n_230) );
XNOR2xp5_ASAP7_75t_L g231 ( .A(n_160), .B(n_150), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_160), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_169), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_180), .B(n_136), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_169), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_158), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_169), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_189), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_189), .B(n_136), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_178), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_178), .B(n_133), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_187), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_187), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_178), .B(n_137), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_192), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_165), .B(n_139), .Y(n_249) );
NOR2xp33_ASAP7_75t_R g250 ( .A(n_173), .B(n_108), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_197), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_199), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_173), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_164), .B(n_139), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_218), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_225), .Y(n_257) );
BUFx12f_ASAP7_75t_L g258 ( .A(n_232), .Y(n_258) );
AND2x4_ASAP7_75t_SL g259 ( .A(n_218), .B(n_164), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_214), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_235), .A2(n_179), .B(n_194), .C(n_196), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_227), .Y(n_263) );
BUFx8_ASAP7_75t_SL g264 ( .A(n_232), .Y(n_264) );
BUFx4f_ASAP7_75t_L g265 ( .A(n_202), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_222), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_207), .A2(n_200), .B(n_164), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_225), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
O2A1O1Ixp5_ASAP7_75t_SL g271 ( .A1(n_246), .A2(n_149), .B(n_151), .C(n_155), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_222), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_244), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_250), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_202), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_212), .A2(n_200), .B(n_188), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_221), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_207), .A2(n_200), .B(n_179), .Y(n_279) );
AO21x1_ASAP7_75t_L g280 ( .A1(n_211), .A2(n_200), .B(n_159), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
AND3x1_ASAP7_75t_SL g282 ( .A(n_231), .B(n_110), .C(n_113), .Y(n_282) );
INVx5_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_254), .B(n_179), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_206), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_249), .B(n_173), .Y(n_286) );
BUFx2_ASAP7_75t_SL g287 ( .A(n_242), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_217), .A2(n_147), .B(n_168), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_214), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_223), .B(n_196), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_241), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_217), .A2(n_147), .B(n_159), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_254), .B(n_193), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_244), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_242), .A2(n_155), .B1(n_149), .B2(n_151), .Y(n_295) );
AND3x4_ASAP7_75t_L g296 ( .A(n_231), .B(n_143), .C(n_127), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_226), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_203), .B(n_195), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_240), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_230), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
O2A1O1Ixp5_ASAP7_75t_SL g302 ( .A1(n_253), .A2(n_117), .B(n_175), .C(n_177), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g303 ( .A1(n_285), .A2(n_224), .B1(n_229), .B2(n_252), .C(n_215), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_268), .A2(n_220), .B(n_243), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_280), .A2(n_247), .B(n_243), .Y(n_305) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_280), .A2(n_171), .B(n_172), .Y(n_306) );
INVx6_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_279), .A2(n_220), .B(n_247), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_302), .A2(n_248), .B(n_182), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_302), .A2(n_182), .B(n_170), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_291), .A2(n_208), .B1(n_237), .B2(n_238), .Y(n_312) );
INVxp33_ASAP7_75t_L g313 ( .A(n_260), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_257), .Y(n_314) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_262), .A2(n_140), .B(n_177), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_292), .A2(n_186), .B(n_182), .Y(n_316) );
BUFx8_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_298), .B(n_221), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_288), .A2(n_186), .B(n_170), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_277), .A2(n_186), .B(n_170), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_271), .A2(n_167), .B(n_245), .Y(n_321) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_262), .A2(n_140), .B(n_175), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_256), .B(n_251), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_261), .A2(n_167), .B(n_245), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_289), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_257), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_259), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
AO31x2_ASAP7_75t_L g329 ( .A1(n_295), .A2(n_145), .A3(n_172), .B(n_171), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_286), .A2(n_167), .B(n_162), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_269), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_298), .A2(n_195), .B1(n_194), .B2(n_198), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_261), .A2(n_162), .B(n_210), .Y(n_333) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_128), .B(n_209), .Y(n_334) );
INVx3_ASAP7_75t_SL g335 ( .A(n_259), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_319), .A2(n_316), .B(n_320), .Y(n_336) );
NOR2x1_ASAP7_75t_SL g337 ( .A(n_332), .B(n_287), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_332), .A2(n_290), .B(n_281), .C(n_275), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_314), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_303), .A2(n_296), .B1(n_263), .B2(n_173), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_313), .A2(n_296), .B1(n_263), .B2(n_173), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_304), .A2(n_290), .B(n_265), .C(n_297), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_307), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_331), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_335), .A2(n_265), .B1(n_299), .B2(n_270), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_318), .A2(n_173), .B1(n_258), .B2(n_300), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_323), .A2(n_156), .B1(n_141), .B2(n_198), .C(n_282), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_318), .B(n_294), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
CKINVDCx12_ASAP7_75t_R g352 ( .A(n_317), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_305), .A2(n_273), .B(n_294), .Y(n_353) );
OAI22x1_ASAP7_75t_L g354 ( .A1(n_335), .A2(n_143), .B1(n_283), .B2(n_293), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_326), .B(n_278), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_312), .A2(n_198), .B1(n_236), .B2(n_239), .C(n_233), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_258), .B1(n_238), .B2(n_237), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_326), .B(n_265), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_317), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_198), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_331), .B(n_278), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_339), .B(n_334), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_337), .A2(n_317), .B1(n_327), .B2(n_307), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_351), .B(n_334), .Y(n_366) );
AOI33xp33_ASAP7_75t_L g367 ( .A1(n_347), .A2(n_88), .A3(n_327), .B1(n_205), .B2(n_204), .B3(n_15), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_351), .B(n_329), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_361), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_361), .B(n_334), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_347), .B(n_329), .Y(n_373) );
OAI221xp5_ASAP7_75t_SL g374 ( .A1(n_340), .A2(n_309), .B1(n_82), .B2(n_80), .C(n_83), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_338), .B(n_315), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_344), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_349), .B(n_315), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_334), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_348), .B(n_329), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_360), .B(n_315), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_341), .A2(n_322), .B1(n_221), .B2(n_284), .C(n_238), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_337), .B(n_308), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_358), .B(n_308), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_358), .B(n_308), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_350), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_360), .B(n_362), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_345), .B(n_264), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_378), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_368), .B(n_329), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_329), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_367), .A2(n_346), .B1(n_357), .B2(n_342), .C(n_356), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_371), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_363), .B(n_322), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_388), .A2(n_359), .B1(n_355), .B2(n_354), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_381), .B(n_322), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_381), .B(n_355), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_364), .A2(n_356), .B1(n_343), .B2(n_307), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_380), .B(n_343), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_353), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_366), .B(n_306), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_373), .A2(n_354), .B1(n_185), .B2(n_161), .C(n_284), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_382), .B(n_306), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_390), .A2(n_307), .B1(n_306), .B2(n_293), .C(n_266), .Y(n_414) );
OAI31xp33_ASAP7_75t_L g415 ( .A1(n_374), .A2(n_393), .A3(n_389), .B(n_380), .Y(n_415) );
OAI321xp33_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_161), .A3(n_185), .B1(n_289), .B2(n_272), .C(n_267), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_376), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_384), .B(n_305), .C(n_325), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_379), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_370), .B(n_306), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_369), .B(n_330), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_370), .Y(n_425) );
NOR2xp33_ASAP7_75t_SL g426 ( .A(n_385), .B(n_264), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_392), .B(n_330), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_385), .B(n_336), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_382), .B(n_336), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_379), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_392), .B(n_330), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_372), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_372), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_386), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_391), .B(n_336), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_391), .B(n_325), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_422), .B(n_391), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_429), .B(n_377), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_425), .B(n_383), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_425), .B(n_383), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_429), .B(n_377), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_403), .B(n_391), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_394), .B(n_372), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_372), .Y(n_445) );
NOR2x1p5_ASAP7_75t_L g446 ( .A(n_420), .B(n_385), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_396), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_395), .B(n_375), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_395), .B(n_385), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_434), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_395), .B(n_387), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_396), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_400), .B(n_410), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_400), .B(n_387), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_387), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_405), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_410), .B(n_387), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_411), .B(n_386), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_405), .B(n_386), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_411), .B(n_386), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_401), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_423), .B(n_319), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_397), .B(n_310), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_401), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_415), .B(n_301), .C(n_261), .D(n_266), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_401), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_432), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_397), .B(n_310), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_423), .B(n_320), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_413), .B(n_321), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_413), .B(n_321), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_402), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_398), .B(n_316), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_407), .B(n_308), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_415), .B(n_301), .C(n_266), .D(n_325), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_426), .B(n_283), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_420), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_398), .B(n_325), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_407), .B(n_283), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_417), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_435), .B(n_324), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_409), .B(n_283), .Y(n_487) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_418), .B(n_289), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_418), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_435), .B(n_324), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_418), .B(n_311), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_408), .A2(n_237), .B1(n_238), .B2(n_333), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_453), .B(n_428), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_438), .B(n_427), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_438), .B(n_431), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_450), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_453), .B(n_406), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_451), .B(n_428), .Y(n_499) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_468), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_451), .B(n_428), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_447), .Y(n_503) );
AND3x2_ASAP7_75t_L g504 ( .A(n_479), .B(n_430), .C(n_419), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
NOR2xp67_ASAP7_75t_L g506 ( .A(n_466), .B(n_416), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_442), .B(n_406), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_454), .B(n_433), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_465), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
NAND2xp33_ASAP7_75t_L g512 ( .A(n_446), .B(n_424), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_452), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_446), .B(n_421), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_454), .B(n_433), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g516 ( .A1(n_459), .A2(n_404), .B1(n_399), .B2(n_414), .C(n_412), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_439), .B(n_421), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_455), .B(n_433), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_476), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_437), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_455), .B(n_421), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_439), .B(n_420), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_443), .B(n_436), .Y(n_523) );
NOR2xp67_ASAP7_75t_SL g524 ( .A(n_478), .B(n_276), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_440), .B(n_311), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_443), .B(n_185), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_478), .A2(n_333), .B1(n_276), .B2(n_161), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_449), .B(n_185), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_442), .B(n_185), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_449), .B(n_185), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_440), .B(n_161), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_452), .B(n_161), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_463), .B(n_17), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_456), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_456), .B(n_161), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_457), .B(n_21), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_461), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_445), .B(n_25), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_483), .B(n_27), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_445), .B(n_28), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_480), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_458), .B(n_32), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_484), .B(n_272), .C(n_267), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_461), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_457), .B(n_460), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_458), .B(n_36), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_464), .B(n_37), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_505), .A2(n_463), .B(n_460), .C(n_492), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_506), .A2(n_488), .B(n_487), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_520), .Y(n_551) );
OAI221xp5_ASAP7_75t_L g552 ( .A1(n_516), .A2(n_463), .B1(n_464), .B2(n_470), .C(n_477), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_500), .A2(n_512), .B(n_548), .C(n_537), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_497), .B(n_463), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_495), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_504), .B(n_470), .C(n_472), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_493), .B(n_448), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_514), .B(n_482), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_512), .A2(n_483), .B(n_476), .C(n_444), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_546), .B(n_448), .Y(n_563) );
OAI31xp33_ASAP7_75t_L g564 ( .A1(n_543), .A2(n_473), .A3(n_472), .B(n_462), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_514), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_543), .A2(n_473), .B1(n_462), .B2(n_471), .Y(n_566) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_548), .A2(n_488), .B(n_469), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_527), .A2(n_469), .B(n_485), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_501), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_540), .A2(n_482), .B1(n_485), .B2(n_489), .Y(n_570) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_514), .B(n_475), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_503), .Y(n_572) );
NAND3x1_ASAP7_75t_L g573 ( .A(n_547), .B(n_490), .C(n_486), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_509), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_547), .A2(n_522), .B1(n_517), .B2(n_496), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_510), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_523), .B(n_471), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_523), .B(n_481), .Y(n_578) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_524), .A2(n_491), .B(n_490), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
OAI21xp33_ASAP7_75t_SL g581 ( .A1(n_493), .A2(n_489), .B(n_481), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_496), .B(n_489), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_539), .A2(n_486), .B(n_481), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_544), .A2(n_475), .B(n_474), .C(n_467), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_539), .A2(n_475), .B(n_474), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_498), .B(n_474), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_494), .B(n_467), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_507), .A2(n_467), .B1(n_276), .B2(n_219), .Y(n_588) );
OAI222xp33_ASAP7_75t_L g589 ( .A1(n_507), .A2(n_44), .B1(n_49), .B2(n_50), .C1(n_53), .C2(n_55), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_564), .A2(n_513), .B1(n_535), .B2(n_545), .C(n_538), .Y(n_590) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_559), .A2(n_510), .B(n_532), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_551), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_576), .Y(n_593) );
OAI221xp5_ASAP7_75t_SL g594 ( .A1(n_552), .A2(n_502), .B1(n_499), .B2(n_541), .C(n_521), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_581), .A2(n_499), .B(n_502), .C(n_541), .Y(n_595) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_585), .A2(n_534), .B(n_521), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_565), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_558), .B(n_508), .Y(n_598) );
NAND2xp33_ASAP7_75t_L g599 ( .A(n_573), .B(n_526), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_558), .B(n_526), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_576), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_571), .B(n_534), .Y(n_602) );
NAND2x1_ASAP7_75t_L g603 ( .A(n_554), .B(n_534), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_553), .A2(n_528), .B(n_530), .C(n_518), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_569), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_578), .B(n_508), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_550), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_555), .B(n_515), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_555), .B(n_515), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_563), .B(n_518), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_580), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_575), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_609), .A2(n_549), .B(n_589), .C(n_562), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_599), .A2(n_584), .B(n_583), .C(n_561), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_605), .B(n_607), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_601), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_614), .B(n_577), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_590), .A2(n_570), .B1(n_582), .B2(n_587), .C(n_567), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_601), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_609), .B(n_560), .Y(n_622) );
OAI22xp33_ASAP7_75t_SL g623 ( .A1(n_594), .A2(n_603), .B1(n_602), .B2(n_592), .Y(n_623) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_596), .B(n_566), .Y(n_624) );
CKINVDCx16_ASAP7_75t_R g625 ( .A(n_600), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_604), .A2(n_579), .B(n_589), .C(n_568), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_595), .A2(n_586), .B(n_588), .C(n_528), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_597), .B(n_530), .Y(n_628) );
AOI21x1_ASAP7_75t_L g629 ( .A1(n_591), .A2(n_531), .B(n_574), .Y(n_629) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_615), .A2(n_591), .B(n_598), .C(n_611), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_617), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_623), .A2(n_598), .B1(n_606), .B2(n_613), .C(n_610), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_616), .A2(n_612), .B(n_593), .C(n_608), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_626), .B(n_525), .C(n_529), .D(n_533), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_624), .A2(n_557), .B1(n_532), .B2(n_529), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_628), .A2(n_536), .B1(n_276), .B2(n_216), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_627), .A2(n_56), .B(n_57), .Y(n_637) );
NOR4xp75_ASAP7_75t_L g638 ( .A(n_629), .B(n_60), .C(n_63), .D(n_67), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_631), .B(n_622), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_636), .Y(n_640) );
AND3x4_ASAP7_75t_L g641 ( .A(n_638), .B(n_625), .C(n_621), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_633), .B(n_618), .C(n_619), .Y(n_642) );
NAND2xp33_ASAP7_75t_SL g643 ( .A(n_635), .B(n_617), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_641), .A2(n_632), .B1(n_630), .B2(n_637), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_640), .B(n_634), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_639), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_646), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_645), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_647), .Y(n_649) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_648), .A2(n_644), .B1(n_642), .B2(n_643), .Y(n_650) );
OAI22xp5_ASAP7_75t_SL g651 ( .A1(n_650), .A2(n_620), .B1(n_70), .B2(n_71), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_651), .B(n_649), .C(n_72), .D(n_75), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_652), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_213), .B(n_69), .Y(n_654) );
endmodule